
module iir_filter ( clk, rst_n, vIn, dIn, coeffs_fb, coeffs_ff, dOut, vOut );
  input [11:0] dIn;
  input [47:0] coeffs_fb;
  input [95:0] coeffs_ff;
  output [11:0] dOut;
  input clk, rst_n, vIn;
  output vOut;
  wire   sw_regs_en_int, delayed_controls_0__1_, delayed_controls_1__0_,
         delayed_controls_1__1_, delayed_controls_2__0_, DP_N17, DP_N16,
         DP_N15, DP_N14, DP_N13, DP_N12, DP_N11, DP_N10, DP_N9, DP_N8, DP_N7,
         DP_N6, DP_N5, DP_N4, DP_N3, DP_N2, DP_y_0_, DP_y_1_, DP_y_2_, DP_y_3_,
         DP_y_4_, DP_y_5_, DP_y_6_, DP_y_7_, DP_y_8_, DP_y_9_, DP_y_10_,
         DP_y_11_, DP_y_23, DP_sw1_0_, DP_sw1_1_, DP_sw1_2_, DP_sw1_3_,
         DP_sw1_4_, DP_sw1_5_, DP_sw1_6_, DP_sw1_7_, DP_sw1_8_, DP_sw1_9_,
         DP_sw1_10_, DP_sw1_11_, DP_sw1_12_, DP_sw1_13_, DP_sw1_14_,
         DP_sw1_15_, DP_sw1_16_, DP_sw1_17_, DP_sw1_18_, DP_sw1_19_,
         DP_sw1_20_, DP_sw1_21_, DP_sw1_22_, DP_sw1_23_, DP_sw0_0_, DP_sw0_1_,
         DP_sw0_2_, DP_sw0_3_, DP_sw0_4_, DP_sw0_5_, DP_sw0_6_, DP_sw0_7_,
         DP_sw0_8_, DP_sw0_9_, DP_sw0_10_, DP_sw0_11_, DP_sw0_12_, DP_sw0_13_,
         DP_sw0_14_, DP_sw0_15_, DP_sw0_16_, DP_sw0_17_, DP_sw0_18_,
         DP_sw0_19_, DP_sw0_20_, DP_sw0_21_, DP_sw0_22_, DP_sw0_23_, DP_w_0_,
         DP_w_1_, DP_w_2_, DP_w_3_, DP_w_4_, DP_w_5_, DP_w_6_, DP_w_7_,
         DP_w_8_, DP_w_9_, DP_w_10_, DP_w_11_, DP_w_12_, DP_w_13_, DP_w_14_,
         DP_w_15_, DP_w_16_, DP_w_17_, DP_w_18_, DP_w_19_, DP_w_20_, DP_w_21_,
         DP_w_22_, DP_w_23_, DP_N1, DP_N0, DP_reg_in_N0,
         DP_reg_coeff_fb_i_1_N0, DP_reg_coeff_fb_i_2_N0, DP_reg_b_i_0_N0,
         DP_reg_b_i_1_N0, DP_reg_b_i_2_N0, DP_reg_b_i_3_N0, DP_reg_sw0_N0,
         DP_reg_sw1_N0, DP_reg_sw2_N0, DP_reg_ret0_N0, DP_reg_ret1_N0,
         DP_reg_pipe00_N0, DP_reg_pipe01_N0, DP_reg_pipe02_N0,
         DP_reg_pipe03_N0, DP_reg_pipe10_N0, DP_reg_pipe11_N0,
         DP_reg_pipe12_N0, DP_reg_pipe13_N0, DP_reg_out_N0, CU_N18, CU_N17,
         CU_N16, CU_N15, CU_N14, CU_N13, CU_N12, CU_N11, CU_N10, CU_N9, CU_N8,
         CU_N7, CU_N6, CU_N5, CU_N4, CU_presentState_0_, CU_presentState_1_,
         CU_N3, CU_N2, CU_N1, CU_N0, reg_delay_0_N0, reg_delay_1_N0;
  wire   [0:23] DP_ff;
  wire   [0:23] DP_ff_part;
  wire   [0:23] DP_fb;
  wire   [0:11] DP_y_out;
  wire   [0:23] DP_pipe13;
  wire   [0:23] DP_pipe0_coeff_pipe03;
  wire   [0:23] DP_pipe12;
  wire   [0:23] DP_pipe0_coeff_pipe02;
  wire   [0:23] DP_pipe11;
  wire   [0:23] DP_pipe0_coeff_pipe01;
  wire   [0:23] DP_pipe10;
  wire   [0:23] DP_pipe0_coeff_pipe00;
  wire   [0:23] DP_pipe03;
  wire   [0:23] DP_pipe02;
  wire   [0:23] DP_pipe01;
  wire   [0:23] DP_pipe00;
  wire   [0:23] DP_ret1;
  wire   [0:23] DP_sw1_coeff_ret1;
  wire   [0:23] DP_ret0;
  wire   [0:23] DP_sw0_coeff_ret0;
  wire   [0:23] DP_sw2;
  wire   [95:0] DP_coeffs_ff_int;
  wire   [47:0] DP_coeffs_fb_int;
  wire   [0:11] DP_x;
  wire   [0:1] CU_nextState;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154;

  GTECH_NOT DP_I_1 ( .A(DP_N4), .Z(DP_N5) );
  GTECH_BUF DP_B_2 ( .A(DP_N3) );
  GTECH_NOT DP_I_0 ( .A(DP_N2), .Z(DP_N3) );
  GTECH_BUF DP_B_1 ( .A(DP_N2), .Z(DP_N1) );
  SELECT_OP DP_C38 ( .DATA1({1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1}), .DATA2({DP_N17, DP_N16, DP_N15, DP_N14, 
        DP_N13, DP_N12, DP_N11, DP_N10, DP_N9, DP_N8, DP_N7, DP_N6}), 
        .CONTROL1(DP_N1), .CONTROL2(DP_N3), .Z({DP_y_out[11], DP_y_out[10], 
        DP_y_out[9], DP_y_out[8], DP_y_out[7], DP_y_out[6], DP_y_out[5], 
        DP_y_out[4], DP_y_out[3], DP_y_out[2], DP_y_out[1], DP_y_out[0]}) );
  GTECH_BUF DP_B_0 ( .A(DP_N4), .Z(DP_N0) );
  SELECT_OP DP_C37 ( .DATA1({1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .DATA2({DP_y_23, DP_y_10_, DP_y_9_, DP_y_8_, 
        DP_y_7_, DP_y_6_, DP_y_5_, DP_y_4_, DP_y_3_, DP_y_2_, DP_y_1_, DP_y_0_}), .CONTROL1(DP_N0), .CONTROL2(DP_N5), .Z({DP_N17, DP_N16, DP_N15, DP_N14, 
        DP_N13, DP_N12, DP_N11, DP_N10, DP_N9, DP_N8, DP_N7, DP_N6}) );
  ADD_TC_OP DP_add_223 ( .A({DP_pipe10[23], DP_pipe10[22], DP_pipe10[21], 
        DP_pipe10[20], DP_pipe10[19], DP_pipe10[18], DP_pipe10[17], 
        DP_pipe10[16], DP_pipe10[15], DP_pipe10[14], DP_pipe10[13], 
        DP_pipe10[12], DP_pipe10[11], DP_pipe10[10], DP_pipe10[9], 
        DP_pipe10[8], DP_pipe10[7], DP_pipe10[6], DP_pipe10[5], DP_pipe10[4], 
        DP_pipe10[3], DP_pipe10[2], DP_pipe10[1], DP_pipe10[0]}), .B({
        DP_ff[23], DP_ff[22], DP_ff[21], DP_ff[20], DP_ff[19], DP_ff[18], 
        DP_ff[17], DP_ff[16], DP_ff[15], DP_ff[14], DP_ff[13], DP_ff[12], 
        DP_ff[11], DP_ff[10], DP_ff[9], DP_ff[8], DP_ff[7], DP_ff[6], DP_ff[5], 
        DP_ff[4], DP_ff[3], DP_ff[2], DP_ff[1], DP_ff[0]}), .Z({DP_y_23, 
        DP_y_11_, DP_y_10_, DP_y_9_, DP_y_8_, DP_y_7_, DP_y_6_, DP_y_5_, 
        DP_y_4_, DP_y_3_, DP_y_2_, DP_y_1_, DP_y_0_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10}) );
  ADD_TC_OP DP_add_216 ( .A({DP_pipe11[23], DP_pipe11[22], DP_pipe11[21], 
        DP_pipe11[20], DP_pipe11[19], DP_pipe11[18], DP_pipe11[17], 
        DP_pipe11[16], DP_pipe11[15], DP_pipe11[14], DP_pipe11[13], 
        DP_pipe11[12], DP_pipe11[11], DP_pipe11[10], DP_pipe11[9], 
        DP_pipe11[8], DP_pipe11[7], DP_pipe11[6], DP_pipe11[5], DP_pipe11[4], 
        DP_pipe11[3], DP_pipe11[2], DP_pipe11[1], DP_pipe11[0]}), .B({
        DP_ff_part[23], DP_ff_part[22], DP_ff_part[21], DP_ff_part[20], 
        DP_ff_part[19], DP_ff_part[18], DP_ff_part[17], DP_ff_part[16], 
        DP_ff_part[15], DP_ff_part[14], DP_ff_part[13], DP_ff_part[12], 
        DP_ff_part[11], DP_ff_part[10], DP_ff_part[9], DP_ff_part[8], 
        DP_ff_part[7], DP_ff_part[6], DP_ff_part[5], DP_ff_part[4], 
        DP_ff_part[3], DP_ff_part[2], DP_ff_part[1], DP_ff_part[0]}), .Z({
        DP_ff[23], DP_ff[22], DP_ff[21], DP_ff[20], DP_ff[19], DP_ff[18], 
        DP_ff[17], DP_ff[16], DP_ff[15], DP_ff[14], DP_ff[13], DP_ff[12], 
        DP_ff[11], DP_ff[10], DP_ff[9], DP_ff[8], DP_ff[7], DP_ff[6], DP_ff[5], 
        DP_ff[4], DP_ff[3], DP_ff[2], DP_ff[1], DP_ff[0]}) );
  SUB_TC_OP DP_sub_217 ( .A({DP_x[11], DP_x[10], DP_x[9], DP_x[8], DP_x[7], 
        DP_x[6], DP_x[5], DP_x[4], DP_x[3], DP_x[2], DP_x[1], DP_x[0], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        DP_fb[23], DP_fb[22], DP_fb[21], DP_fb[20], DP_fb[19], DP_fb[18], 
        DP_fb[17], DP_fb[16], DP_fb[15], DP_fb[14], DP_fb[13], DP_fb[12], 
        DP_fb[11], DP_fb[10], DP_fb[9], DP_fb[8], DP_fb[7], DP_fb[6], DP_fb[5], 
        DP_fb[4], DP_fb[3], DP_fb[2], DP_fb[1], DP_fb[0]}), .Z({DP_w_23_, 
        DP_w_22_, DP_w_21_, DP_w_20_, DP_w_19_, DP_w_18_, DP_w_17_, DP_w_16_, 
        DP_w_15_, DP_w_14_, DP_w_13_, DP_w_12_, DP_w_11_, DP_w_10_, DP_w_9_, 
        DP_w_8_, DP_w_7_, DP_w_6_, DP_w_5_, DP_w_4_, DP_w_3_, DP_w_2_, DP_w_1_, 
        DP_w_0_}) );
  ADD_TC_OP DP_add_215 ( .A({DP_pipe12[23], DP_pipe12[22], DP_pipe12[21], 
        DP_pipe12[20], DP_pipe12[19], DP_pipe12[18], DP_pipe12[17], 
        DP_pipe12[16], DP_pipe12[15], DP_pipe12[14], DP_pipe12[13], 
        DP_pipe12[12], DP_pipe12[11], DP_pipe12[10], DP_pipe12[9], 
        DP_pipe12[8], DP_pipe12[7], DP_pipe12[6], DP_pipe12[5], DP_pipe12[4], 
        DP_pipe12[3], DP_pipe12[2], DP_pipe12[1], DP_pipe12[0]}), .B({
        DP_pipe13[23], DP_pipe13[22], DP_pipe13[21], DP_pipe13[20], 
        DP_pipe13[19], DP_pipe13[18], DP_pipe13[17], DP_pipe13[16], 
        DP_pipe13[15], DP_pipe13[14], DP_pipe13[13], DP_pipe13[12], 
        DP_pipe13[11], DP_pipe13[10], DP_pipe13[9], DP_pipe13[8], DP_pipe13[7], 
        DP_pipe13[6], DP_pipe13[5], DP_pipe13[4], DP_pipe13[3], DP_pipe13[2], 
        DP_pipe13[1], DP_pipe13[0]}), .Z({DP_ff_part[23], DP_ff_part[22], 
        DP_ff_part[21], DP_ff_part[20], DP_ff_part[19], DP_ff_part[18], 
        DP_ff_part[17], DP_ff_part[16], DP_ff_part[15], DP_ff_part[14], 
        DP_ff_part[13], DP_ff_part[12], DP_ff_part[11], DP_ff_part[10], 
        DP_ff_part[9], DP_ff_part[8], DP_ff_part[7], DP_ff_part[6], 
        DP_ff_part[5], DP_ff_part[4], DP_ff_part[3], DP_ff_part[2], 
        DP_ff_part[1], DP_ff_part[0]}) );
  LT_TC_OP DP_lt_228 ( .A({DP_y_23, DP_y_23, DP_y_23, DP_y_23, DP_y_23, 
        DP_y_23, DP_y_23, DP_y_23, DP_y_23, DP_y_23, DP_y_23, DP_y_23, 
        DP_y_11_, DP_y_10_, DP_y_9_, DP_y_8_, DP_y_7_, DP_y_6_, DP_y_5_, 
        DP_y_4_, DP_y_3_, DP_y_2_, DP_y_1_, DP_y_0_}), .B({1'b1, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Z(DP_N4) );
  GT_TC_OP DP_gt_226 ( .A({DP_y_23, DP_y_23, DP_y_23, DP_y_23, DP_y_23, 
        DP_y_23, DP_y_23, DP_y_23, DP_y_23, DP_y_23, DP_y_23, DP_y_23, 
        DP_y_11_, DP_y_10_, DP_y_9_, DP_y_8_, DP_y_7_, DP_y_6_, DP_y_5_, 
        DP_y_4_, DP_y_3_, DP_y_2_, DP_y_1_, DP_y_0_}), .B({1'b0, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .Z(DP_N2) );
  ADD_TC_OP DP_add_214 ( .A({DP_ret0[23], DP_ret0[22], DP_ret0[21], 
        DP_ret0[20], DP_ret0[19], DP_ret0[18], DP_ret0[17], DP_ret0[16], 
        DP_ret0[15], DP_ret0[14], DP_ret0[13], DP_ret0[12], DP_ret0[11], 
        DP_ret0[10], DP_ret0[9], DP_ret0[8], DP_ret0[7], DP_ret0[6], 
        DP_ret0[5], DP_ret0[4], DP_ret0[3], DP_ret0[2], DP_ret0[1], DP_ret0[0]}), .B({DP_ret1[23], DP_ret1[22], DP_ret1[21], DP_ret1[20], DP_ret1[19], 
        DP_ret1[18], DP_ret1[17], DP_ret1[16], DP_ret1[15], DP_ret1[14], 
        DP_ret1[13], DP_ret1[12], DP_ret1[11], DP_ret1[10], DP_ret1[9], 
        DP_ret1[8], DP_ret1[7], DP_ret1[6], DP_ret1[5], DP_ret1[4], DP_ret1[3], 
        DP_ret1[2], DP_ret1[1], DP_ret1[0]}), .Z({DP_fb[23], DP_fb[22], 
        DP_fb[21], DP_fb[20], DP_fb[19], DP_fb[18], DP_fb[17], DP_fb[16], 
        DP_fb[15], DP_fb[14], DP_fb[13], DP_fb[12], DP_fb[11], DP_fb[10], 
        DP_fb[9], DP_fb[8], DP_fb[7], DP_fb[6], DP_fb[5], DP_fb[4], DP_fb[3], 
        DP_fb[2], DP_fb[1], DP_fb[0]}) );
  MULT_TC_OP DP_mult_209 ( .A({DP_coeffs_ff_int[72], DP_coeffs_ff_int[73], 
        DP_coeffs_ff_int[74], DP_coeffs_ff_int[75], DP_coeffs_ff_int[76], 
        DP_coeffs_ff_int[77], DP_coeffs_ff_int[78], DP_coeffs_ff_int[79], 
        DP_coeffs_ff_int[80], DP_coeffs_ff_int[81], DP_coeffs_ff_int[82], 
        DP_coeffs_ff_int[83], DP_coeffs_ff_int[84], DP_coeffs_ff_int[85], 
        DP_coeffs_ff_int[86], DP_coeffs_ff_int[87], DP_coeffs_ff_int[88], 
        DP_coeffs_ff_int[89], DP_coeffs_ff_int[90], DP_coeffs_ff_int[91], 
        DP_coeffs_ff_int[92], DP_coeffs_ff_int[93], DP_coeffs_ff_int[94], 
        DP_coeffs_ff_int[95]}), .B({DP_pipe03[23], DP_pipe03[22], 
        DP_pipe03[21], DP_pipe03[20], DP_pipe03[19], DP_pipe03[18], 
        DP_pipe03[17], DP_pipe03[16], DP_pipe03[15], DP_pipe03[14], 
        DP_pipe03[13], DP_pipe03[12], DP_pipe03[11], DP_pipe03[10], 
        DP_pipe03[9], DP_pipe03[8], DP_pipe03[7], DP_pipe03[6], DP_pipe03[5], 
        DP_pipe03[4], DP_pipe03[3], DP_pipe03[2], DP_pipe03[1], DP_pipe03[0]}), 
        .Z({DP_pipe0_coeff_pipe03[23], SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, DP_pipe0_coeff_pipe03[22], 
        DP_pipe0_coeff_pipe03[21], DP_pipe0_coeff_pipe03[20], 
        DP_pipe0_coeff_pipe03[19], DP_pipe0_coeff_pipe03[18], 
        DP_pipe0_coeff_pipe03[17], DP_pipe0_coeff_pipe03[16], 
        DP_pipe0_coeff_pipe03[15], DP_pipe0_coeff_pipe03[14], 
        DP_pipe0_coeff_pipe03[13], DP_pipe0_coeff_pipe03[12], 
        DP_pipe0_coeff_pipe03[11], DP_pipe0_coeff_pipe03[10], 
        DP_pipe0_coeff_pipe03[9], DP_pipe0_coeff_pipe03[8], 
        DP_pipe0_coeff_pipe03[7], DP_pipe0_coeff_pipe03[6], 
        DP_pipe0_coeff_pipe03[5], DP_pipe0_coeff_pipe03[4], 
        DP_pipe0_coeff_pipe03[3], DP_pipe0_coeff_pipe03[2], 
        DP_pipe0_coeff_pipe03[1], DP_pipe0_coeff_pipe03[0], 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34}) );
  MULT_TC_OP DP_mult_208 ( .A({DP_coeffs_ff_int[48], DP_coeffs_ff_int[49], 
        DP_coeffs_ff_int[50], DP_coeffs_ff_int[51], DP_coeffs_ff_int[52], 
        DP_coeffs_ff_int[53], DP_coeffs_ff_int[54], DP_coeffs_ff_int[55], 
        DP_coeffs_ff_int[56], DP_coeffs_ff_int[57], DP_coeffs_ff_int[58], 
        DP_coeffs_ff_int[59], DP_coeffs_ff_int[60], DP_coeffs_ff_int[61], 
        DP_coeffs_ff_int[62], DP_coeffs_ff_int[63], DP_coeffs_ff_int[64], 
        DP_coeffs_ff_int[65], DP_coeffs_ff_int[66], DP_coeffs_ff_int[67], 
        DP_coeffs_ff_int[68], DP_coeffs_ff_int[69], DP_coeffs_ff_int[70], 
        DP_coeffs_ff_int[71]}), .B({DP_pipe02[23], DP_pipe02[22], 
        DP_pipe02[21], DP_pipe02[20], DP_pipe02[19], DP_pipe02[18], 
        DP_pipe02[17], DP_pipe02[16], DP_pipe02[15], DP_pipe02[14], 
        DP_pipe02[13], DP_pipe02[12], DP_pipe02[11], DP_pipe02[10], 
        DP_pipe02[9], DP_pipe02[8], DP_pipe02[7], DP_pipe02[6], DP_pipe02[5], 
        DP_pipe02[4], DP_pipe02[3], DP_pipe02[2], DP_pipe02[1], DP_pipe02[0]}), 
        .Z({DP_pipe0_coeff_pipe02[23], SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, DP_pipe0_coeff_pipe02[22], 
        DP_pipe0_coeff_pipe02[21], DP_pipe0_coeff_pipe02[20], 
        DP_pipe0_coeff_pipe02[19], DP_pipe0_coeff_pipe02[18], 
        DP_pipe0_coeff_pipe02[17], DP_pipe0_coeff_pipe02[16], 
        DP_pipe0_coeff_pipe02[15], DP_pipe0_coeff_pipe02[14], 
        DP_pipe0_coeff_pipe02[13], DP_pipe0_coeff_pipe02[12], 
        DP_pipe0_coeff_pipe02[11], DP_pipe0_coeff_pipe02[10], 
        DP_pipe0_coeff_pipe02[9], DP_pipe0_coeff_pipe02[8], 
        DP_pipe0_coeff_pipe02[7], DP_pipe0_coeff_pipe02[6], 
        DP_pipe0_coeff_pipe02[5], DP_pipe0_coeff_pipe02[4], 
        DP_pipe0_coeff_pipe02[3], DP_pipe0_coeff_pipe02[2], 
        DP_pipe0_coeff_pipe02[1], DP_pipe0_coeff_pipe02[0], 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, 
        SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48, 
        SYNOPSYS_UNCONNECTED__49, SYNOPSYS_UNCONNECTED__50, 
        SYNOPSYS_UNCONNECTED__51, SYNOPSYS_UNCONNECTED__52, 
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54, 
        SYNOPSYS_UNCONNECTED__55, SYNOPSYS_UNCONNECTED__56, 
        SYNOPSYS_UNCONNECTED__57, SYNOPSYS_UNCONNECTED__58}) );
  MULT_TC_OP DP_mult_207 ( .A({DP_coeffs_ff_int[24], DP_coeffs_ff_int[25], 
        DP_coeffs_ff_int[26], DP_coeffs_ff_int[27], DP_coeffs_ff_int[28], 
        DP_coeffs_ff_int[29], DP_coeffs_ff_int[30], DP_coeffs_ff_int[31], 
        DP_coeffs_ff_int[32], DP_coeffs_ff_int[33], DP_coeffs_ff_int[34], 
        DP_coeffs_ff_int[35], DP_coeffs_ff_int[36], DP_coeffs_ff_int[37], 
        DP_coeffs_ff_int[38], DP_coeffs_ff_int[39], DP_coeffs_ff_int[40], 
        DP_coeffs_ff_int[41], DP_coeffs_ff_int[42], DP_coeffs_ff_int[43], 
        DP_coeffs_ff_int[44], DP_coeffs_ff_int[45], DP_coeffs_ff_int[46], 
        DP_coeffs_ff_int[47]}), .B({DP_pipe01[23], DP_pipe01[22], 
        DP_pipe01[21], DP_pipe01[20], DP_pipe01[19], DP_pipe01[18], 
        DP_pipe01[17], DP_pipe01[16], DP_pipe01[15], DP_pipe01[14], 
        DP_pipe01[13], DP_pipe01[12], DP_pipe01[11], DP_pipe01[10], 
        DP_pipe01[9], DP_pipe01[8], DP_pipe01[7], DP_pipe01[6], DP_pipe01[5], 
        DP_pipe01[4], DP_pipe01[3], DP_pipe01[2], DP_pipe01[1], DP_pipe01[0]}), 
        .Z({DP_pipe0_coeff_pipe01[23], SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, DP_pipe0_coeff_pipe01[22], 
        DP_pipe0_coeff_pipe01[21], DP_pipe0_coeff_pipe01[20], 
        DP_pipe0_coeff_pipe01[19], DP_pipe0_coeff_pipe01[18], 
        DP_pipe0_coeff_pipe01[17], DP_pipe0_coeff_pipe01[16], 
        DP_pipe0_coeff_pipe01[15], DP_pipe0_coeff_pipe01[14], 
        DP_pipe0_coeff_pipe01[13], DP_pipe0_coeff_pipe01[12], 
        DP_pipe0_coeff_pipe01[11], DP_pipe0_coeff_pipe01[10], 
        DP_pipe0_coeff_pipe01[9], DP_pipe0_coeff_pipe01[8], 
        DP_pipe0_coeff_pipe01[7], DP_pipe0_coeff_pipe01[6], 
        DP_pipe0_coeff_pipe01[5], DP_pipe0_coeff_pipe01[4], 
        DP_pipe0_coeff_pipe01[3], DP_pipe0_coeff_pipe01[2], 
        DP_pipe0_coeff_pipe01[1], DP_pipe0_coeff_pipe01[0], 
        SYNOPSYS_UNCONNECTED__61, SYNOPSYS_UNCONNECTED__62, 
        SYNOPSYS_UNCONNECTED__63, SYNOPSYS_UNCONNECTED__64, 
        SYNOPSYS_UNCONNECTED__65, SYNOPSYS_UNCONNECTED__66, 
        SYNOPSYS_UNCONNECTED__67, SYNOPSYS_UNCONNECTED__68, 
        SYNOPSYS_UNCONNECTED__69, SYNOPSYS_UNCONNECTED__70, 
        SYNOPSYS_UNCONNECTED__71, SYNOPSYS_UNCONNECTED__72, 
        SYNOPSYS_UNCONNECTED__73, SYNOPSYS_UNCONNECTED__74, 
        SYNOPSYS_UNCONNECTED__75, SYNOPSYS_UNCONNECTED__76, 
        SYNOPSYS_UNCONNECTED__77, SYNOPSYS_UNCONNECTED__78, 
        SYNOPSYS_UNCONNECTED__79, SYNOPSYS_UNCONNECTED__80, 
        SYNOPSYS_UNCONNECTED__81, SYNOPSYS_UNCONNECTED__82}) );
  MULT_TC_OP DP_mult_206 ( .A({DP_coeffs_ff_int[0], DP_coeffs_ff_int[1], 
        DP_coeffs_ff_int[2], DP_coeffs_ff_int[3], DP_coeffs_ff_int[4], 
        DP_coeffs_ff_int[5], DP_coeffs_ff_int[6], DP_coeffs_ff_int[7], 
        DP_coeffs_ff_int[8], DP_coeffs_ff_int[9], DP_coeffs_ff_int[10], 
        DP_coeffs_ff_int[11], DP_coeffs_ff_int[12], DP_coeffs_ff_int[13], 
        DP_coeffs_ff_int[14], DP_coeffs_ff_int[15], DP_coeffs_ff_int[16], 
        DP_coeffs_ff_int[17], DP_coeffs_ff_int[18], DP_coeffs_ff_int[19], 
        DP_coeffs_ff_int[20], DP_coeffs_ff_int[21], DP_coeffs_ff_int[22], 
        DP_coeffs_ff_int[23]}), .B({DP_pipe00[23], DP_pipe00[22], 
        DP_pipe00[21], DP_pipe00[20], DP_pipe00[19], DP_pipe00[18], 
        DP_pipe00[17], DP_pipe00[16], DP_pipe00[15], DP_pipe00[14], 
        DP_pipe00[13], DP_pipe00[12], DP_pipe00[11], DP_pipe00[10], 
        DP_pipe00[9], DP_pipe00[8], DP_pipe00[7], DP_pipe00[6], DP_pipe00[5], 
        DP_pipe00[4], DP_pipe00[3], DP_pipe00[2], DP_pipe00[1], DP_pipe00[0]}), 
        .Z({DP_pipe0_coeff_pipe00[23], SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, DP_pipe0_coeff_pipe00[22], 
        DP_pipe0_coeff_pipe00[21], DP_pipe0_coeff_pipe00[20], 
        DP_pipe0_coeff_pipe00[19], DP_pipe0_coeff_pipe00[18], 
        DP_pipe0_coeff_pipe00[17], DP_pipe0_coeff_pipe00[16], 
        DP_pipe0_coeff_pipe00[15], DP_pipe0_coeff_pipe00[14], 
        DP_pipe0_coeff_pipe00[13], DP_pipe0_coeff_pipe00[12], 
        DP_pipe0_coeff_pipe00[11], DP_pipe0_coeff_pipe00[10], 
        DP_pipe0_coeff_pipe00[9], DP_pipe0_coeff_pipe00[8], 
        DP_pipe0_coeff_pipe00[7], DP_pipe0_coeff_pipe00[6], 
        DP_pipe0_coeff_pipe00[5], DP_pipe0_coeff_pipe00[4], 
        DP_pipe0_coeff_pipe00[3], DP_pipe0_coeff_pipe00[2], 
        DP_pipe0_coeff_pipe00[1], DP_pipe0_coeff_pipe00[0], 
        SYNOPSYS_UNCONNECTED__85, SYNOPSYS_UNCONNECTED__86, 
        SYNOPSYS_UNCONNECTED__87, SYNOPSYS_UNCONNECTED__88, 
        SYNOPSYS_UNCONNECTED__89, SYNOPSYS_UNCONNECTED__90, 
        SYNOPSYS_UNCONNECTED__91, SYNOPSYS_UNCONNECTED__92, 
        SYNOPSYS_UNCONNECTED__93, SYNOPSYS_UNCONNECTED__94, 
        SYNOPSYS_UNCONNECTED__95, SYNOPSYS_UNCONNECTED__96, 
        SYNOPSYS_UNCONNECTED__97, SYNOPSYS_UNCONNECTED__98, 
        SYNOPSYS_UNCONNECTED__99, SYNOPSYS_UNCONNECTED__100, 
        SYNOPSYS_UNCONNECTED__101, SYNOPSYS_UNCONNECTED__102, 
        SYNOPSYS_UNCONNECTED__103, SYNOPSYS_UNCONNECTED__104, 
        SYNOPSYS_UNCONNECTED__105, SYNOPSYS_UNCONNECTED__106}) );
  MULT_TC_OP DP_mult_205 ( .A({DP_coeffs_fb_int[24], DP_coeffs_fb_int[25], 
        DP_coeffs_fb_int[26], DP_coeffs_fb_int[27], DP_coeffs_fb_int[28], 
        DP_coeffs_fb_int[29], DP_coeffs_fb_int[30], DP_coeffs_fb_int[31], 
        DP_coeffs_fb_int[32], DP_coeffs_fb_int[33], DP_coeffs_fb_int[34], 
        DP_coeffs_fb_int[35], DP_coeffs_fb_int[36], DP_coeffs_fb_int[37], 
        DP_coeffs_fb_int[38], DP_coeffs_fb_int[39], DP_coeffs_fb_int[40], 
        DP_coeffs_fb_int[41], DP_coeffs_fb_int[42], DP_coeffs_fb_int[43], 
        DP_coeffs_fb_int[44], DP_coeffs_fb_int[45], DP_coeffs_fb_int[46], 
        DP_coeffs_fb_int[47]}), .B({DP_sw1_23_, DP_sw1_22_, DP_sw1_21_, 
        DP_sw1_20_, DP_sw1_19_, DP_sw1_18_, DP_sw1_17_, DP_sw1_16_, DP_sw1_15_, 
        DP_sw1_14_, DP_sw1_13_, DP_sw1_12_, DP_sw1_11_, DP_sw1_10_, DP_sw1_9_, 
        DP_sw1_8_, DP_sw1_7_, DP_sw1_6_, DP_sw1_5_, DP_sw1_4_, DP_sw1_3_, 
        DP_sw1_2_, DP_sw1_1_, DP_sw1_0_}), .Z({DP_sw1_coeff_ret1[23], 
        SYNOPSYS_UNCONNECTED__107, SYNOPSYS_UNCONNECTED__108, 
        DP_sw1_coeff_ret1[22], DP_sw1_coeff_ret1[21], DP_sw1_coeff_ret1[20], 
        DP_sw1_coeff_ret1[19], DP_sw1_coeff_ret1[18], DP_sw1_coeff_ret1[17], 
        DP_sw1_coeff_ret1[16], DP_sw1_coeff_ret1[15], DP_sw1_coeff_ret1[14], 
        DP_sw1_coeff_ret1[13], DP_sw1_coeff_ret1[12], DP_sw1_coeff_ret1[11], 
        DP_sw1_coeff_ret1[10], DP_sw1_coeff_ret1[9], DP_sw1_coeff_ret1[8], 
        DP_sw1_coeff_ret1[7], DP_sw1_coeff_ret1[6], DP_sw1_coeff_ret1[5], 
        DP_sw1_coeff_ret1[4], DP_sw1_coeff_ret1[3], DP_sw1_coeff_ret1[2], 
        DP_sw1_coeff_ret1[1], DP_sw1_coeff_ret1[0], SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130}) );
  MULT_TC_OP DP_mult_204 ( .A({DP_coeffs_fb_int[0], DP_coeffs_fb_int[1], 
        DP_coeffs_fb_int[2], DP_coeffs_fb_int[3], DP_coeffs_fb_int[4], 
        DP_coeffs_fb_int[5], DP_coeffs_fb_int[6], DP_coeffs_fb_int[7], 
        DP_coeffs_fb_int[8], DP_coeffs_fb_int[9], DP_coeffs_fb_int[10], 
        DP_coeffs_fb_int[11], DP_coeffs_fb_int[12], DP_coeffs_fb_int[13], 
        DP_coeffs_fb_int[14], DP_coeffs_fb_int[15], DP_coeffs_fb_int[16], 
        DP_coeffs_fb_int[17], DP_coeffs_fb_int[18], DP_coeffs_fb_int[19], 
        DP_coeffs_fb_int[20], DP_coeffs_fb_int[21], DP_coeffs_fb_int[22], 
        DP_coeffs_fb_int[23]}), .B({DP_sw0_23_, DP_sw0_22_, DP_sw0_21_, 
        DP_sw0_20_, DP_sw0_19_, DP_sw0_18_, DP_sw0_17_, DP_sw0_16_, DP_sw0_15_, 
        DP_sw0_14_, DP_sw0_13_, DP_sw0_12_, DP_sw0_11_, DP_sw0_10_, DP_sw0_9_, 
        DP_sw0_8_, DP_sw0_7_, DP_sw0_6_, DP_sw0_5_, DP_sw0_4_, DP_sw0_3_, 
        DP_sw0_2_, DP_sw0_1_, DP_sw0_0_}), .Z({DP_sw0_coeff_ret0[23], 
        SYNOPSYS_UNCONNECTED__131, SYNOPSYS_UNCONNECTED__132, 
        DP_sw0_coeff_ret0[22], DP_sw0_coeff_ret0[21], DP_sw0_coeff_ret0[20], 
        DP_sw0_coeff_ret0[19], DP_sw0_coeff_ret0[18], DP_sw0_coeff_ret0[17], 
        DP_sw0_coeff_ret0[16], DP_sw0_coeff_ret0[15], DP_sw0_coeff_ret0[14], 
        DP_sw0_coeff_ret0[13], DP_sw0_coeff_ret0[12], DP_sw0_coeff_ret0[11], 
        DP_sw0_coeff_ret0[10], DP_sw0_coeff_ret0[9], DP_sw0_coeff_ret0[8], 
        DP_sw0_coeff_ret0[7], DP_sw0_coeff_ret0[6], DP_sw0_coeff_ret0[5], 
        DP_sw0_coeff_ret0[4], DP_sw0_coeff_ret0[3], DP_sw0_coeff_ret0[2], 
        DP_sw0_coeff_ret0[1], DP_sw0_coeff_ret0[0], SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154}) );
  GTECH_NOT DP_reg_in_I_0 ( .A(rst_n), .Z(DP_reg_in_N0) );
  \**SEQGEN**  DP_reg_in_Q_reg_0_ ( .clear(DP_reg_in_N0), .preset(1'b0), 
        .next_state(dIn[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_x[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_in_Q_reg_1_ ( .clear(DP_reg_in_N0), .preset(1'b0), 
        .next_state(dIn[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_x[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_in_Q_reg_2_ ( .clear(DP_reg_in_N0), .preset(1'b0), 
        .next_state(dIn[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_x[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_in_Q_reg_3_ ( .clear(DP_reg_in_N0), .preset(1'b0), 
        .next_state(dIn[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_x[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_in_Q_reg_4_ ( .clear(DP_reg_in_N0), .preset(1'b0), 
        .next_state(dIn[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_x[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_in_Q_reg_5_ ( .clear(DP_reg_in_N0), .preset(1'b0), 
        .next_state(dIn[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_x[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_in_Q_reg_6_ ( .clear(DP_reg_in_N0), .preset(1'b0), 
        .next_state(dIn[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_x[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_in_Q_reg_7_ ( .clear(DP_reg_in_N0), .preset(1'b0), 
        .next_state(dIn[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_x[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_in_Q_reg_8_ ( .clear(DP_reg_in_N0), .preset(1'b0), 
        .next_state(dIn[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_x[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_in_Q_reg_9_ ( .clear(DP_reg_in_N0), .preset(1'b0), 
        .next_state(dIn[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_x[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_in_Q_reg_10_ ( .clear(DP_reg_in_N0), .preset(1'b0), 
        .next_state(dIn[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_x[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_in_Q_reg_11_ ( .clear(DP_reg_in_N0), .preset(1'b0), 
        .next_state(dIn[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_x[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(vIn) );
  GTECH_NOT DP_reg_coeff_fb_i_1_I_0 ( .A(rst_n), .Z(DP_reg_coeff_fb_i_1_N0) );
  \**SEQGEN**  DP_reg_coeff_fb_i_1_Q_reg_0_ ( .clear(DP_reg_coeff_fb_i_1_N0), 
        .preset(1'b0), .next_state(coeffs_fb[24]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[23]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_1_Q_reg_1_ ( .clear(DP_reg_coeff_fb_i_1_N0), 
        .preset(1'b0), .next_state(coeffs_fb[25]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[22]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_1_Q_reg_2_ ( .clear(DP_reg_coeff_fb_i_1_N0), 
        .preset(1'b0), .next_state(coeffs_fb[26]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[21]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_1_Q_reg_3_ ( .clear(DP_reg_coeff_fb_i_1_N0), 
        .preset(1'b0), .next_state(coeffs_fb[27]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[20]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_1_Q_reg_4_ ( .clear(DP_reg_coeff_fb_i_1_N0), 
        .preset(1'b0), .next_state(coeffs_fb[28]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[19]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_1_Q_reg_5_ ( .clear(DP_reg_coeff_fb_i_1_N0), 
        .preset(1'b0), .next_state(coeffs_fb[29]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[18]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_1_Q_reg_6_ ( .clear(DP_reg_coeff_fb_i_1_N0), 
        .preset(1'b0), .next_state(coeffs_fb[30]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[17]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_1_Q_reg_7_ ( .clear(DP_reg_coeff_fb_i_1_N0), 
        .preset(1'b0), .next_state(coeffs_fb[31]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[16]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_1_Q_reg_8_ ( .clear(DP_reg_coeff_fb_i_1_N0), 
        .preset(1'b0), .next_state(coeffs_fb[32]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[15]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_1_Q_reg_9_ ( .clear(DP_reg_coeff_fb_i_1_N0), 
        .preset(1'b0), .next_state(coeffs_fb[33]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[14]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_1_Q_reg_10_ ( .clear(DP_reg_coeff_fb_i_1_N0), 
        .preset(1'b0), .next_state(coeffs_fb[34]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[13]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_1_Q_reg_11_ ( .clear(DP_reg_coeff_fb_i_1_N0), 
        .preset(1'b0), .next_state(coeffs_fb[35]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[12]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_1_Q_reg_12_ ( .clear(DP_reg_coeff_fb_i_1_N0), 
        .preset(1'b0), .next_state(coeffs_fb[36]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[11]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_1_Q_reg_13_ ( .clear(DP_reg_coeff_fb_i_1_N0), 
        .preset(1'b0), .next_state(coeffs_fb[37]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[10]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_1_Q_reg_14_ ( .clear(DP_reg_coeff_fb_i_1_N0), 
        .preset(1'b0), .next_state(coeffs_fb[38]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[9]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_1_Q_reg_15_ ( .clear(DP_reg_coeff_fb_i_1_N0), 
        .preset(1'b0), .next_state(coeffs_fb[39]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[8]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_1_Q_reg_16_ ( .clear(DP_reg_coeff_fb_i_1_N0), 
        .preset(1'b0), .next_state(coeffs_fb[40]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[7]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_1_Q_reg_17_ ( .clear(DP_reg_coeff_fb_i_1_N0), 
        .preset(1'b0), .next_state(coeffs_fb[41]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[6]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_1_Q_reg_18_ ( .clear(DP_reg_coeff_fb_i_1_N0), 
        .preset(1'b0), .next_state(coeffs_fb[42]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[5]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_1_Q_reg_19_ ( .clear(DP_reg_coeff_fb_i_1_N0), 
        .preset(1'b0), .next_state(coeffs_fb[43]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[4]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_1_Q_reg_20_ ( .clear(DP_reg_coeff_fb_i_1_N0), 
        .preset(1'b0), .next_state(coeffs_fb[44]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[3]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_1_Q_reg_21_ ( .clear(DP_reg_coeff_fb_i_1_N0), 
        .preset(1'b0), .next_state(coeffs_fb[45]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[2]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_1_Q_reg_22_ ( .clear(DP_reg_coeff_fb_i_1_N0), 
        .preset(1'b0), .next_state(coeffs_fb[46]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[1]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_1_Q_reg_23_ ( .clear(DP_reg_coeff_fb_i_1_N0), 
        .preset(1'b0), .next_state(coeffs_fb[47]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[0]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  GTECH_NOT DP_reg_coeff_fb_i_2_I_0 ( .A(rst_n), .Z(DP_reg_coeff_fb_i_2_N0) );
  \**SEQGEN**  DP_reg_coeff_fb_i_2_Q_reg_0_ ( .clear(DP_reg_coeff_fb_i_2_N0), 
        .preset(1'b0), .next_state(coeffs_fb[0]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[47]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_2_Q_reg_1_ ( .clear(DP_reg_coeff_fb_i_2_N0), 
        .preset(1'b0), .next_state(coeffs_fb[1]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[46]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_2_Q_reg_2_ ( .clear(DP_reg_coeff_fb_i_2_N0), 
        .preset(1'b0), .next_state(coeffs_fb[2]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[45]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_2_Q_reg_3_ ( .clear(DP_reg_coeff_fb_i_2_N0), 
        .preset(1'b0), .next_state(coeffs_fb[3]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[44]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_2_Q_reg_4_ ( .clear(DP_reg_coeff_fb_i_2_N0), 
        .preset(1'b0), .next_state(coeffs_fb[4]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[43]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_2_Q_reg_5_ ( .clear(DP_reg_coeff_fb_i_2_N0), 
        .preset(1'b0), .next_state(coeffs_fb[5]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[42]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_2_Q_reg_6_ ( .clear(DP_reg_coeff_fb_i_2_N0), 
        .preset(1'b0), .next_state(coeffs_fb[6]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[41]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_2_Q_reg_7_ ( .clear(DP_reg_coeff_fb_i_2_N0), 
        .preset(1'b0), .next_state(coeffs_fb[7]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[40]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_2_Q_reg_8_ ( .clear(DP_reg_coeff_fb_i_2_N0), 
        .preset(1'b0), .next_state(coeffs_fb[8]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[39]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_2_Q_reg_9_ ( .clear(DP_reg_coeff_fb_i_2_N0), 
        .preset(1'b0), .next_state(coeffs_fb[9]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[38]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_2_Q_reg_10_ ( .clear(DP_reg_coeff_fb_i_2_N0), 
        .preset(1'b0), .next_state(coeffs_fb[10]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[37]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_2_Q_reg_11_ ( .clear(DP_reg_coeff_fb_i_2_N0), 
        .preset(1'b0), .next_state(coeffs_fb[11]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[36]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_2_Q_reg_12_ ( .clear(DP_reg_coeff_fb_i_2_N0), 
        .preset(1'b0), .next_state(coeffs_fb[12]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[35]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_2_Q_reg_13_ ( .clear(DP_reg_coeff_fb_i_2_N0), 
        .preset(1'b0), .next_state(coeffs_fb[13]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[34]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_2_Q_reg_14_ ( .clear(DP_reg_coeff_fb_i_2_N0), 
        .preset(1'b0), .next_state(coeffs_fb[14]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[33]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_2_Q_reg_15_ ( .clear(DP_reg_coeff_fb_i_2_N0), 
        .preset(1'b0), .next_state(coeffs_fb[15]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[32]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_2_Q_reg_16_ ( .clear(DP_reg_coeff_fb_i_2_N0), 
        .preset(1'b0), .next_state(coeffs_fb[16]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[31]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_2_Q_reg_17_ ( .clear(DP_reg_coeff_fb_i_2_N0), 
        .preset(1'b0), .next_state(coeffs_fb[17]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[30]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_2_Q_reg_18_ ( .clear(DP_reg_coeff_fb_i_2_N0), 
        .preset(1'b0), .next_state(coeffs_fb[18]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[29]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_2_Q_reg_19_ ( .clear(DP_reg_coeff_fb_i_2_N0), 
        .preset(1'b0), .next_state(coeffs_fb[19]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[28]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_2_Q_reg_20_ ( .clear(DP_reg_coeff_fb_i_2_N0), 
        .preset(1'b0), .next_state(coeffs_fb[20]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[27]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_2_Q_reg_21_ ( .clear(DP_reg_coeff_fb_i_2_N0), 
        .preset(1'b0), .next_state(coeffs_fb[21]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[26]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_2_Q_reg_22_ ( .clear(DP_reg_coeff_fb_i_2_N0), 
        .preset(1'b0), .next_state(coeffs_fb[22]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[25]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_coeff_fb_i_2_Q_reg_23_ ( .clear(DP_reg_coeff_fb_i_2_N0), 
        .preset(1'b0), .next_state(coeffs_fb[23]), .clocked_on(clk), .data_in(
        1'b0), .enable(1'b0), .Q(DP_coeffs_fb_int[24]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  GTECH_NOT DP_reg_b_i_0_I_0 ( .A(rst_n), .Z(DP_reg_b_i_0_N0) );
  \**SEQGEN**  DP_reg_b_i_0_Q_reg_0_ ( .clear(DP_reg_b_i_0_N0), .preset(1'b0), 
        .next_state(coeffs_ff[72]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[23]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_0_Q_reg_1_ ( .clear(DP_reg_b_i_0_N0), .preset(1'b0), 
        .next_state(coeffs_ff[73]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[22]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_0_Q_reg_2_ ( .clear(DP_reg_b_i_0_N0), .preset(1'b0), 
        .next_state(coeffs_ff[74]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[21]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_0_Q_reg_3_ ( .clear(DP_reg_b_i_0_N0), .preset(1'b0), 
        .next_state(coeffs_ff[75]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[20]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_0_Q_reg_4_ ( .clear(DP_reg_b_i_0_N0), .preset(1'b0), 
        .next_state(coeffs_ff[76]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[19]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_0_Q_reg_5_ ( .clear(DP_reg_b_i_0_N0), .preset(1'b0), 
        .next_state(coeffs_ff[77]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[18]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_0_Q_reg_6_ ( .clear(DP_reg_b_i_0_N0), .preset(1'b0), 
        .next_state(coeffs_ff[78]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[17]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_0_Q_reg_7_ ( .clear(DP_reg_b_i_0_N0), .preset(1'b0), 
        .next_state(coeffs_ff[79]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[16]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_0_Q_reg_8_ ( .clear(DP_reg_b_i_0_N0), .preset(1'b0), 
        .next_state(coeffs_ff[80]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[15]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_0_Q_reg_9_ ( .clear(DP_reg_b_i_0_N0), .preset(1'b0), 
        .next_state(coeffs_ff[81]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[14]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_0_Q_reg_10_ ( .clear(DP_reg_b_i_0_N0), .preset(1'b0), 
        .next_state(coeffs_ff[82]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[13]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_0_Q_reg_11_ ( .clear(DP_reg_b_i_0_N0), .preset(1'b0), 
        .next_state(coeffs_ff[83]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[12]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_0_Q_reg_12_ ( .clear(DP_reg_b_i_0_N0), .preset(1'b0), 
        .next_state(coeffs_ff[84]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[11]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_0_Q_reg_13_ ( .clear(DP_reg_b_i_0_N0), .preset(1'b0), 
        .next_state(coeffs_ff[85]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[10]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_0_Q_reg_14_ ( .clear(DP_reg_b_i_0_N0), .preset(1'b0), 
        .next_state(coeffs_ff[86]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_0_Q_reg_15_ ( .clear(DP_reg_b_i_0_N0), .preset(1'b0), 
        .next_state(coeffs_ff[87]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_0_Q_reg_16_ ( .clear(DP_reg_b_i_0_N0), .preset(1'b0), 
        .next_state(coeffs_ff[88]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_0_Q_reg_17_ ( .clear(DP_reg_b_i_0_N0), .preset(1'b0), 
        .next_state(coeffs_ff[89]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_0_Q_reg_18_ ( .clear(DP_reg_b_i_0_N0), .preset(1'b0), 
        .next_state(coeffs_ff[90]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_0_Q_reg_19_ ( .clear(DP_reg_b_i_0_N0), .preset(1'b0), 
        .next_state(coeffs_ff[91]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_0_Q_reg_20_ ( .clear(DP_reg_b_i_0_N0), .preset(1'b0), 
        .next_state(coeffs_ff[92]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_0_Q_reg_21_ ( .clear(DP_reg_b_i_0_N0), .preset(1'b0), 
        .next_state(coeffs_ff[93]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_0_Q_reg_22_ ( .clear(DP_reg_b_i_0_N0), .preset(1'b0), 
        .next_state(coeffs_ff[94]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_0_Q_reg_23_ ( .clear(DP_reg_b_i_0_N0), .preset(1'b0), 
        .next_state(coeffs_ff[95]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  GTECH_NOT DP_reg_b_i_1_I_0 ( .A(rst_n), .Z(DP_reg_b_i_1_N0) );
  \**SEQGEN**  DP_reg_b_i_1_Q_reg_0_ ( .clear(DP_reg_b_i_1_N0), .preset(1'b0), 
        .next_state(coeffs_ff[48]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[47]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_1_Q_reg_1_ ( .clear(DP_reg_b_i_1_N0), .preset(1'b0), 
        .next_state(coeffs_ff[49]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[46]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_1_Q_reg_2_ ( .clear(DP_reg_b_i_1_N0), .preset(1'b0), 
        .next_state(coeffs_ff[50]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[45]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_1_Q_reg_3_ ( .clear(DP_reg_b_i_1_N0), .preset(1'b0), 
        .next_state(coeffs_ff[51]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[44]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_1_Q_reg_4_ ( .clear(DP_reg_b_i_1_N0), .preset(1'b0), 
        .next_state(coeffs_ff[52]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[43]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_1_Q_reg_5_ ( .clear(DP_reg_b_i_1_N0), .preset(1'b0), 
        .next_state(coeffs_ff[53]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[42]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_1_Q_reg_6_ ( .clear(DP_reg_b_i_1_N0), .preset(1'b0), 
        .next_state(coeffs_ff[54]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[41]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_1_Q_reg_7_ ( .clear(DP_reg_b_i_1_N0), .preset(1'b0), 
        .next_state(coeffs_ff[55]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[40]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_1_Q_reg_8_ ( .clear(DP_reg_b_i_1_N0), .preset(1'b0), 
        .next_state(coeffs_ff[56]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[39]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_1_Q_reg_9_ ( .clear(DP_reg_b_i_1_N0), .preset(1'b0), 
        .next_state(coeffs_ff[57]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[38]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_1_Q_reg_10_ ( .clear(DP_reg_b_i_1_N0), .preset(1'b0), 
        .next_state(coeffs_ff[58]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[37]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_1_Q_reg_11_ ( .clear(DP_reg_b_i_1_N0), .preset(1'b0), 
        .next_state(coeffs_ff[59]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[36]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_1_Q_reg_12_ ( .clear(DP_reg_b_i_1_N0), .preset(1'b0), 
        .next_state(coeffs_ff[60]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[35]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_1_Q_reg_13_ ( .clear(DP_reg_b_i_1_N0), .preset(1'b0), 
        .next_state(coeffs_ff[61]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[34]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_1_Q_reg_14_ ( .clear(DP_reg_b_i_1_N0), .preset(1'b0), 
        .next_state(coeffs_ff[62]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[33]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_1_Q_reg_15_ ( .clear(DP_reg_b_i_1_N0), .preset(1'b0), 
        .next_state(coeffs_ff[63]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[32]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_1_Q_reg_16_ ( .clear(DP_reg_b_i_1_N0), .preset(1'b0), 
        .next_state(coeffs_ff[64]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[31]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_1_Q_reg_17_ ( .clear(DP_reg_b_i_1_N0), .preset(1'b0), 
        .next_state(coeffs_ff[65]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[30]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_1_Q_reg_18_ ( .clear(DP_reg_b_i_1_N0), .preset(1'b0), 
        .next_state(coeffs_ff[66]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[29]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_1_Q_reg_19_ ( .clear(DP_reg_b_i_1_N0), .preset(1'b0), 
        .next_state(coeffs_ff[67]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[28]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_1_Q_reg_20_ ( .clear(DP_reg_b_i_1_N0), .preset(1'b0), 
        .next_state(coeffs_ff[68]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[27]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_1_Q_reg_21_ ( .clear(DP_reg_b_i_1_N0), .preset(1'b0), 
        .next_state(coeffs_ff[69]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[26]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_1_Q_reg_22_ ( .clear(DP_reg_b_i_1_N0), .preset(1'b0), 
        .next_state(coeffs_ff[70]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[25]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_1_Q_reg_23_ ( .clear(DP_reg_b_i_1_N0), .preset(1'b0), 
        .next_state(coeffs_ff[71]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[24]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  GTECH_NOT DP_reg_b_i_2_I_0 ( .A(rst_n), .Z(DP_reg_b_i_2_N0) );
  \**SEQGEN**  DP_reg_b_i_2_Q_reg_0_ ( .clear(DP_reg_b_i_2_N0), .preset(1'b0), 
        .next_state(coeffs_ff[24]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[71]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_2_Q_reg_1_ ( .clear(DP_reg_b_i_2_N0), .preset(1'b0), 
        .next_state(coeffs_ff[25]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[70]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_2_Q_reg_2_ ( .clear(DP_reg_b_i_2_N0), .preset(1'b0), 
        .next_state(coeffs_ff[26]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[69]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_2_Q_reg_3_ ( .clear(DP_reg_b_i_2_N0), .preset(1'b0), 
        .next_state(coeffs_ff[27]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[68]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_2_Q_reg_4_ ( .clear(DP_reg_b_i_2_N0), .preset(1'b0), 
        .next_state(coeffs_ff[28]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[67]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_2_Q_reg_5_ ( .clear(DP_reg_b_i_2_N0), .preset(1'b0), 
        .next_state(coeffs_ff[29]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[66]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_2_Q_reg_6_ ( .clear(DP_reg_b_i_2_N0), .preset(1'b0), 
        .next_state(coeffs_ff[30]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[65]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_2_Q_reg_7_ ( .clear(DP_reg_b_i_2_N0), .preset(1'b0), 
        .next_state(coeffs_ff[31]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[64]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_2_Q_reg_8_ ( .clear(DP_reg_b_i_2_N0), .preset(1'b0), 
        .next_state(coeffs_ff[32]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[63]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_2_Q_reg_9_ ( .clear(DP_reg_b_i_2_N0), .preset(1'b0), 
        .next_state(coeffs_ff[33]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[62]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_2_Q_reg_10_ ( .clear(DP_reg_b_i_2_N0), .preset(1'b0), 
        .next_state(coeffs_ff[34]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[61]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_2_Q_reg_11_ ( .clear(DP_reg_b_i_2_N0), .preset(1'b0), 
        .next_state(coeffs_ff[35]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[60]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_2_Q_reg_12_ ( .clear(DP_reg_b_i_2_N0), .preset(1'b0), 
        .next_state(coeffs_ff[36]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[59]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_2_Q_reg_13_ ( .clear(DP_reg_b_i_2_N0), .preset(1'b0), 
        .next_state(coeffs_ff[37]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[58]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_2_Q_reg_14_ ( .clear(DP_reg_b_i_2_N0), .preset(1'b0), 
        .next_state(coeffs_ff[38]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[57]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_2_Q_reg_15_ ( .clear(DP_reg_b_i_2_N0), .preset(1'b0), 
        .next_state(coeffs_ff[39]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[56]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_2_Q_reg_16_ ( .clear(DP_reg_b_i_2_N0), .preset(1'b0), 
        .next_state(coeffs_ff[40]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[55]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_2_Q_reg_17_ ( .clear(DP_reg_b_i_2_N0), .preset(1'b0), 
        .next_state(coeffs_ff[41]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[54]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_2_Q_reg_18_ ( .clear(DP_reg_b_i_2_N0), .preset(1'b0), 
        .next_state(coeffs_ff[42]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[53]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_2_Q_reg_19_ ( .clear(DP_reg_b_i_2_N0), .preset(1'b0), 
        .next_state(coeffs_ff[43]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[52]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_2_Q_reg_20_ ( .clear(DP_reg_b_i_2_N0), .preset(1'b0), 
        .next_state(coeffs_ff[44]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[51]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_2_Q_reg_21_ ( .clear(DP_reg_b_i_2_N0), .preset(1'b0), 
        .next_state(coeffs_ff[45]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[50]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_2_Q_reg_22_ ( .clear(DP_reg_b_i_2_N0), .preset(1'b0), 
        .next_state(coeffs_ff[46]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[49]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_2_Q_reg_23_ ( .clear(DP_reg_b_i_2_N0), .preset(1'b0), 
        .next_state(coeffs_ff[47]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[48]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  GTECH_NOT DP_reg_b_i_3_I_0 ( .A(rst_n), .Z(DP_reg_b_i_3_N0) );
  \**SEQGEN**  DP_reg_b_i_3_Q_reg_0_ ( .clear(DP_reg_b_i_3_N0), .preset(1'b0), 
        .next_state(coeffs_ff[0]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[95]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_3_Q_reg_1_ ( .clear(DP_reg_b_i_3_N0), .preset(1'b0), 
        .next_state(coeffs_ff[1]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[94]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_3_Q_reg_2_ ( .clear(DP_reg_b_i_3_N0), .preset(1'b0), 
        .next_state(coeffs_ff[2]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[93]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_3_Q_reg_3_ ( .clear(DP_reg_b_i_3_N0), .preset(1'b0), 
        .next_state(coeffs_ff[3]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[92]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_3_Q_reg_4_ ( .clear(DP_reg_b_i_3_N0), .preset(1'b0), 
        .next_state(coeffs_ff[4]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[91]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_3_Q_reg_5_ ( .clear(DP_reg_b_i_3_N0), .preset(1'b0), 
        .next_state(coeffs_ff[5]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[90]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_3_Q_reg_6_ ( .clear(DP_reg_b_i_3_N0), .preset(1'b0), 
        .next_state(coeffs_ff[6]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[89]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_3_Q_reg_7_ ( .clear(DP_reg_b_i_3_N0), .preset(1'b0), 
        .next_state(coeffs_ff[7]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[88]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_3_Q_reg_8_ ( .clear(DP_reg_b_i_3_N0), .preset(1'b0), 
        .next_state(coeffs_ff[8]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[87]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_3_Q_reg_9_ ( .clear(DP_reg_b_i_3_N0), .preset(1'b0), 
        .next_state(coeffs_ff[9]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[86]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_3_Q_reg_10_ ( .clear(DP_reg_b_i_3_N0), .preset(1'b0), 
        .next_state(coeffs_ff[10]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[85]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_3_Q_reg_11_ ( .clear(DP_reg_b_i_3_N0), .preset(1'b0), 
        .next_state(coeffs_ff[11]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[84]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_3_Q_reg_12_ ( .clear(DP_reg_b_i_3_N0), .preset(1'b0), 
        .next_state(coeffs_ff[12]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[83]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_3_Q_reg_13_ ( .clear(DP_reg_b_i_3_N0), .preset(1'b0), 
        .next_state(coeffs_ff[13]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[82]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_3_Q_reg_14_ ( .clear(DP_reg_b_i_3_N0), .preset(1'b0), 
        .next_state(coeffs_ff[14]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[81]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_3_Q_reg_15_ ( .clear(DP_reg_b_i_3_N0), .preset(1'b0), 
        .next_state(coeffs_ff[15]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[80]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_3_Q_reg_16_ ( .clear(DP_reg_b_i_3_N0), .preset(1'b0), 
        .next_state(coeffs_ff[16]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[79]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_3_Q_reg_17_ ( .clear(DP_reg_b_i_3_N0), .preset(1'b0), 
        .next_state(coeffs_ff[17]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[78]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_3_Q_reg_18_ ( .clear(DP_reg_b_i_3_N0), .preset(1'b0), 
        .next_state(coeffs_ff[18]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[77]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_3_Q_reg_19_ ( .clear(DP_reg_b_i_3_N0), .preset(1'b0), 
        .next_state(coeffs_ff[19]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[76]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_3_Q_reg_20_ ( .clear(DP_reg_b_i_3_N0), .preset(1'b0), 
        .next_state(coeffs_ff[20]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[75]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_3_Q_reg_21_ ( .clear(DP_reg_b_i_3_N0), .preset(1'b0), 
        .next_state(coeffs_ff[21]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[74]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_3_Q_reg_22_ ( .clear(DP_reg_b_i_3_N0), .preset(1'b0), 
        .next_state(coeffs_ff[22]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[73]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  \**SEQGEN**  DP_reg_b_i_3_Q_reg_23_ ( .clear(DP_reg_b_i_3_N0), .preset(1'b0), 
        .next_state(coeffs_ff[23]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_coeffs_ff_int[72]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(vIn) );
  GTECH_NOT DP_reg_sw0_I_0 ( .A(rst_n), .Z(DP_reg_sw0_N0) );
  \**SEQGEN**  DP_reg_sw0_Q_reg_0_ ( .clear(DP_reg_sw0_N0), .preset(1'b0), 
        .next_state(DP_w_0_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_sw0_0_), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw0_Q_reg_1_ ( .clear(DP_reg_sw0_N0), .preset(1'b0), 
        .next_state(DP_w_1_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_sw0_1_), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw0_Q_reg_2_ ( .clear(DP_reg_sw0_N0), .preset(1'b0), 
        .next_state(DP_w_2_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_sw0_2_), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw0_Q_reg_3_ ( .clear(DP_reg_sw0_N0), .preset(1'b0), 
        .next_state(DP_w_3_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_sw0_3_), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw0_Q_reg_4_ ( .clear(DP_reg_sw0_N0), .preset(1'b0), 
        .next_state(DP_w_4_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_sw0_4_), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw0_Q_reg_5_ ( .clear(DP_reg_sw0_N0), .preset(1'b0), 
        .next_state(DP_w_5_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_sw0_5_), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw0_Q_reg_6_ ( .clear(DP_reg_sw0_N0), .preset(1'b0), 
        .next_state(DP_w_6_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_sw0_6_), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw0_Q_reg_7_ ( .clear(DP_reg_sw0_N0), .preset(1'b0), 
        .next_state(DP_w_7_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_sw0_7_), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw0_Q_reg_8_ ( .clear(DP_reg_sw0_N0), .preset(1'b0), 
        .next_state(DP_w_8_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_sw0_8_), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw0_Q_reg_9_ ( .clear(DP_reg_sw0_N0), .preset(1'b0), 
        .next_state(DP_w_9_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_sw0_9_), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw0_Q_reg_10_ ( .clear(DP_reg_sw0_N0), .preset(1'b0), 
        .next_state(DP_w_10_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_sw0_10_), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw0_Q_reg_11_ ( .clear(DP_reg_sw0_N0), .preset(1'b0), 
        .next_state(DP_w_11_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_sw0_11_), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw0_Q_reg_12_ ( .clear(DP_reg_sw0_N0), .preset(1'b0), 
        .next_state(DP_w_12_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_sw0_12_), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw0_Q_reg_13_ ( .clear(DP_reg_sw0_N0), .preset(1'b0), 
        .next_state(DP_w_13_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_sw0_13_), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw0_Q_reg_14_ ( .clear(DP_reg_sw0_N0), .preset(1'b0), 
        .next_state(DP_w_14_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_sw0_14_), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw0_Q_reg_15_ ( .clear(DP_reg_sw0_N0), .preset(1'b0), 
        .next_state(DP_w_15_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_sw0_15_), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw0_Q_reg_16_ ( .clear(DP_reg_sw0_N0), .preset(1'b0), 
        .next_state(DP_w_16_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_sw0_16_), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw0_Q_reg_17_ ( .clear(DP_reg_sw0_N0), .preset(1'b0), 
        .next_state(DP_w_17_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_sw0_17_), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw0_Q_reg_18_ ( .clear(DP_reg_sw0_N0), .preset(1'b0), 
        .next_state(DP_w_18_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_sw0_18_), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw0_Q_reg_19_ ( .clear(DP_reg_sw0_N0), .preset(1'b0), 
        .next_state(DP_w_19_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_sw0_19_), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw0_Q_reg_20_ ( .clear(DP_reg_sw0_N0), .preset(1'b0), 
        .next_state(DP_w_20_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_sw0_20_), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw0_Q_reg_21_ ( .clear(DP_reg_sw0_N0), .preset(1'b0), 
        .next_state(DP_w_21_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_sw0_21_), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw0_Q_reg_22_ ( .clear(DP_reg_sw0_N0), .preset(1'b0), 
        .next_state(DP_w_22_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_sw0_22_), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw0_Q_reg_23_ ( .clear(DP_reg_sw0_N0), .preset(1'b0), 
        .next_state(DP_w_23_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), 
        .Q(DP_sw0_23_), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  GTECH_NOT DP_reg_sw1_I_0 ( .A(rst_n), .Z(DP_reg_sw1_N0) );
  \**SEQGEN**  DP_reg_sw1_Q_reg_0_ ( .clear(DP_reg_sw1_N0), .preset(1'b0), 
        .next_state(DP_sw0_0_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(DP_sw1_0_), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw1_Q_reg_1_ ( .clear(DP_reg_sw1_N0), .preset(1'b0), 
        .next_state(DP_sw0_1_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(DP_sw1_1_), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw1_Q_reg_2_ ( .clear(DP_reg_sw1_N0), .preset(1'b0), 
        .next_state(DP_sw0_2_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(DP_sw1_2_), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw1_Q_reg_3_ ( .clear(DP_reg_sw1_N0), .preset(1'b0), 
        .next_state(DP_sw0_3_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(DP_sw1_3_), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw1_Q_reg_4_ ( .clear(DP_reg_sw1_N0), .preset(1'b0), 
        .next_state(DP_sw0_4_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(DP_sw1_4_), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw1_Q_reg_5_ ( .clear(DP_reg_sw1_N0), .preset(1'b0), 
        .next_state(DP_sw0_5_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(DP_sw1_5_), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw1_Q_reg_6_ ( .clear(DP_reg_sw1_N0), .preset(1'b0), 
        .next_state(DP_sw0_6_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(DP_sw1_6_), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw1_Q_reg_7_ ( .clear(DP_reg_sw1_N0), .preset(1'b0), 
        .next_state(DP_sw0_7_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(DP_sw1_7_), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw1_Q_reg_8_ ( .clear(DP_reg_sw1_N0), .preset(1'b0), 
        .next_state(DP_sw0_8_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(DP_sw1_8_), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw1_Q_reg_9_ ( .clear(DP_reg_sw1_N0), .preset(1'b0), 
        .next_state(DP_sw0_9_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(DP_sw1_9_), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw1_Q_reg_10_ ( .clear(DP_reg_sw1_N0), .preset(1'b0), 
        .next_state(DP_sw0_10_), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_sw1_10_), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw1_Q_reg_11_ ( .clear(DP_reg_sw1_N0), .preset(1'b0), 
        .next_state(DP_sw0_11_), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_sw1_11_), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw1_Q_reg_12_ ( .clear(DP_reg_sw1_N0), .preset(1'b0), 
        .next_state(DP_sw0_12_), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_sw1_12_), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw1_Q_reg_13_ ( .clear(DP_reg_sw1_N0), .preset(1'b0), 
        .next_state(DP_sw0_13_), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_sw1_13_), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw1_Q_reg_14_ ( .clear(DP_reg_sw1_N0), .preset(1'b0), 
        .next_state(DP_sw0_14_), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_sw1_14_), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw1_Q_reg_15_ ( .clear(DP_reg_sw1_N0), .preset(1'b0), 
        .next_state(DP_sw0_15_), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_sw1_15_), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw1_Q_reg_16_ ( .clear(DP_reg_sw1_N0), .preset(1'b0), 
        .next_state(DP_sw0_16_), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_sw1_16_), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw1_Q_reg_17_ ( .clear(DP_reg_sw1_N0), .preset(1'b0), 
        .next_state(DP_sw0_17_), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_sw1_17_), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw1_Q_reg_18_ ( .clear(DP_reg_sw1_N0), .preset(1'b0), 
        .next_state(DP_sw0_18_), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_sw1_18_), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw1_Q_reg_19_ ( .clear(DP_reg_sw1_N0), .preset(1'b0), 
        .next_state(DP_sw0_19_), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_sw1_19_), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw1_Q_reg_20_ ( .clear(DP_reg_sw1_N0), .preset(1'b0), 
        .next_state(DP_sw0_20_), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_sw1_20_), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw1_Q_reg_21_ ( .clear(DP_reg_sw1_N0), .preset(1'b0), 
        .next_state(DP_sw0_21_), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_sw1_21_), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw1_Q_reg_22_ ( .clear(DP_reg_sw1_N0), .preset(1'b0), 
        .next_state(DP_sw0_22_), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_sw1_22_), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw1_Q_reg_23_ ( .clear(DP_reg_sw1_N0), .preset(1'b0), 
        .next_state(DP_sw0_23_), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_sw1_23_), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  GTECH_NOT DP_reg_sw2_I_0 ( .A(rst_n), .Z(DP_reg_sw2_N0) );
  \**SEQGEN**  DP_reg_sw2_Q_reg_0_ ( .clear(DP_reg_sw2_N0), .preset(1'b0), 
        .next_state(DP_sw1_0_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(DP_sw2[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw2_Q_reg_1_ ( .clear(DP_reg_sw2_N0), .preset(1'b0), 
        .next_state(DP_sw1_1_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(DP_sw2[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw2_Q_reg_2_ ( .clear(DP_reg_sw2_N0), .preset(1'b0), 
        .next_state(DP_sw1_2_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(DP_sw2[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw2_Q_reg_3_ ( .clear(DP_reg_sw2_N0), .preset(1'b0), 
        .next_state(DP_sw1_3_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(DP_sw2[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw2_Q_reg_4_ ( .clear(DP_reg_sw2_N0), .preset(1'b0), 
        .next_state(DP_sw1_4_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(DP_sw2[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw2_Q_reg_5_ ( .clear(DP_reg_sw2_N0), .preset(1'b0), 
        .next_state(DP_sw1_5_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(DP_sw2[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw2_Q_reg_6_ ( .clear(DP_reg_sw2_N0), .preset(1'b0), 
        .next_state(DP_sw1_6_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(DP_sw2[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw2_Q_reg_7_ ( .clear(DP_reg_sw2_N0), .preset(1'b0), 
        .next_state(DP_sw1_7_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(DP_sw2[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw2_Q_reg_8_ ( .clear(DP_reg_sw2_N0), .preset(1'b0), 
        .next_state(DP_sw1_8_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(DP_sw2[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw2_Q_reg_9_ ( .clear(DP_reg_sw2_N0), .preset(1'b0), 
        .next_state(DP_sw1_9_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(DP_sw2[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw2_Q_reg_10_ ( .clear(DP_reg_sw2_N0), .preset(1'b0), 
        .next_state(DP_sw1_10_), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_sw2[10]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw2_Q_reg_11_ ( .clear(DP_reg_sw2_N0), .preset(1'b0), 
        .next_state(DP_sw1_11_), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_sw2[11]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw2_Q_reg_12_ ( .clear(DP_reg_sw2_N0), .preset(1'b0), 
        .next_state(DP_sw1_12_), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_sw2[12]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw2_Q_reg_13_ ( .clear(DP_reg_sw2_N0), .preset(1'b0), 
        .next_state(DP_sw1_13_), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_sw2[13]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw2_Q_reg_14_ ( .clear(DP_reg_sw2_N0), .preset(1'b0), 
        .next_state(DP_sw1_14_), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_sw2[14]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw2_Q_reg_15_ ( .clear(DP_reg_sw2_N0), .preset(1'b0), 
        .next_state(DP_sw1_15_), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_sw2[15]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw2_Q_reg_16_ ( .clear(DP_reg_sw2_N0), .preset(1'b0), 
        .next_state(DP_sw1_16_), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_sw2[16]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw2_Q_reg_17_ ( .clear(DP_reg_sw2_N0), .preset(1'b0), 
        .next_state(DP_sw1_17_), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_sw2[17]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw2_Q_reg_18_ ( .clear(DP_reg_sw2_N0), .preset(1'b0), 
        .next_state(DP_sw1_18_), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_sw2[18]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw2_Q_reg_19_ ( .clear(DP_reg_sw2_N0), .preset(1'b0), 
        .next_state(DP_sw1_19_), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_sw2[19]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw2_Q_reg_20_ ( .clear(DP_reg_sw2_N0), .preset(1'b0), 
        .next_state(DP_sw1_20_), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_sw2[20]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw2_Q_reg_21_ ( .clear(DP_reg_sw2_N0), .preset(1'b0), 
        .next_state(DP_sw1_21_), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_sw2[21]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw2_Q_reg_22_ ( .clear(DP_reg_sw2_N0), .preset(1'b0), 
        .next_state(DP_sw1_22_), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_sw2[22]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  \**SEQGEN**  DP_reg_sw2_Q_reg_23_ ( .clear(DP_reg_sw2_N0), .preset(1'b0), 
        .next_state(DP_sw1_23_), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(DP_sw2[23]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(sw_regs_en_int) );
  GTECH_NOT DP_reg_ret0_I_0 ( .A(rst_n), .Z(DP_reg_ret0_N0) );
  \**SEQGEN**  DP_reg_ret0_Q_reg_0_ ( .clear(DP_reg_ret0_N0), .preset(1'b0), 
        .next_state(DP_sw0_coeff_ret0[0]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret0[0]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret0_Q_reg_1_ ( .clear(DP_reg_ret0_N0), .preset(1'b0), 
        .next_state(DP_sw0_coeff_ret0[1]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret0[1]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret0_Q_reg_2_ ( .clear(DP_reg_ret0_N0), .preset(1'b0), 
        .next_state(DP_sw0_coeff_ret0[2]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret0[2]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret0_Q_reg_3_ ( .clear(DP_reg_ret0_N0), .preset(1'b0), 
        .next_state(DP_sw0_coeff_ret0[3]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret0[3]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret0_Q_reg_4_ ( .clear(DP_reg_ret0_N0), .preset(1'b0), 
        .next_state(DP_sw0_coeff_ret0[4]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret0[4]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret0_Q_reg_5_ ( .clear(DP_reg_ret0_N0), .preset(1'b0), 
        .next_state(DP_sw0_coeff_ret0[5]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret0[5]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret0_Q_reg_6_ ( .clear(DP_reg_ret0_N0), .preset(1'b0), 
        .next_state(DP_sw0_coeff_ret0[6]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret0[6]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret0_Q_reg_7_ ( .clear(DP_reg_ret0_N0), .preset(1'b0), 
        .next_state(DP_sw0_coeff_ret0[7]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret0[7]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret0_Q_reg_8_ ( .clear(DP_reg_ret0_N0), .preset(1'b0), 
        .next_state(DP_sw0_coeff_ret0[8]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret0[8]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret0_Q_reg_9_ ( .clear(DP_reg_ret0_N0), .preset(1'b0), 
        .next_state(DP_sw0_coeff_ret0[9]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret0[9]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret0_Q_reg_10_ ( .clear(DP_reg_ret0_N0), .preset(1'b0), 
        .next_state(DP_sw0_coeff_ret0[10]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret0[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret0_Q_reg_11_ ( .clear(DP_reg_ret0_N0), .preset(1'b0), 
        .next_state(DP_sw0_coeff_ret0[11]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret0[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret0_Q_reg_12_ ( .clear(DP_reg_ret0_N0), .preset(1'b0), 
        .next_state(DP_sw0_coeff_ret0[12]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret0[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret0_Q_reg_13_ ( .clear(DP_reg_ret0_N0), .preset(1'b0), 
        .next_state(DP_sw0_coeff_ret0[13]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret0[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret0_Q_reg_14_ ( .clear(DP_reg_ret0_N0), .preset(1'b0), 
        .next_state(DP_sw0_coeff_ret0[14]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret0[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret0_Q_reg_15_ ( .clear(DP_reg_ret0_N0), .preset(1'b0), 
        .next_state(DP_sw0_coeff_ret0[15]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret0[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret0_Q_reg_16_ ( .clear(DP_reg_ret0_N0), .preset(1'b0), 
        .next_state(DP_sw0_coeff_ret0[16]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret0[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret0_Q_reg_17_ ( .clear(DP_reg_ret0_N0), .preset(1'b0), 
        .next_state(DP_sw0_coeff_ret0[17]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret0[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret0_Q_reg_18_ ( .clear(DP_reg_ret0_N0), .preset(1'b0), 
        .next_state(DP_sw0_coeff_ret0[18]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret0[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret0_Q_reg_19_ ( .clear(DP_reg_ret0_N0), .preset(1'b0), 
        .next_state(DP_sw0_coeff_ret0[19]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret0[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret0_Q_reg_20_ ( .clear(DP_reg_ret0_N0), .preset(1'b0), 
        .next_state(DP_sw0_coeff_ret0[20]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret0[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret0_Q_reg_21_ ( .clear(DP_reg_ret0_N0), .preset(1'b0), 
        .next_state(DP_sw0_coeff_ret0[21]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret0[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret0_Q_reg_22_ ( .clear(DP_reg_ret0_N0), .preset(1'b0), 
        .next_state(DP_sw0_coeff_ret0[22]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret0[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret0_Q_reg_23_ ( .clear(DP_reg_ret0_N0), .preset(1'b0), 
        .next_state(DP_sw0_coeff_ret0[23]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret0[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  GTECH_NOT DP_reg_ret1_I_0 ( .A(rst_n), .Z(DP_reg_ret1_N0) );
  \**SEQGEN**  DP_reg_ret1_Q_reg_0_ ( .clear(DP_reg_ret1_N0), .preset(1'b0), 
        .next_state(DP_sw1_coeff_ret1[0]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret1[0]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret1_Q_reg_1_ ( .clear(DP_reg_ret1_N0), .preset(1'b0), 
        .next_state(DP_sw1_coeff_ret1[1]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret1[1]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret1_Q_reg_2_ ( .clear(DP_reg_ret1_N0), .preset(1'b0), 
        .next_state(DP_sw1_coeff_ret1[2]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret1[2]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret1_Q_reg_3_ ( .clear(DP_reg_ret1_N0), .preset(1'b0), 
        .next_state(DP_sw1_coeff_ret1[3]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret1[3]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret1_Q_reg_4_ ( .clear(DP_reg_ret1_N0), .preset(1'b0), 
        .next_state(DP_sw1_coeff_ret1[4]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret1[4]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret1_Q_reg_5_ ( .clear(DP_reg_ret1_N0), .preset(1'b0), 
        .next_state(DP_sw1_coeff_ret1[5]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret1[5]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret1_Q_reg_6_ ( .clear(DP_reg_ret1_N0), .preset(1'b0), 
        .next_state(DP_sw1_coeff_ret1[6]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret1[6]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret1_Q_reg_7_ ( .clear(DP_reg_ret1_N0), .preset(1'b0), 
        .next_state(DP_sw1_coeff_ret1[7]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret1[7]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret1_Q_reg_8_ ( .clear(DP_reg_ret1_N0), .preset(1'b0), 
        .next_state(DP_sw1_coeff_ret1[8]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret1[8]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret1_Q_reg_9_ ( .clear(DP_reg_ret1_N0), .preset(1'b0), 
        .next_state(DP_sw1_coeff_ret1[9]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret1[9]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret1_Q_reg_10_ ( .clear(DP_reg_ret1_N0), .preset(1'b0), 
        .next_state(DP_sw1_coeff_ret1[10]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret1[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret1_Q_reg_11_ ( .clear(DP_reg_ret1_N0), .preset(1'b0), 
        .next_state(DP_sw1_coeff_ret1[11]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret1[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret1_Q_reg_12_ ( .clear(DP_reg_ret1_N0), .preset(1'b0), 
        .next_state(DP_sw1_coeff_ret1[12]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret1[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret1_Q_reg_13_ ( .clear(DP_reg_ret1_N0), .preset(1'b0), 
        .next_state(DP_sw1_coeff_ret1[13]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret1[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret1_Q_reg_14_ ( .clear(DP_reg_ret1_N0), .preset(1'b0), 
        .next_state(DP_sw1_coeff_ret1[14]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret1[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret1_Q_reg_15_ ( .clear(DP_reg_ret1_N0), .preset(1'b0), 
        .next_state(DP_sw1_coeff_ret1[15]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret1[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret1_Q_reg_16_ ( .clear(DP_reg_ret1_N0), .preset(1'b0), 
        .next_state(DP_sw1_coeff_ret1[16]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret1[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret1_Q_reg_17_ ( .clear(DP_reg_ret1_N0), .preset(1'b0), 
        .next_state(DP_sw1_coeff_ret1[17]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret1[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret1_Q_reg_18_ ( .clear(DP_reg_ret1_N0), .preset(1'b0), 
        .next_state(DP_sw1_coeff_ret1[18]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret1[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret1_Q_reg_19_ ( .clear(DP_reg_ret1_N0), .preset(1'b0), 
        .next_state(DP_sw1_coeff_ret1[19]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret1[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret1_Q_reg_20_ ( .clear(DP_reg_ret1_N0), .preset(1'b0), 
        .next_state(DP_sw1_coeff_ret1[20]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret1[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret1_Q_reg_21_ ( .clear(DP_reg_ret1_N0), .preset(1'b0), 
        .next_state(DP_sw1_coeff_ret1[21]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret1[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret1_Q_reg_22_ ( .clear(DP_reg_ret1_N0), .preset(1'b0), 
        .next_state(DP_sw1_coeff_ret1[22]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret1[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_ret1_Q_reg_23_ ( .clear(DP_reg_ret1_N0), .preset(1'b0), 
        .next_state(DP_sw1_coeff_ret1[23]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_ret1[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  GTECH_NOT DP_reg_pipe00_I_0 ( .A(rst_n), .Z(DP_reg_pipe00_N0) );
  \**SEQGEN**  DP_reg_pipe00_Q_reg_0_ ( .clear(DP_reg_pipe00_N0), .preset(1'b0), .next_state(DP_w_0_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe00[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe00_Q_reg_1_ ( .clear(DP_reg_pipe00_N0), .preset(1'b0), .next_state(DP_w_1_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe00[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe00_Q_reg_2_ ( .clear(DP_reg_pipe00_N0), .preset(1'b0), .next_state(DP_w_2_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe00[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe00_Q_reg_3_ ( .clear(DP_reg_pipe00_N0), .preset(1'b0), .next_state(DP_w_3_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe00[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe00_Q_reg_4_ ( .clear(DP_reg_pipe00_N0), .preset(1'b0), .next_state(DP_w_4_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe00[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe00_Q_reg_5_ ( .clear(DP_reg_pipe00_N0), .preset(1'b0), .next_state(DP_w_5_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe00[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe00_Q_reg_6_ ( .clear(DP_reg_pipe00_N0), .preset(1'b0), .next_state(DP_w_6_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe00[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe00_Q_reg_7_ ( .clear(DP_reg_pipe00_N0), .preset(1'b0), .next_state(DP_w_7_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe00[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe00_Q_reg_8_ ( .clear(DP_reg_pipe00_N0), .preset(1'b0), .next_state(DP_w_8_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe00[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe00_Q_reg_9_ ( .clear(DP_reg_pipe00_N0), .preset(1'b0), .next_state(DP_w_9_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe00[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe00_Q_reg_10_ ( .clear(DP_reg_pipe00_N0), .preset(
        1'b0), .next_state(DP_w_10_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe00[10]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe00_Q_reg_11_ ( .clear(DP_reg_pipe00_N0), .preset(
        1'b0), .next_state(DP_w_11_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe00[11]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe00_Q_reg_12_ ( .clear(DP_reg_pipe00_N0), .preset(
        1'b0), .next_state(DP_w_12_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe00[12]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe00_Q_reg_13_ ( .clear(DP_reg_pipe00_N0), .preset(
        1'b0), .next_state(DP_w_13_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe00[13]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe00_Q_reg_14_ ( .clear(DP_reg_pipe00_N0), .preset(
        1'b0), .next_state(DP_w_14_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe00[14]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe00_Q_reg_15_ ( .clear(DP_reg_pipe00_N0), .preset(
        1'b0), .next_state(DP_w_15_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe00[15]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe00_Q_reg_16_ ( .clear(DP_reg_pipe00_N0), .preset(
        1'b0), .next_state(DP_w_16_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe00[16]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe00_Q_reg_17_ ( .clear(DP_reg_pipe00_N0), .preset(
        1'b0), .next_state(DP_w_17_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe00[17]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe00_Q_reg_18_ ( .clear(DP_reg_pipe00_N0), .preset(
        1'b0), .next_state(DP_w_18_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe00[18]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe00_Q_reg_19_ ( .clear(DP_reg_pipe00_N0), .preset(
        1'b0), .next_state(DP_w_19_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe00[19]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe00_Q_reg_20_ ( .clear(DP_reg_pipe00_N0), .preset(
        1'b0), .next_state(DP_w_20_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe00[20]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe00_Q_reg_21_ ( .clear(DP_reg_pipe00_N0), .preset(
        1'b0), .next_state(DP_w_21_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe00[21]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe00_Q_reg_22_ ( .clear(DP_reg_pipe00_N0), .preset(
        1'b0), .next_state(DP_w_22_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe00[22]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe00_Q_reg_23_ ( .clear(DP_reg_pipe00_N0), .preset(
        1'b0), .next_state(DP_w_23_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe00[23]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  GTECH_NOT DP_reg_pipe01_I_0 ( .A(rst_n), .Z(DP_reg_pipe01_N0) );
  \**SEQGEN**  DP_reg_pipe01_Q_reg_0_ ( .clear(DP_reg_pipe01_N0), .preset(1'b0), .next_state(DP_sw0_0_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe01[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe01_Q_reg_1_ ( .clear(DP_reg_pipe01_N0), .preset(1'b0), .next_state(DP_sw0_1_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe01[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe01_Q_reg_2_ ( .clear(DP_reg_pipe01_N0), .preset(1'b0), .next_state(DP_sw0_2_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe01[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe01_Q_reg_3_ ( .clear(DP_reg_pipe01_N0), .preset(1'b0), .next_state(DP_sw0_3_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe01[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe01_Q_reg_4_ ( .clear(DP_reg_pipe01_N0), .preset(1'b0), .next_state(DP_sw0_4_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe01[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe01_Q_reg_5_ ( .clear(DP_reg_pipe01_N0), .preset(1'b0), .next_state(DP_sw0_5_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe01[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe01_Q_reg_6_ ( .clear(DP_reg_pipe01_N0), .preset(1'b0), .next_state(DP_sw0_6_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe01[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe01_Q_reg_7_ ( .clear(DP_reg_pipe01_N0), .preset(1'b0), .next_state(DP_sw0_7_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe01[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe01_Q_reg_8_ ( .clear(DP_reg_pipe01_N0), .preset(1'b0), .next_state(DP_sw0_8_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe01[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe01_Q_reg_9_ ( .clear(DP_reg_pipe01_N0), .preset(1'b0), .next_state(DP_sw0_9_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe01[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe01_Q_reg_10_ ( .clear(DP_reg_pipe01_N0), .preset(
        1'b0), .next_state(DP_sw0_10_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe01[10]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe01_Q_reg_11_ ( .clear(DP_reg_pipe01_N0), .preset(
        1'b0), .next_state(DP_sw0_11_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe01[11]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe01_Q_reg_12_ ( .clear(DP_reg_pipe01_N0), .preset(
        1'b0), .next_state(DP_sw0_12_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe01[12]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe01_Q_reg_13_ ( .clear(DP_reg_pipe01_N0), .preset(
        1'b0), .next_state(DP_sw0_13_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe01[13]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe01_Q_reg_14_ ( .clear(DP_reg_pipe01_N0), .preset(
        1'b0), .next_state(DP_sw0_14_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe01[14]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe01_Q_reg_15_ ( .clear(DP_reg_pipe01_N0), .preset(
        1'b0), .next_state(DP_sw0_15_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe01[15]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe01_Q_reg_16_ ( .clear(DP_reg_pipe01_N0), .preset(
        1'b0), .next_state(DP_sw0_16_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe01[16]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe01_Q_reg_17_ ( .clear(DP_reg_pipe01_N0), .preset(
        1'b0), .next_state(DP_sw0_17_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe01[17]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe01_Q_reg_18_ ( .clear(DP_reg_pipe01_N0), .preset(
        1'b0), .next_state(DP_sw0_18_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe01[18]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe01_Q_reg_19_ ( .clear(DP_reg_pipe01_N0), .preset(
        1'b0), .next_state(DP_sw0_19_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe01[19]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe01_Q_reg_20_ ( .clear(DP_reg_pipe01_N0), .preset(
        1'b0), .next_state(DP_sw0_20_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe01[20]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe01_Q_reg_21_ ( .clear(DP_reg_pipe01_N0), .preset(
        1'b0), .next_state(DP_sw0_21_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe01[21]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe01_Q_reg_22_ ( .clear(DP_reg_pipe01_N0), .preset(
        1'b0), .next_state(DP_sw0_22_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe01[22]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe01_Q_reg_23_ ( .clear(DP_reg_pipe01_N0), .preset(
        1'b0), .next_state(DP_sw0_23_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe01[23]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  GTECH_NOT DP_reg_pipe02_I_0 ( .A(rst_n), .Z(DP_reg_pipe02_N0) );
  \**SEQGEN**  DP_reg_pipe02_Q_reg_0_ ( .clear(DP_reg_pipe02_N0), .preset(1'b0), .next_state(DP_sw1_0_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe02[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe02_Q_reg_1_ ( .clear(DP_reg_pipe02_N0), .preset(1'b0), .next_state(DP_sw1_1_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe02[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe02_Q_reg_2_ ( .clear(DP_reg_pipe02_N0), .preset(1'b0), .next_state(DP_sw1_2_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe02[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe02_Q_reg_3_ ( .clear(DP_reg_pipe02_N0), .preset(1'b0), .next_state(DP_sw1_3_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe02[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe02_Q_reg_4_ ( .clear(DP_reg_pipe02_N0), .preset(1'b0), .next_state(DP_sw1_4_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe02[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe02_Q_reg_5_ ( .clear(DP_reg_pipe02_N0), .preset(1'b0), .next_state(DP_sw1_5_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe02[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe02_Q_reg_6_ ( .clear(DP_reg_pipe02_N0), .preset(1'b0), .next_state(DP_sw1_6_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe02[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe02_Q_reg_7_ ( .clear(DP_reg_pipe02_N0), .preset(1'b0), .next_state(DP_sw1_7_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe02[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe02_Q_reg_8_ ( .clear(DP_reg_pipe02_N0), .preset(1'b0), .next_state(DP_sw1_8_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe02[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe02_Q_reg_9_ ( .clear(DP_reg_pipe02_N0), .preset(1'b0), .next_state(DP_sw1_9_), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe02[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe02_Q_reg_10_ ( .clear(DP_reg_pipe02_N0), .preset(
        1'b0), .next_state(DP_sw1_10_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe02[10]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe02_Q_reg_11_ ( .clear(DP_reg_pipe02_N0), .preset(
        1'b0), .next_state(DP_sw1_11_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe02[11]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe02_Q_reg_12_ ( .clear(DP_reg_pipe02_N0), .preset(
        1'b0), .next_state(DP_sw1_12_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe02[12]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe02_Q_reg_13_ ( .clear(DP_reg_pipe02_N0), .preset(
        1'b0), .next_state(DP_sw1_13_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe02[13]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe02_Q_reg_14_ ( .clear(DP_reg_pipe02_N0), .preset(
        1'b0), .next_state(DP_sw1_14_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe02[14]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe02_Q_reg_15_ ( .clear(DP_reg_pipe02_N0), .preset(
        1'b0), .next_state(DP_sw1_15_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe02[15]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe02_Q_reg_16_ ( .clear(DP_reg_pipe02_N0), .preset(
        1'b0), .next_state(DP_sw1_16_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe02[16]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe02_Q_reg_17_ ( .clear(DP_reg_pipe02_N0), .preset(
        1'b0), .next_state(DP_sw1_17_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe02[17]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe02_Q_reg_18_ ( .clear(DP_reg_pipe02_N0), .preset(
        1'b0), .next_state(DP_sw1_18_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe02[18]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe02_Q_reg_19_ ( .clear(DP_reg_pipe02_N0), .preset(
        1'b0), .next_state(DP_sw1_19_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe02[19]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe02_Q_reg_20_ ( .clear(DP_reg_pipe02_N0), .preset(
        1'b0), .next_state(DP_sw1_20_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe02[20]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe02_Q_reg_21_ ( .clear(DP_reg_pipe02_N0), .preset(
        1'b0), .next_state(DP_sw1_21_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe02[21]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe02_Q_reg_22_ ( .clear(DP_reg_pipe02_N0), .preset(
        1'b0), .next_state(DP_sw1_22_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe02[22]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe02_Q_reg_23_ ( .clear(DP_reg_pipe02_N0), .preset(
        1'b0), .next_state(DP_sw1_23_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe02[23]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  GTECH_NOT DP_reg_pipe03_I_0 ( .A(rst_n), .Z(DP_reg_pipe03_N0) );
  \**SEQGEN**  DP_reg_pipe03_Q_reg_0_ ( .clear(DP_reg_pipe03_N0), .preset(1'b0), .next_state(DP_sw2[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe03[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe03_Q_reg_1_ ( .clear(DP_reg_pipe03_N0), .preset(1'b0), .next_state(DP_sw2[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe03[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe03_Q_reg_2_ ( .clear(DP_reg_pipe03_N0), .preset(1'b0), .next_state(DP_sw2[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe03[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe03_Q_reg_3_ ( .clear(DP_reg_pipe03_N0), .preset(1'b0), .next_state(DP_sw2[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe03[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe03_Q_reg_4_ ( .clear(DP_reg_pipe03_N0), .preset(1'b0), .next_state(DP_sw2[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe03[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe03_Q_reg_5_ ( .clear(DP_reg_pipe03_N0), .preset(1'b0), .next_state(DP_sw2[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe03[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe03_Q_reg_6_ ( .clear(DP_reg_pipe03_N0), .preset(1'b0), .next_state(DP_sw2[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe03[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe03_Q_reg_7_ ( .clear(DP_reg_pipe03_N0), .preset(1'b0), .next_state(DP_sw2[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe03[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe03_Q_reg_8_ ( .clear(DP_reg_pipe03_N0), .preset(1'b0), .next_state(DP_sw2[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe03[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe03_Q_reg_9_ ( .clear(DP_reg_pipe03_N0), .preset(1'b0), .next_state(DP_sw2[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        DP_pipe03[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe03_Q_reg_10_ ( .clear(DP_reg_pipe03_N0), .preset(
        1'b0), .next_state(DP_sw2[10]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe03[10]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe03_Q_reg_11_ ( .clear(DP_reg_pipe03_N0), .preset(
        1'b0), .next_state(DP_sw2[11]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe03[11]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe03_Q_reg_12_ ( .clear(DP_reg_pipe03_N0), .preset(
        1'b0), .next_state(DP_sw2[12]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe03[12]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe03_Q_reg_13_ ( .clear(DP_reg_pipe03_N0), .preset(
        1'b0), .next_state(DP_sw2[13]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe03[13]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe03_Q_reg_14_ ( .clear(DP_reg_pipe03_N0), .preset(
        1'b0), .next_state(DP_sw2[14]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe03[14]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe03_Q_reg_15_ ( .clear(DP_reg_pipe03_N0), .preset(
        1'b0), .next_state(DP_sw2[15]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe03[15]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe03_Q_reg_16_ ( .clear(DP_reg_pipe03_N0), .preset(
        1'b0), .next_state(DP_sw2[16]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe03[16]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe03_Q_reg_17_ ( .clear(DP_reg_pipe03_N0), .preset(
        1'b0), .next_state(DP_sw2[17]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe03[17]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe03_Q_reg_18_ ( .clear(DP_reg_pipe03_N0), .preset(
        1'b0), .next_state(DP_sw2[18]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe03[18]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe03_Q_reg_19_ ( .clear(DP_reg_pipe03_N0), .preset(
        1'b0), .next_state(DP_sw2[19]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe03[19]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe03_Q_reg_20_ ( .clear(DP_reg_pipe03_N0), .preset(
        1'b0), .next_state(DP_sw2[20]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe03[20]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe03_Q_reg_21_ ( .clear(DP_reg_pipe03_N0), .preset(
        1'b0), .next_state(DP_sw2[21]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe03[21]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe03_Q_reg_22_ ( .clear(DP_reg_pipe03_N0), .preset(
        1'b0), .next_state(DP_sw2[22]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe03[22]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe03_Q_reg_23_ ( .clear(DP_reg_pipe03_N0), .preset(
        1'b0), .next_state(DP_sw2[23]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe03[23]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  GTECH_NOT DP_reg_pipe10_I_0 ( .A(rst_n), .Z(DP_reg_pipe10_N0) );
  \**SEQGEN**  DP_reg_pipe10_Q_reg_0_ ( .clear(DP_reg_pipe10_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe00[0]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe10[0]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe10_Q_reg_1_ ( .clear(DP_reg_pipe10_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe00[1]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe10[1]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe10_Q_reg_2_ ( .clear(DP_reg_pipe10_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe00[2]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe10[2]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe10_Q_reg_3_ ( .clear(DP_reg_pipe10_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe00[3]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe10[3]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe10_Q_reg_4_ ( .clear(DP_reg_pipe10_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe00[4]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe10[4]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe10_Q_reg_5_ ( .clear(DP_reg_pipe10_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe00[5]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe10[5]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe10_Q_reg_6_ ( .clear(DP_reg_pipe10_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe00[6]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe10[6]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe10_Q_reg_7_ ( .clear(DP_reg_pipe10_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe00[7]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe10[7]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe10_Q_reg_8_ ( .clear(DP_reg_pipe10_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe00[8]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe10[8]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe10_Q_reg_9_ ( .clear(DP_reg_pipe10_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe00[9]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe10[9]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe10_Q_reg_10_ ( .clear(DP_reg_pipe10_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe00[10]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe10[10]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe10_Q_reg_11_ ( .clear(DP_reg_pipe10_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe00[11]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe10[11]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe10_Q_reg_12_ ( .clear(DP_reg_pipe10_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe00[12]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe10[12]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe10_Q_reg_13_ ( .clear(DP_reg_pipe10_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe00[13]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe10[13]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe10_Q_reg_14_ ( .clear(DP_reg_pipe10_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe00[14]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe10[14]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe10_Q_reg_15_ ( .clear(DP_reg_pipe10_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe00[15]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe10[15]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe10_Q_reg_16_ ( .clear(DP_reg_pipe10_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe00[16]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe10[16]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe10_Q_reg_17_ ( .clear(DP_reg_pipe10_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe00[17]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe10[17]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe10_Q_reg_18_ ( .clear(DP_reg_pipe10_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe00[18]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe10[18]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe10_Q_reg_19_ ( .clear(DP_reg_pipe10_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe00[19]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe10[19]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe10_Q_reg_20_ ( .clear(DP_reg_pipe10_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe00[20]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe10[20]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe10_Q_reg_21_ ( .clear(DP_reg_pipe10_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe00[21]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe10[21]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe10_Q_reg_22_ ( .clear(DP_reg_pipe10_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe00[22]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe10[22]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe10_Q_reg_23_ ( .clear(DP_reg_pipe10_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe00[23]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe10[23]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  GTECH_NOT DP_reg_pipe11_I_0 ( .A(rst_n), .Z(DP_reg_pipe11_N0) );
  \**SEQGEN**  DP_reg_pipe11_Q_reg_0_ ( .clear(DP_reg_pipe11_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe01[0]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe11[0]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe11_Q_reg_1_ ( .clear(DP_reg_pipe11_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe01[1]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe11[1]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe11_Q_reg_2_ ( .clear(DP_reg_pipe11_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe01[2]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe11[2]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe11_Q_reg_3_ ( .clear(DP_reg_pipe11_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe01[3]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe11[3]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe11_Q_reg_4_ ( .clear(DP_reg_pipe11_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe01[4]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe11[4]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe11_Q_reg_5_ ( .clear(DP_reg_pipe11_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe01[5]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe11[5]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe11_Q_reg_6_ ( .clear(DP_reg_pipe11_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe01[6]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe11[6]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe11_Q_reg_7_ ( .clear(DP_reg_pipe11_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe01[7]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe11[7]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe11_Q_reg_8_ ( .clear(DP_reg_pipe11_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe01[8]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe11[8]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe11_Q_reg_9_ ( .clear(DP_reg_pipe11_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe01[9]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe11[9]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe11_Q_reg_10_ ( .clear(DP_reg_pipe11_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe01[10]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe11[10]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe11_Q_reg_11_ ( .clear(DP_reg_pipe11_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe01[11]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe11[11]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe11_Q_reg_12_ ( .clear(DP_reg_pipe11_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe01[12]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe11[12]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe11_Q_reg_13_ ( .clear(DP_reg_pipe11_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe01[13]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe11[13]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe11_Q_reg_14_ ( .clear(DP_reg_pipe11_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe01[14]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe11[14]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe11_Q_reg_15_ ( .clear(DP_reg_pipe11_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe01[15]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe11[15]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe11_Q_reg_16_ ( .clear(DP_reg_pipe11_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe01[16]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe11[16]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe11_Q_reg_17_ ( .clear(DP_reg_pipe11_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe01[17]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe11[17]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe11_Q_reg_18_ ( .clear(DP_reg_pipe11_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe01[18]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe11[18]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe11_Q_reg_19_ ( .clear(DP_reg_pipe11_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe01[19]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe11[19]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe11_Q_reg_20_ ( .clear(DP_reg_pipe11_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe01[20]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe11[20]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe11_Q_reg_21_ ( .clear(DP_reg_pipe11_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe01[21]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe11[21]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe11_Q_reg_22_ ( .clear(DP_reg_pipe11_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe01[22]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe11[22]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe11_Q_reg_23_ ( .clear(DP_reg_pipe11_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe01[23]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe11[23]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  GTECH_NOT DP_reg_pipe12_I_0 ( .A(rst_n), .Z(DP_reg_pipe12_N0) );
  \**SEQGEN**  DP_reg_pipe12_Q_reg_0_ ( .clear(DP_reg_pipe12_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe02[0]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe12[0]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe12_Q_reg_1_ ( .clear(DP_reg_pipe12_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe02[1]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe12[1]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe12_Q_reg_2_ ( .clear(DP_reg_pipe12_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe02[2]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe12[2]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe12_Q_reg_3_ ( .clear(DP_reg_pipe12_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe02[3]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe12[3]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe12_Q_reg_4_ ( .clear(DP_reg_pipe12_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe02[4]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe12[4]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe12_Q_reg_5_ ( .clear(DP_reg_pipe12_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe02[5]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe12[5]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe12_Q_reg_6_ ( .clear(DP_reg_pipe12_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe02[6]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe12[6]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe12_Q_reg_7_ ( .clear(DP_reg_pipe12_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe02[7]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe12[7]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe12_Q_reg_8_ ( .clear(DP_reg_pipe12_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe02[8]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe12[8]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe12_Q_reg_9_ ( .clear(DP_reg_pipe12_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe02[9]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe12[9]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe12_Q_reg_10_ ( .clear(DP_reg_pipe12_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe02[10]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe12[10]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe12_Q_reg_11_ ( .clear(DP_reg_pipe12_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe02[11]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe12[11]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe12_Q_reg_12_ ( .clear(DP_reg_pipe12_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe02[12]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe12[12]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe12_Q_reg_13_ ( .clear(DP_reg_pipe12_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe02[13]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe12[13]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe12_Q_reg_14_ ( .clear(DP_reg_pipe12_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe02[14]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe12[14]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe12_Q_reg_15_ ( .clear(DP_reg_pipe12_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe02[15]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe12[15]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe12_Q_reg_16_ ( .clear(DP_reg_pipe12_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe02[16]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe12[16]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe12_Q_reg_17_ ( .clear(DP_reg_pipe12_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe02[17]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe12[17]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe12_Q_reg_18_ ( .clear(DP_reg_pipe12_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe02[18]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe12[18]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe12_Q_reg_19_ ( .clear(DP_reg_pipe12_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe02[19]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe12[19]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe12_Q_reg_20_ ( .clear(DP_reg_pipe12_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe02[20]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe12[20]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe12_Q_reg_21_ ( .clear(DP_reg_pipe12_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe02[21]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe12[21]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe12_Q_reg_22_ ( .clear(DP_reg_pipe12_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe02[22]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe12[22]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe12_Q_reg_23_ ( .clear(DP_reg_pipe12_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe02[23]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe12[23]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  GTECH_NOT DP_reg_pipe13_I_0 ( .A(rst_n), .Z(DP_reg_pipe13_N0) );
  \**SEQGEN**  DP_reg_pipe13_Q_reg_0_ ( .clear(DP_reg_pipe13_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe03[0]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe13[0]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe13_Q_reg_1_ ( .clear(DP_reg_pipe13_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe03[1]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe13[1]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe13_Q_reg_2_ ( .clear(DP_reg_pipe13_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe03[2]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe13[2]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe13_Q_reg_3_ ( .clear(DP_reg_pipe13_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe03[3]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe13[3]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe13_Q_reg_4_ ( .clear(DP_reg_pipe13_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe03[4]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe13[4]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe13_Q_reg_5_ ( .clear(DP_reg_pipe13_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe03[5]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe13[5]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe13_Q_reg_6_ ( .clear(DP_reg_pipe13_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe03[6]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe13[6]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe13_Q_reg_7_ ( .clear(DP_reg_pipe13_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe03[7]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe13[7]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe13_Q_reg_8_ ( .clear(DP_reg_pipe13_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe03[8]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe13[8]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe13_Q_reg_9_ ( .clear(DP_reg_pipe13_N0), .preset(1'b0), .next_state(DP_pipe0_coeff_pipe03[9]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(DP_pipe13[9]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe13_Q_reg_10_ ( .clear(DP_reg_pipe13_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe03[10]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe13[10]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe13_Q_reg_11_ ( .clear(DP_reg_pipe13_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe03[11]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe13[11]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe13_Q_reg_12_ ( .clear(DP_reg_pipe13_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe03[12]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe13[12]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe13_Q_reg_13_ ( .clear(DP_reg_pipe13_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe03[13]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe13[13]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe13_Q_reg_14_ ( .clear(DP_reg_pipe13_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe03[14]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe13[14]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe13_Q_reg_15_ ( .clear(DP_reg_pipe13_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe03[15]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe13[15]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe13_Q_reg_16_ ( .clear(DP_reg_pipe13_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe03[16]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe13[16]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe13_Q_reg_17_ ( .clear(DP_reg_pipe13_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe03[17]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe13[17]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe13_Q_reg_18_ ( .clear(DP_reg_pipe13_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe03[18]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe13[18]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe13_Q_reg_19_ ( .clear(DP_reg_pipe13_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe03[19]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe13[19]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe13_Q_reg_20_ ( .clear(DP_reg_pipe13_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe03[20]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe13[20]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe13_Q_reg_21_ ( .clear(DP_reg_pipe13_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe03[21]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe13[21]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe13_Q_reg_22_ ( .clear(DP_reg_pipe13_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe03[22]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe13[22]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DP_reg_pipe13_Q_reg_23_ ( .clear(DP_reg_pipe13_N0), .preset(
        1'b0), .next_state(DP_pipe0_coeff_pipe03[23]), .clocked_on(clk), 
        .data_in(1'b0), .enable(1'b0), .Q(DP_pipe13[23]), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  GTECH_NOT DP_reg_out_I_0 ( .A(rst_n), .Z(DP_reg_out_N0) );
  \**SEQGEN**  DP_reg_out_Q_reg_0_ ( .clear(DP_reg_out_N0), .preset(1'b0), 
        .next_state(DP_y_out[0]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(dOut[0]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(delayed_controls_2__0_) );
  \**SEQGEN**  DP_reg_out_Q_reg_1_ ( .clear(DP_reg_out_N0), .preset(1'b0), 
        .next_state(DP_y_out[1]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(dOut[1]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(delayed_controls_2__0_) );
  \**SEQGEN**  DP_reg_out_Q_reg_2_ ( .clear(DP_reg_out_N0), .preset(1'b0), 
        .next_state(DP_y_out[2]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(dOut[2]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(delayed_controls_2__0_) );
  \**SEQGEN**  DP_reg_out_Q_reg_3_ ( .clear(DP_reg_out_N0), .preset(1'b0), 
        .next_state(DP_y_out[3]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(dOut[3]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(delayed_controls_2__0_) );
  \**SEQGEN**  DP_reg_out_Q_reg_4_ ( .clear(DP_reg_out_N0), .preset(1'b0), 
        .next_state(DP_y_out[4]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(dOut[4]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(delayed_controls_2__0_) );
  \**SEQGEN**  DP_reg_out_Q_reg_5_ ( .clear(DP_reg_out_N0), .preset(1'b0), 
        .next_state(DP_y_out[5]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(dOut[5]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(delayed_controls_2__0_) );
  \**SEQGEN**  DP_reg_out_Q_reg_6_ ( .clear(DP_reg_out_N0), .preset(1'b0), 
        .next_state(DP_y_out[6]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(dOut[6]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(delayed_controls_2__0_) );
  \**SEQGEN**  DP_reg_out_Q_reg_7_ ( .clear(DP_reg_out_N0), .preset(1'b0), 
        .next_state(DP_y_out[7]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(dOut[7]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(delayed_controls_2__0_) );
  \**SEQGEN**  DP_reg_out_Q_reg_8_ ( .clear(DP_reg_out_N0), .preset(1'b0), 
        .next_state(DP_y_out[8]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(dOut[8]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(delayed_controls_2__0_) );
  \**SEQGEN**  DP_reg_out_Q_reg_9_ ( .clear(DP_reg_out_N0), .preset(1'b0), 
        .next_state(DP_y_out[9]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(dOut[9]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(delayed_controls_2__0_) );
  \**SEQGEN**  DP_reg_out_Q_reg_10_ ( .clear(DP_reg_out_N0), .preset(1'b0), 
        .next_state(DP_y_out[10]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(dOut[10]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(delayed_controls_2__0_) );
  \**SEQGEN**  DP_reg_out_Q_reg_11_ ( .clear(DP_reg_out_N0), .preset(1'b0), 
        .next_state(DP_y_out[11]), .clocked_on(clk), .data_in(1'b0), .enable(
        1'b0), .Q(dOut[11]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(delayed_controls_2__0_) );
  GTECH_AND2 CU_C91 ( .A(CU_presentState_1_), .B(CU_presentState_0_), .Z(
        CU_N11) );
  GTECH_OR2 CU_C89 ( .A(CU_N13), .B(CU_presentState_0_), .Z(CU_N18) );
  GTECH_NOT CU_I_7 ( .A(CU_N18), .Z(CU_N10) );
  GTECH_OR2 CU_C86 ( .A(CU_presentState_1_), .B(CU_N14), .Z(CU_N17) );
  GTECH_NOT CU_I_6 ( .A(CU_N17), .Z(CU_N9) );
  GTECH_NOT CU_I_5 ( .A(vIn), .Z(CU_N8) );
  GTECH_AND2 CU_C82 ( .A(CU_presentState_1_), .B(CU_presentState_0_), .Z(CU_N7) );
  GTECH_OR2 CU_C80 ( .A(CU_N13), .B(CU_presentState_0_), .Z(CU_N16) );
  GTECH_NOT CU_I_4 ( .A(CU_N16), .Z(CU_N6) );
  GTECH_OR2 CU_C77 ( .A(CU_presentState_1_), .B(CU_N14), .Z(CU_N15) );
  GTECH_NOT CU_I_3 ( .A(CU_N15), .Z(CU_N5) );
  GTECH_NOT CU_I_2 ( .A(CU_presentState_0_), .Z(CU_N14) );
  GTECH_NOT CU_I_1 ( .A(CU_presentState_1_), .Z(CU_N13) );
  GTECH_AND2 CU_C73 ( .A(CU_N13), .B(CU_N14), .Z(CU_N4) );
  GTECH_BUF CU_B_3 ( .A(CU_N7), .Z(CU_N3) );
  GTECH_BUF CU_B_2 ( .A(CU_N6), .Z(CU_N2) );
  GTECH_BUF CU_B_1 ( .A(CU_N5), .Z(CU_N1) );
  GTECH_BUF CU_B_0 ( .A(CU_N4), .Z(CU_N0) );
  SELECT_OP CU_C70 ( .DATA1(vIn), .DATA2(CU_N8), .DATA3(CU_N8), .DATA4(vIn), 
        .CONTROL1(CU_N0), .CONTROL2(CU_N1), .CONTROL3(CU_N2), .CONTROL4(CU_N3), 
        .Z(CU_nextState[0]) );
  GTECH_OR2 CU_C68 ( .A(CU_N10), .B(CU_N11), .Z(delayed_controls_0__1_) );
  GTECH_OR2 CU_C62 ( .A(CU_N9), .B(CU_N10), .Z(sw_regs_en_int) );
  GTECH_OR2 CU_C59 ( .A(CU_N5), .B(CU_N6), .Z(CU_nextState[1]) );
  GTECH_NOT CU_I_0 ( .A(rst_n), .Z(CU_N12) );
  \**SEQGEN**  CU_presentState_reg_0_ ( .clear(CU_N12), .preset(1'b0), 
        .next_state(CU_nextState[0]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(CU_presentState_0_), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  CU_presentState_reg_1_ ( .clear(CU_N12), .preset(1'b0), 
        .next_state(CU_nextState[1]), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(CU_presentState_1_), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  GTECH_NOT reg_delay_0_I_0 ( .A(rst_n), .Z(reg_delay_0_N0) );
  \**SEQGEN**  reg_delay_0_Q_reg_0_ ( .clear(reg_delay_0_N0), .preset(1'b0), 
        .next_state(delayed_controls_0__1_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(delayed_controls_1__1_), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  reg_delay_0_Q_reg_1_ ( .clear(reg_delay_0_N0), .preset(1'b0), 
        .next_state(sw_regs_en_int), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(delayed_controls_1__0_), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  GTECH_NOT reg_delay_1_I_0 ( .A(rst_n), .Z(reg_delay_1_N0) );
  \**SEQGEN**  reg_delay_1_Q_reg_0_ ( .clear(reg_delay_1_N0), .preset(1'b0), 
        .next_state(delayed_controls_1__1_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vOut), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  reg_delay_1_Q_reg_1_ ( .clear(reg_delay_1_N0), .preset(1'b0), 
        .next_state(delayed_controls_1__0_), .clocked_on(clk), .data_in(1'b0), 
        .enable(1'b0), .Q(delayed_controls_2__0_), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
endmodule

