----------------------------- 
-- COLUMN 0
----------------------------- 
-- full adder c0, number 0
0_FA_0: fullAdder
	port map (
		i0 => grid5(0)(0),
		i1 => grid5(1)(0),
		ci => grid5(2)(0),
		s => grid4(0)(0),
		co => grid4(0)(1) );

-- full adder c0, number 1
0_FA_1: fullAdder
	port map (
		i0 => grid5(3)(0),
		i1 => grid5(4)(0),
		ci => grid5(5)(0),
		s => grid4(1)(0),
		co => grid4(1)(1) );

-- half adder c0, number 0
0_HA_0: halfAdder
	port map (
		i0 => grid5(6)(0),
		i1 => grid5(7)(0),
		s => grid4(2)(0),
		co => grid4(2)(1) );

-- move the other elements of the column
grid4(3)(0) <= grid5(8)(0);
grid4(4)(0) <= grid5(9)(0);
grid4(5)(0) <= grid5(10)(0);
grid4(6)(0) <= grid5(11)(0);

----------------------------- 
-- COLUMN 1
----------------------------- 
-- full adder c1, number 0
1_FA_0: fullAdder
	port map (
		i0 => grid5(0)(1),
		i1 => grid5(1)(1),
		ci => grid5(2)(1),
		s => grid4(3)(1),
		co => grid4(0)(2) );

-- full adder c1, number 1
1_FA_1: fullAdder
	port map (
		i0 => grid5(3)(1),
		i1 => grid5(4)(1),
		ci => grid5(5)(1),
		s => grid4(4)(1),
		co => grid4(1)(2) );

-- half adder c1, number 0
1_HA_0: halfAdder
	port map (
		i0 => grid5(6)(1),
		i1 => grid5(7)(1),
		s => grid4(5)(1),
		co => grid4(2)(2) );

-- move the other elements of the column
grid4(6)(1) <= grid5(8)(1);
grid4(7)(1) <= grid5(9)(1);
grid4(8)(1) <= grid5(10)(1);
grid4(9)(1) <= grid5(11)(1);

----------------------------- 
-- COLUMN 2
----------------------------- 
-- full adder c2, number 0
2_FA_0: fullAdder
	port map (
		i0 => grid5(0)(2),
		i1 => grid5(1)(2),
		ci => grid5(2)(2),
		s => grid4(3)(2),
		co => grid4(0)(3) );

-- full adder c2, number 1
2_FA_1: fullAdder
	port map (
		i0 => grid5(3)(2),
		i1 => grid5(4)(2),
		ci => grid5(5)(2),
		s => grid4(4)(2),
		co => grid4(1)(3) );

-- half adder c2, number 0
2_HA_0: halfAdder
	port map (
		i0 => grid5(6)(2),
		i1 => grid5(7)(2),
		s => grid4(5)(2),
		co => grid4(2)(3) );

-- move the other elements of the column
grid4(6)(2) <= grid5(8)(2);
grid4(7)(2) <= grid5(9)(2);
grid4(8)(2) <= grid5(10)(2);
grid4(9)(2) <= grid5(11)(2);

----------------------------- 
-- COLUMN 3
----------------------------- 
-- full adder c3, number 0
3_FA_0: fullAdder
	port map (
		i0 => grid5(0)(3),
		i1 => grid5(1)(3),
		ci => grid5(2)(3),
		s => grid4(3)(3),
		co => grid4(0)(4) );

-- full adder c3, number 1
3_FA_1: fullAdder
	port map (
		i0 => grid5(3)(3),
		i1 => grid5(4)(3),
		ci => grid5(5)(3),
		s => grid4(4)(3),
		co => grid4(1)(4) );

-- half adder c3, number 0
3_HA_0: halfAdder
	port map (
		i0 => grid5(6)(3),
		i1 => grid5(7)(3),
		s => grid4(5)(3),
		co => grid4(2)(4) );

-- move the other elements of the column
grid4(6)(3) <= grid5(8)(3);
grid4(7)(3) <= grid5(9)(3);
grid4(8)(3) <= grid5(10)(3);
grid4(9)(3) <= grid5(11)(3);

----------------------------- 
-- COLUMN 4
----------------------------- 
-- full adder c4, number 0
4_FA_0: fullAdder
	port map (
		i0 => grid5(0)(4),
		i1 => grid5(1)(4),
		ci => grid5(2)(4),
		s => grid4(3)(4),
		co => grid4(0)(5) );

-- full adder c4, number 1
4_FA_1: fullAdder
	port map (
		i0 => grid5(3)(4),
		i1 => grid5(4)(4),
		ci => grid5(5)(4),
		s => grid4(4)(4),
		co => grid4(1)(5) );

-- half adder c4, number 0
4_HA_0: halfAdder
	port map (
		i0 => grid5(6)(4),
		i1 => grid5(7)(4),
		s => grid4(5)(4),
		co => grid4(2)(5) );

-- move the other elements of the column
grid4(6)(4) <= grid5(8)(4);
grid4(7)(4) <= grid5(9)(4);
grid4(8)(4) <= grid5(10)(4);
grid4(9)(4) <= grid5(11)(4);

----------------------------- 
-- COLUMN 5
----------------------------- 
-- full adder c5, number 0
5_FA_0: fullAdder
	port map (
		i0 => grid5(0)(5),
		i1 => grid5(1)(5),
		ci => grid5(2)(5),
		s => grid4(3)(5),
		co => grid4(0)(6) );

-- full adder c5, number 1
5_FA_1: fullAdder
	port map (
		i0 => grid5(3)(5),
		i1 => grid5(4)(5),
		ci => grid5(5)(5),
		s => grid4(4)(5),
		co => grid4(1)(6) );

-- half adder c5, number 0
5_HA_0: halfAdder
	port map (
		i0 => grid5(6)(5),
		i1 => grid5(7)(5),
		s => grid4(5)(5),
		co => grid4(2)(6) );

-- move the other elements of the column
grid4(6)(5) <= grid5(8)(5);
grid4(7)(5) <= grid5(9)(5);
grid4(8)(5) <= grid5(10)(5);
grid4(9)(5) <= grid5(11)(5);

----------------------------- 
-- COLUMN 6
----------------------------- 
-- full adder c6, number 0
6_FA_0: fullAdder
	port map (
		i0 => grid5(0)(6),
		i1 => grid5(1)(6),
		ci => grid5(2)(6),
		s => grid4(3)(6),
		co => grid4(0)(7) );

-- full adder c6, number 1
6_FA_1: fullAdder
	port map (
		i0 => grid5(3)(6),
		i1 => grid5(4)(6),
		ci => grid5(5)(6),
		s => grid4(4)(6),
		co => grid4(1)(7) );

-- half adder c6, number 0
6_HA_0: halfAdder
	port map (
		i0 => grid5(6)(6),
		i1 => grid5(7)(6),
		s => grid4(5)(6),
		co => grid4(2)(7) );

-- move the other elements of the column
grid4(6)(6) <= grid5(8)(6);
grid4(7)(6) <= grid5(9)(6);
grid4(8)(6) <= grid5(10)(6);
grid4(9)(6) <= grid5(11)(6);

----------------------------- 
-- COLUMN 7
----------------------------- 
-- full adder c7, number 0
7_FA_0: fullAdder
	port map (
		i0 => grid5(0)(7),
		i1 => grid5(1)(7),
		ci => grid5(2)(7),
		s => grid4(3)(7),
		co => grid4(0)(8) );

-- full adder c7, number 1
7_FA_1: fullAdder
	port map (
		i0 => grid5(3)(7),
		i1 => grid5(4)(7),
		ci => grid5(5)(7),
		s => grid4(4)(7),
		co => grid4(1)(8) );

-- half adder c7, number 0
7_HA_0: halfAdder
	port map (
		i0 => grid5(6)(7),
		i1 => grid5(7)(7),
		s => grid4(5)(7),
		co => grid4(2)(8) );

-- move the other elements of the column
grid4(6)(7) <= grid5(8)(7);
grid4(7)(7) <= grid5(9)(7);
grid4(8)(7) <= grid5(10)(7);
grid4(9)(7) <= grid5(11)(7);

----------------------------- 
-- COLUMN 8
----------------------------- 
-- full adder c8, number 0
8_FA_0: fullAdder
	port map (
		i0 => grid5(0)(8),
		i1 => grid5(1)(8),
		ci => grid5(2)(8),
		s => grid4(3)(8),
		co => grid4(0)(9) );

-- full adder c8, number 1
8_FA_1: fullAdder
	port map (
		i0 => grid5(3)(8),
		i1 => grid5(4)(8),
		ci => grid5(5)(8),
		s => grid4(4)(8),
		co => grid4(1)(9) );

-- half adder c8, number 0
8_HA_0: halfAdder
	port map (
		i0 => grid5(6)(8),
		i1 => grid5(7)(8),
		s => grid4(5)(8),
		co => grid4(2)(9) );

-- move the other elements of the column
grid4(6)(8) <= grid5(8)(8);
grid4(7)(8) <= grid5(9)(8);
grid4(8)(8) <= grid5(10)(8);
grid4(9)(8) <= grid5(11)(8);

----------------------------- 
-- COLUMN 9
----------------------------- 
-- full adder c9, number 0
9_FA_0: fullAdder
	port map (
		i0 => grid5(0)(9),
		i1 => grid5(1)(9),
		ci => grid5(2)(9),
		s => grid4(3)(9),
		co => grid4(0)(10) );

-- full adder c9, number 1
9_FA_1: fullAdder
	port map (
		i0 => grid5(3)(9),
		i1 => grid5(4)(9),
		ci => grid5(5)(9),
		s => grid4(4)(9),
		co => grid4(1)(10) );

-- half adder c9, number 0
9_HA_0: halfAdder
	port map (
		i0 => grid5(6)(9),
		i1 => grid5(7)(9),
		s => grid4(5)(9),
		co => grid4(2)(10) );

-- move the other elements of the column
grid4(6)(9) <= grid5(8)(9);
grid4(7)(9) <= grid5(9)(9);
grid4(8)(9) <= grid5(10)(9);
grid4(9)(9) <= grid5(11)(9);

----------------------------- 
-- COLUMN 10
----------------------------- 
-- full adder c10, number 0
10_FA_0: fullAdder
	port map (
		i0 => grid5(0)(10),
		i1 => grid5(1)(10),
		ci => grid5(2)(10),
		s => grid4(3)(10),
		co => grid4(0)(11) );

-- full adder c10, number 1
10_FA_1: fullAdder
	port map (
		i0 => grid5(3)(10),
		i1 => grid5(4)(10),
		ci => grid5(5)(10),
		s => grid4(4)(10),
		co => grid4(1)(11) );

-- half adder c10, number 0
10_HA_0: halfAdder
	port map (
		i0 => grid5(6)(10),
		i1 => grid5(7)(10),
		s => grid4(5)(10),
		co => grid4(2)(11) );

-- move the other elements of the column
grid4(6)(10) <= grid5(8)(10);
grid4(7)(10) <= grid5(9)(10);
grid4(8)(10) <= grid5(10)(10);
grid4(9)(10) <= grid5(11)(10);

----------------------------- 
-- COLUMN 11
----------------------------- 
-- full adder c11, number 0
11_FA_0: fullAdder
	port map (
		i0 => grid5(0)(11),
		i1 => grid5(1)(11),
		ci => grid5(2)(11),
		s => grid4(3)(11),
		co => grid4(0)(12) );

-- full adder c11, number 1
11_FA_1: fullAdder
	port map (
		i0 => grid5(3)(11),
		i1 => grid5(4)(11),
		ci => grid5(5)(11),
		s => grid4(4)(11),
		co => grid4(1)(12) );

-- half adder c11, number 0
11_HA_0: halfAdder
	port map (
		i0 => grid5(6)(11),
		i1 => grid5(7)(11),
		s => grid4(5)(11),
		co => grid4(2)(12) );

-- move the other elements of the column
grid4(6)(11) <= grid5(8)(11);
grid4(7)(11) <= grid5(9)(11);
grid4(8)(11) <= grid5(10)(11);
grid4(9)(11) <= grid5(11)(11);

----------------------------- 
-- COLUMN 12
----------------------------- 
-- full adder c12, number 0
12_FA_0: fullAdder
	port map (
		i0 => grid5(0)(12),
		i1 => grid5(1)(12),
		ci => grid5(2)(12),
		s => grid4(3)(12),
		co => grid4(0)(13) );

-- full adder c12, number 1
12_FA_1: fullAdder
	port map (
		i0 => grid5(3)(12),
		i1 => grid5(4)(12),
		ci => grid5(5)(12),
		s => grid4(4)(12),
		co => grid4(1)(13) );

-- half adder c12, number 0
12_HA_0: halfAdder
	port map (
		i0 => grid5(6)(12),
		i1 => grid5(7)(12),
		s => grid4(5)(12),
		co => grid4(2)(13) );

-- move the other elements of the column
grid4(6)(12) <= grid5(8)(12);
grid4(7)(12) <= grid5(9)(12);
grid4(8)(12) <= grid5(10)(12);
grid4(9)(12) <= grid5(11)(12);

----------------------------- 
-- COLUMN 13
----------------------------- 
-- full adder c13, number 0
13_FA_0: fullAdder
	port map (
		i0 => grid5(0)(13),
		i1 => grid5(1)(13),
		ci => grid5(2)(13),
		s => grid4(3)(13),
		co => grid4(0)(14) );

-- full adder c13, number 1
13_FA_1: fullAdder
	port map (
		i0 => grid5(3)(13),
		i1 => grid5(4)(13),
		ci => grid5(5)(13),
		s => grid4(4)(13),
		co => grid4(1)(14) );

-- half adder c13, number 0
13_HA_0: halfAdder
	port map (
		i0 => grid5(6)(13),
		i1 => grid5(7)(13),
		s => grid4(5)(13),
		co => grid4(2)(14) );

-- move the other elements of the column
grid4(6)(13) <= grid5(8)(13);
grid4(7)(13) <= grid5(9)(13);
grid4(8)(13) <= grid5(10)(13);
grid4(9)(13) <= grid5(11)(13);

----------------------------- 
-- COLUMN 14
----------------------------- 
-- full adder c14, number 0
14_FA_0: fullAdder
	port map (
		i0 => grid5(0)(14),
		i1 => grid5(1)(14),
		ci => grid5(2)(14),
		s => grid4(3)(14),
		co => grid4(0)(15) );

-- full adder c14, number 1
14_FA_1: fullAdder
	port map (
		i0 => grid5(3)(14),
		i1 => grid5(4)(14),
		ci => grid5(5)(14),
		s => grid4(4)(14),
		co => grid4(1)(15) );

-- half adder c14, number 0
14_HA_0: halfAdder
	port map (
		i0 => grid5(6)(14),
		i1 => grid5(7)(14),
		s => grid4(5)(14),
		co => grid4(2)(15) );

-- move the other elements of the column
grid4(6)(14) <= grid5(8)(14);
grid4(7)(14) <= grid5(9)(14);
grid4(8)(14) <= grid5(10)(14);
grid4(9)(14) <= grid5(11)(14);

----------------------------- 
-- COLUMN 15
----------------------------- 
-- full adder c15, number 0
15_FA_0: fullAdder
	port map (
		i0 => grid5(0)(15),
		i1 => grid5(1)(15),
		ci => grid5(2)(15),
		s => grid4(3)(15),
		co => grid4(0)(16) );

-- full adder c15, number 1
15_FA_1: fullAdder
	port map (
		i0 => grid5(3)(15),
		i1 => grid5(4)(15),
		ci => grid5(5)(15),
		s => grid4(4)(15),
		co => grid4(1)(16) );

-- half adder c15, number 0
15_HA_0: halfAdder
	port map (
		i0 => grid5(6)(15),
		i1 => grid5(7)(15),
		s => grid4(5)(15),
		co => grid4(2)(16) );

-- move the other elements of the column
grid4(6)(15) <= grid5(8)(15);
grid4(7)(15) <= grid5(9)(15);
grid4(8)(15) <= grid5(10)(15);
grid4(9)(15) <= grid5(11)(15);

----------------------------- 
-- COLUMN 16
----------------------------- 
-- full adder c16, number 0
16_FA_0: fullAdder
	port map (
		i0 => grid5(0)(16),
		i1 => grid5(1)(16),
		ci => grid5(2)(16),
		s => grid4(3)(16),
		co => grid4(0)(17) );

-- full adder c16, number 1
16_FA_1: fullAdder
	port map (
		i0 => grid5(3)(16),
		i1 => grid5(4)(16),
		ci => grid5(5)(16),
		s => grid4(4)(16),
		co => grid4(1)(17) );

-- half adder c16, number 0
16_HA_0: halfAdder
	port map (
		i0 => grid5(6)(16),
		i1 => grid5(7)(16),
		s => grid4(5)(16),
		co => grid4(2)(17) );

-- move the other elements of the column
grid4(6)(16) <= grid5(8)(16);
grid4(7)(16) <= grid5(9)(16);
grid4(8)(16) <= grid5(10)(16);
grid4(9)(16) <= grid5(11)(16);

----------------------------- 
-- COLUMN 17
----------------------------- 
-- full adder c17, number 0
17_FA_0: fullAdder
	port map (
		i0 => grid5(0)(17),
		i1 => grid5(1)(17),
		ci => grid5(2)(17),
		s => grid4(3)(17),
		co => grid4(0)(18) );

-- full adder c17, number 1
17_FA_1: fullAdder
	port map (
		i0 => grid5(3)(17),
		i1 => grid5(4)(17),
		ci => grid5(5)(17),
		s => grid4(4)(17),
		co => grid4(1)(18) );

-- half adder c17, number 0
17_HA_0: halfAdder
	port map (
		i0 => grid5(6)(17),
		i1 => grid5(7)(17),
		s => grid4(5)(17),
		co => grid4(2)(18) );

-- move the other elements of the column
grid4(6)(17) <= grid5(8)(17);
grid4(7)(17) <= grid5(9)(17);
grid4(8)(17) <= grid5(10)(17);
grid4(9)(17) <= grid5(11)(17);

----------------------------- 
-- COLUMN 18
----------------------------- 
-- full adder c18, number 0
18_FA_0: fullAdder
	port map (
		i0 => grid5(0)(18),
		i1 => grid5(1)(18),
		ci => grid5(2)(18),
		s => grid4(3)(18),
		co => grid4(0)(19) );

-- full adder c18, number 1
18_FA_1: fullAdder
	port map (
		i0 => grid5(3)(18),
		i1 => grid5(4)(18),
		ci => grid5(5)(18),
		s => grid4(4)(18),
		co => grid4(1)(19) );

-- half adder c18, number 0
18_HA_0: halfAdder
	port map (
		i0 => grid5(6)(18),
		i1 => grid5(7)(18),
		s => grid4(5)(18),
		co => grid4(2)(19) );

-- move the other elements of the column
grid4(6)(18) <= grid5(8)(18);
grid4(7)(18) <= grid5(9)(18);
grid4(8)(18) <= grid5(10)(18);
grid4(9)(18) <= grid5(11)(18);

----------------------------- 
-- COLUMN 19
----------------------------- 
-- full adder c19, number 0
19_FA_0: fullAdder
	port map (
		i0 => grid5(0)(19),
		i1 => grid5(1)(19),
		ci => grid5(2)(19),
		s => grid4(3)(19),
		co => grid4(0)(20) );

-- full adder c19, number 1
19_FA_1: fullAdder
	port map (
		i0 => grid5(3)(19),
		i1 => grid5(4)(19),
		ci => grid5(5)(19),
		s => grid4(4)(19),
		co => grid4(1)(20) );

-- half adder c19, number 0
19_HA_0: halfAdder
	port map (
		i0 => grid5(6)(19),
		i1 => grid5(7)(19),
		s => grid4(5)(19),
		co => grid4(2)(20) );

-- move the other elements of the column
grid4(6)(19) <= grid5(8)(19);
grid4(7)(19) <= grid5(9)(19);
grid4(8)(19) <= grid5(10)(19);
grid4(9)(19) <= grid5(11)(19);

----------------------------- 
-- COLUMN 20
----------------------------- 
-- full adder c20, number 0
20_FA_0: fullAdder
	port map (
		i0 => grid5(0)(20),
		i1 => grid5(1)(20),
		ci => grid5(2)(20),
		s => grid4(3)(20),
		co => grid4(0)(21) );

-- full adder c20, number 1
20_FA_1: fullAdder
	port map (
		i0 => grid5(3)(20),
		i1 => grid5(4)(20),
		ci => grid5(5)(20),
		s => grid4(4)(20),
		co => grid4(1)(21) );

-- half adder c20, number 0
20_HA_0: halfAdder
	port map (
		i0 => grid5(6)(20),
		i1 => grid5(7)(20),
		s => grid4(5)(20),
		co => grid4(2)(21) );

-- move the other elements of the column
grid4(6)(20) <= grid5(8)(20);
grid4(7)(20) <= grid5(9)(20);
grid4(8)(20) <= grid5(10)(20);
grid4(9)(20) <= grid5(11)(20);

----------------------------- 
-- COLUMN 21
----------------------------- 
-- full adder c21, number 0
21_FA_0: fullAdder
	port map (
		i0 => grid5(0)(21),
		i1 => grid5(1)(21),
		ci => grid5(2)(21),
		s => grid4(3)(21),
		co => grid4(0)(22) );

-- full adder c21, number 1
21_FA_1: fullAdder
	port map (
		i0 => grid5(3)(21),
		i1 => grid5(4)(21),
		ci => grid5(5)(21),
		s => grid4(4)(21),
		co => grid4(1)(22) );

-- half adder c21, number 0
21_HA_0: halfAdder
	port map (
		i0 => grid5(6)(21),
		i1 => grid5(7)(21),
		s => grid4(5)(21),
		co => grid4(2)(22) );

-- move the other elements of the column
grid4(6)(21) <= grid5(8)(21);
grid4(7)(21) <= grid5(9)(21);
grid4(8)(21) <= grid5(10)(21);
grid4(9)(21) <= grid5(11)(21);

----------------------------- 
-- COLUMN 22
----------------------------- 
-- full adder c22, number 0
22_FA_0: fullAdder
	port map (
		i0 => grid5(0)(22),
		i1 => grid5(1)(22),
		ci => grid5(2)(22),
		s => grid4(3)(22),
		co => grid4(0)(23) );

-- full adder c22, number 1
22_FA_1: fullAdder
	port map (
		i0 => grid5(3)(22),
		i1 => grid5(4)(22),
		ci => grid5(5)(22),
		s => grid4(4)(22),
		co => grid4(1)(23) );

-- half adder c22, number 0
22_HA_0: halfAdder
	port map (
		i0 => grid5(6)(22),
		i1 => grid5(7)(22),
		s => grid4(5)(22),
		co => grid4(2)(23) );

-- move the other elements of the column
grid4(6)(22) <= grid5(8)(22);
grid4(7)(22) <= grid5(9)(22);
grid4(8)(22) <= grid5(10)(22);
grid4(9)(22) <= grid5(11)(22);

----------------------------- 
-- COLUMN 23
----------------------------- 
-- full adder c23, number 0
23_FA_0: fullAdder
	port map (
		i0 => grid5(0)(23),
		i1 => grid5(1)(23),
		ci => grid5(2)(23),
		s => grid4(3)(23),
		co => grid4(0)(24) );

-- full adder c23, number 1
23_FA_1: fullAdder
	port map (
		i0 => grid5(3)(23),
		i1 => grid5(4)(23),
		ci => grid5(5)(23),
		s => grid4(4)(23),
		co => grid4(1)(24) );

-- half adder c23, number 0
23_HA_0: halfAdder
	port map (
		i0 => grid5(6)(23),
		i1 => grid5(7)(23),
		s => grid4(5)(23),
		co => grid4(2)(24) );

-- move the other elements of the column
grid4(6)(23) <= grid5(8)(23);
grid4(7)(23) <= grid5(9)(23);
grid4(8)(23) <= grid5(10)(23);
grid4(9)(23) <= grid5(11)(23);

----------------------------- 
-- COLUMN 24
----------------------------- 
-- full adder c24, number 0
24_FA_0: fullAdder
	port map (
		i0 => grid5(0)(24),
		i1 => grid5(1)(24),
		ci => grid5(2)(24),
		s => grid4(3)(24),
		co => grid4(0)(25) );

-- full adder c24, number 1
24_FA_1: fullAdder
	port map (
		i0 => grid5(3)(24),
		i1 => grid5(4)(24),
		ci => grid5(5)(24),
		s => grid4(4)(24),
		co => grid4(1)(25) );

-- half adder c24, number 0
24_HA_0: halfAdder
	port map (
		i0 => grid5(6)(24),
		i1 => grid5(7)(24),
		s => grid4(5)(24),
		co => grid4(2)(25) );

-- move the other elements of the column
grid4(6)(24) <= grid5(8)(24);
grid4(7)(24) <= grid5(9)(24);
grid4(8)(24) <= grid5(10)(24);
grid4(9)(24) <= grid5(11)(24);

----------------------------- 
-- COLUMN 25
----------------------------- 
-- full adder c25, number 0
25_FA_0: fullAdder
	port map (
		i0 => grid5(0)(25),
		i1 => grid5(1)(25),
		ci => grid5(2)(25),
		s => grid4(3)(25),
		co => grid4(0)(26) );

-- full adder c25, number 1
25_FA_1: fullAdder
	port map (
		i0 => grid5(3)(25),
		i1 => grid5(4)(25),
		ci => grid5(5)(25),
		s => grid4(4)(25),
		co => grid4(1)(26) );

-- half adder c25, number 0
25_HA_0: halfAdder
	port map (
		i0 => grid5(6)(25),
		i1 => grid5(7)(25),
		s => grid4(5)(25),
		co => grid4(2)(26) );

-- move the other elements of the column
grid4(6)(25) <= grid5(8)(25);
grid4(7)(25) <= grid5(9)(25);
grid4(8)(25) <= grid5(10)(25);
grid4(9)(25) <= grid5(11)(25);

----------------------------- 
-- COLUMN 26
----------------------------- 
-- full adder c26, number 0
26_FA_0: fullAdder
	port map (
		i0 => grid5(0)(26),
		i1 => grid5(1)(26),
		ci => grid5(2)(26),
		s => grid4(3)(26),
		co => grid4(0)(27) );

-- full adder c26, number 1
26_FA_1: fullAdder
	port map (
		i0 => grid5(3)(26),
		i1 => grid5(4)(26),
		ci => grid5(5)(26),
		s => grid4(4)(26),
		co => grid4(1)(27) );

-- half adder c26, number 0
26_HA_0: halfAdder
	port map (
		i0 => grid5(6)(26),
		i1 => grid5(7)(26),
		s => grid4(5)(26),
		co => grid4(2)(27) );

-- move the other elements of the column
grid4(6)(26) <= grid5(8)(26);
grid4(7)(26) <= grid5(9)(26);
grid4(8)(26) <= grid5(10)(26);
grid4(9)(26) <= grid5(11)(26);

----------------------------- 
-- COLUMN 27
----------------------------- 
-- full adder c27, number 0
27_FA_0: fullAdder
	port map (
		i0 => grid5(0)(27),
		i1 => grid5(1)(27),
		ci => grid5(2)(27),
		s => grid4(3)(27),
		co => grid4(0)(28) );

-- full adder c27, number 1
27_FA_1: fullAdder
	port map (
		i0 => grid5(3)(27),
		i1 => grid5(4)(27),
		ci => grid5(5)(27),
		s => grid4(4)(27),
		co => grid4(1)(28) );

-- half adder c27, number 0
27_HA_0: halfAdder
	port map (
		i0 => grid5(6)(27),
		i1 => grid5(7)(27),
		s => grid4(5)(27),
		co => grid4(2)(28) );

-- move the other elements of the column
grid4(6)(27) <= grid5(8)(27);
grid4(7)(27) <= grid5(9)(27);
grid4(8)(27) <= grid5(10)(27);
grid4(9)(27) <= grid5(11)(27);

----------------------------- 
-- COLUMN 28
----------------------------- 
-- full adder c28, number 0
28_FA_0: fullAdder
	port map (
		i0 => grid5(0)(28),
		i1 => grid5(1)(28),
		ci => grid5(2)(28),
		s => grid4(3)(28),
		co => grid4(0)(29) );

-- full adder c28, number 1
28_FA_1: fullAdder
	port map (
		i0 => grid5(3)(28),
		i1 => grid5(4)(28),
		ci => grid5(5)(28),
		s => grid4(4)(28),
		co => grid4(1)(29) );

-- half adder c28, number 0
28_HA_0: halfAdder
	port map (
		i0 => grid5(6)(28),
		i1 => grid5(7)(28),
		s => grid4(5)(28),
		co => grid4(2)(29) );

-- move the other elements of the column
grid4(6)(28) <= grid5(8)(28);
grid4(7)(28) <= grid5(9)(28);
grid4(8)(28) <= grid5(10)(28);
grid4(9)(28) <= grid5(11)(28);

----------------------------- 
-- COLUMN 29
----------------------------- 
-- full adder c29, number 0
29_FA_0: fullAdder
	port map (
		i0 => grid5(0)(29),
		i1 => grid5(1)(29),
		ci => grid5(2)(29),
		s => grid4(3)(29),
		co => grid4(0)(30) );

-- full adder c29, number 1
29_FA_1: fullAdder
	port map (
		i0 => grid5(3)(29),
		i1 => grid5(4)(29),
		ci => grid5(5)(29),
		s => grid4(4)(29),
		co => grid4(1)(30) );

-- half adder c29, number 0
29_HA_0: halfAdder
	port map (
		i0 => grid5(6)(29),
		i1 => grid5(7)(29),
		s => grid4(5)(29),
		co => grid4(2)(30) );

-- move the other elements of the column
grid4(6)(29) <= grid5(8)(29);
grid4(7)(29) <= grid5(9)(29);
grid4(8)(29) <= grid5(10)(29);
grid4(9)(29) <= grid5(11)(29);

----------------------------- 
-- COLUMN 30
----------------------------- 
-- full adder c30, number 0
30_FA_0: fullAdder
	port map (
		i0 => grid5(0)(30),
		i1 => grid5(1)(30),
		ci => grid5(2)(30),
		s => grid4(3)(30),
		co => grid4(0)(31) );

-- full adder c30, number 1
30_FA_1: fullAdder
	port map (
		i0 => grid5(3)(30),
		i1 => grid5(4)(30),
		ci => grid5(5)(30),
		s => grid4(4)(30),
		co => grid4(1)(31) );

-- half adder c30, number 0
30_HA_0: halfAdder
	port map (
		i0 => grid5(6)(30),
		i1 => grid5(7)(30),
		s => grid4(5)(30),
		co => grid4(2)(31) );

-- move the other elements of the column
grid4(6)(30) <= grid5(8)(30);
grid4(7)(30) <= grid5(9)(30);
grid4(8)(30) <= grid5(10)(30);
grid4(9)(30) <= grid5(11)(30);

----------------------------- 
-- COLUMN 31
----------------------------- 
-- full adder c31, number 0
31_FA_0: fullAdder
	port map (
		i0 => grid5(0)(31),
		i1 => grid5(1)(31),
		ci => grid5(2)(31),
		s => grid4(3)(31),
		co => grid4(0)(32) );

-- full adder c31, number 1
31_FA_1: fullAdder
	port map (
		i0 => grid5(3)(31),
		i1 => grid5(4)(31),
		ci => grid5(5)(31),
		s => grid4(4)(31),
		co => grid4(1)(32) );

-- half adder c31, number 0
31_HA_0: halfAdder
	port map (
		i0 => grid5(6)(31),
		i1 => grid5(7)(31),
		s => grid4(5)(31),
		co => grid4(2)(32) );

-- move the other elements of the column
grid4(6)(31) <= grid5(8)(31);
grid4(7)(31) <= grid5(9)(31);
grid4(8)(31) <= grid5(10)(31);
grid4(9)(31) <= grid5(11)(31);

----------------------------- 
-- COLUMN 32
----------------------------- 
-- full adder c32, number 0
32_FA_0: fullAdder
	port map (
		i0 => grid5(0)(32),
		i1 => grid5(1)(32),
		ci => grid5(2)(32),
		s => grid4(3)(32),
		co => grid4(0)(33) );

-- full adder c32, number 1
32_FA_1: fullAdder
	port map (
		i0 => grid5(3)(32),
		i1 => grid5(4)(32),
		ci => grid5(5)(32),
		s => grid4(4)(32),
		co => grid4(1)(33) );

-- half adder c32, number 0
32_HA_0: halfAdder
	port map (
		i0 => grid5(6)(32),
		i1 => grid5(7)(32),
		s => grid4(5)(32),
		co => grid4(2)(33) );

-- move the other elements of the column
grid4(6)(32) <= grid5(8)(32);
grid4(7)(32) <= grid5(9)(32);
grid4(8)(32) <= grid5(10)(32);
grid4(9)(32) <= grid5(11)(32);

----------------------------- 
-- COLUMN 33
----------------------------- 
-- full adder c33, number 0
33_FA_0: fullAdder
	port map (
		i0 => grid5(0)(33),
		i1 => grid5(1)(33),
		ci => grid5(2)(33),
		s => grid4(3)(33),
		co => grid4(0)(34) );

-- full adder c33, number 1
33_FA_1: fullAdder
	port map (
		i0 => grid5(3)(33),
		i1 => grid5(4)(33),
		ci => grid5(5)(33),
		s => grid4(4)(33),
		co => grid4(1)(34) );

-- half adder c33, number 0
33_HA_0: halfAdder
	port map (
		i0 => grid5(6)(33),
		i1 => grid5(7)(33),
		s => grid4(5)(33),
		co => grid4(2)(34) );

-- move the other elements of the column
grid4(6)(33) <= grid5(8)(33);
grid4(7)(33) <= grid5(9)(33);
grid4(8)(33) <= grid5(10)(33);
grid4(9)(33) <= grid5(11)(33);

----------------------------- 
-- COLUMN 34
----------------------------- 
-- full adder c34, number 0
34_FA_0: fullAdder
	port map (
		i0 => grid5(0)(34),
		i1 => grid5(1)(34),
		ci => grid5(2)(34),
		s => grid4(3)(34),
		co => grid4(0)(35) );

-- full adder c34, number 1
34_FA_1: fullAdder
	port map (
		i0 => grid5(3)(34),
		i1 => grid5(4)(34),
		ci => grid5(5)(34),
		s => grid4(4)(34),
		co => grid4(1)(35) );

-- half adder c34, number 0
34_HA_0: halfAdder
	port map (
		i0 => grid5(6)(34),
		i1 => grid5(7)(34),
		s => grid4(5)(34),
		co => grid4(2)(35) );

-- move the other elements of the column
grid4(6)(34) <= grid5(8)(34);
grid4(7)(34) <= grid5(9)(34);
grid4(8)(34) <= grid5(10)(34);
grid4(9)(34) <= grid5(11)(34);

----------------------------- 
-- COLUMN 35
----------------------------- 
-- full adder c35, number 0
35_FA_0: fullAdder
	port map (
		i0 => grid5(0)(35),
		i1 => grid5(1)(35),
		ci => grid5(2)(35),
		s => grid4(3)(35),
		co => grid4(0)(36) );

-- full adder c35, number 1
35_FA_1: fullAdder
	port map (
		i0 => grid5(3)(35),
		i1 => grid5(4)(35),
		ci => grid5(5)(35),
		s => grid4(4)(35),
		co => grid4(1)(36) );

-- half adder c35, number 0
35_HA_0: halfAdder
	port map (
		i0 => grid5(6)(35),
		i1 => grid5(7)(35),
		s => grid4(5)(35),
		co => grid4(2)(36) );

-- move the other elements of the column
grid4(6)(35) <= grid5(8)(35);
grid4(7)(35) <= grid5(9)(35);
grid4(8)(35) <= grid5(10)(35);
grid4(9)(35) <= grid5(11)(35);

----------------------------- 
-- COLUMN 36
----------------------------- 
-- full adder c36, number 0
36_FA_0: fullAdder
	port map (
		i0 => grid5(0)(36),
		i1 => grid5(1)(36),
		ci => grid5(2)(36),
		s => grid4(3)(36),
		co => grid4(0)(37) );

-- full adder c36, number 1
36_FA_1: fullAdder
	port map (
		i0 => grid5(3)(36),
		i1 => grid5(4)(36),
		ci => grid5(5)(36),
		s => grid4(4)(36),
		co => grid4(1)(37) );

-- half adder c36, number 0
36_HA_0: halfAdder
	port map (
		i0 => grid5(6)(36),
		i1 => grid5(7)(36),
		s => grid4(5)(36),
		co => grid4(2)(37) );

-- move the other elements of the column
grid4(6)(36) <= grid5(8)(36);
grid4(7)(36) <= grid5(9)(36);
grid4(8)(36) <= grid5(10)(36);
grid4(9)(36) <= grid5(11)(36);

----------------------------- 
-- COLUMN 37
----------------------------- 
-- full adder c37, number 0
37_FA_0: fullAdder
	port map (
		i0 => grid5(0)(37),
		i1 => grid5(1)(37),
		ci => grid5(2)(37),
		s => grid4(3)(37),
		co => grid4(0)(38) );

-- full adder c37, number 1
37_FA_1: fullAdder
	port map (
		i0 => grid5(3)(37),
		i1 => grid5(4)(37),
		ci => grid5(5)(37),
		s => grid4(4)(37),
		co => grid4(1)(38) );

-- half adder c37, number 0
37_HA_0: halfAdder
	port map (
		i0 => grid5(6)(37),
		i1 => grid5(7)(37),
		s => grid4(5)(37),
		co => grid4(2)(38) );

-- move the other elements of the column
grid4(6)(37) <= grid5(8)(37);
grid4(7)(37) <= grid5(9)(37);
grid4(8)(37) <= grid5(10)(37);
grid4(9)(37) <= grid5(11)(37);

----------------------------- 
-- COLUMN 38
----------------------------- 
-- full adder c38, number 0
38_FA_0: fullAdder
	port map (
		i0 => grid5(0)(38),
		i1 => grid5(1)(38),
		ci => grid5(2)(38),
		s => grid4(3)(38),
		co => grid4(0)(39) );

-- full adder c38, number 1
38_FA_1: fullAdder
	port map (
		i0 => grid5(3)(38),
		i1 => grid5(4)(38),
		ci => grid5(5)(38),
		s => grid4(4)(38),
		co => grid4(1)(39) );

-- half adder c38, number 0
38_HA_0: halfAdder
	port map (
		i0 => grid5(6)(38),
		i1 => grid5(7)(38),
		s => grid4(5)(38),
		co => grid4(2)(39) );

-- move the other elements of the column
grid4(6)(38) <= grid5(8)(38);
grid4(7)(38) <= grid5(9)(38);
grid4(8)(38) <= grid5(10)(38);
grid4(9)(38) <= grid5(11)(38);

----------------------------- 
-- COLUMN 39
----------------------------- 
-- full adder c39, number 0
39_FA_0: fullAdder
	port map (
		i0 => grid5(0)(39),
		i1 => grid5(1)(39),
		ci => grid5(2)(39),
		s => grid4(3)(39),
		co => grid4(0)(40) );

-- full adder c39, number 1
39_FA_1: fullAdder
	port map (
		i0 => grid5(3)(39),
		i1 => grid5(4)(39),
		ci => grid5(5)(39),
		s => grid4(4)(39),
		co => grid4(1)(40) );

-- half adder c39, number 0
39_HA_0: halfAdder
	port map (
		i0 => grid5(6)(39),
		i1 => grid5(7)(39),
		s => grid4(5)(39),
		co => grid4(2)(40) );

-- move the other elements of the column
grid4(6)(39) <= grid5(8)(39);
grid4(7)(39) <= grid5(9)(39);
grid4(8)(39) <= grid5(10)(39);
grid4(9)(39) <= grid5(11)(39);

----------------------------- 
-- COLUMN 40
----------------------------- 
-- full adder c40, number 0
40_FA_0: fullAdder
	port map (
		i0 => grid5(0)(40),
		i1 => grid5(1)(40),
		ci => grid5(2)(40),
		s => grid4(3)(40),
		co => grid4(0)(41) );

-- full adder c40, number 1
40_FA_1: fullAdder
	port map (
		i0 => grid5(3)(40),
		i1 => grid5(4)(40),
		ci => grid5(5)(40),
		s => grid4(4)(40),
		co => grid4(1)(41) );

-- half adder c40, number 0
40_HA_0: halfAdder
	port map (
		i0 => grid5(6)(40),
		i1 => grid5(7)(40),
		s => grid4(5)(40),
		co => grid4(2)(41) );

-- move the other elements of the column
grid4(6)(40) <= grid5(8)(40);
grid4(7)(40) <= grid5(9)(40);
grid4(8)(40) <= grid5(10)(40);
grid4(9)(40) <= grid5(11)(40);

----------------------------- 
-- COLUMN 41
----------------------------- 
-- full adder c41, number 0
41_FA_0: fullAdder
	port map (
		i0 => grid5(0)(41),
		i1 => grid5(1)(41),
		ci => grid5(2)(41),
		s => grid4(3)(41),
		co => grid4(0)(42) );

-- full adder c41, number 1
41_FA_1: fullAdder
	port map (
		i0 => grid5(3)(41),
		i1 => grid5(4)(41),
		ci => grid5(5)(41),
		s => grid4(4)(41),
		co => grid4(1)(42) );

-- half adder c41, number 0
41_HA_0: halfAdder
	port map (
		i0 => grid5(6)(41),
		i1 => grid5(7)(41),
		s => grid4(5)(41),
		co => grid4(2)(42) );

-- move the other elements of the column
grid4(6)(41) <= grid5(8)(41);
grid4(7)(41) <= grid5(9)(41);
grid4(8)(41) <= grid5(10)(41);
grid4(9)(41) <= grid5(11)(41);

----------------------------- 
-- COLUMN 42
----------------------------- 
-- full adder c42, number 0
42_FA_0: fullAdder
	port map (
		i0 => grid5(0)(42),
		i1 => grid5(1)(42),
		ci => grid5(2)(42),
		s => grid4(3)(42),
		co => grid4(0)(43) );

-- full adder c42, number 1
42_FA_1: fullAdder
	port map (
		i0 => grid5(3)(42),
		i1 => grid5(4)(42),
		ci => grid5(5)(42),
		s => grid4(4)(42),
		co => grid4(1)(43) );

-- half adder c42, number 0
42_HA_0: halfAdder
	port map (
		i0 => grid5(6)(42),
		i1 => grid5(7)(42),
		s => grid4(5)(42),
		co => grid4(2)(43) );

-- move the other elements of the column
grid4(6)(42) <= grid5(8)(42);
grid4(7)(42) <= grid5(9)(42);
grid4(8)(42) <= grid5(10)(42);
grid4(9)(42) <= grid5(11)(42);

----------------------------- 
-- COLUMN 43
----------------------------- 
-- full adder c43, number 0
43_FA_0: fullAdder
	port map (
		i0 => grid5(0)(43),
		i1 => grid5(1)(43),
		ci => grid5(2)(43),
		s => grid4(3)(43),
		co => grid4(0)(44) );

-- full adder c43, number 1
43_FA_1: fullAdder
	port map (
		i0 => grid5(3)(43),
		i1 => grid5(4)(43),
		ci => grid5(5)(43),
		s => grid4(4)(43),
		co => grid4(1)(44) );

-- half adder c43, number 0
43_HA_0: halfAdder
	port map (
		i0 => grid5(6)(43),
		i1 => grid5(7)(43),
		s => grid4(5)(43),
		co => grid4(2)(44) );

-- move the other elements of the column
grid4(6)(43) <= grid5(8)(43);
grid4(7)(43) <= grid5(9)(43);
grid4(8)(43) <= grid5(10)(43);
grid4(9)(43) <= grid5(11)(43);

----------------------------- 
-- COLUMN 44
----------------------------- 
-- full adder c44, number 0
44_FA_0: fullAdder
	port map (
		i0 => grid5(0)(44),
		i1 => grid5(1)(44),
		ci => grid5(2)(44),
		s => grid4(3)(44),
		co => grid4(0)(45) );

-- full adder c44, number 1
44_FA_1: fullAdder
	port map (
		i0 => grid5(3)(44),
		i1 => grid5(4)(44),
		ci => grid5(5)(44),
		s => grid4(4)(44),
		co => grid4(1)(45) );

-- half adder c44, number 0
44_HA_0: halfAdder
	port map (
		i0 => grid5(6)(44),
		i1 => grid5(7)(44),
		s => grid4(5)(44),
		co => grid4(2)(45) );

-- move the other elements of the column
grid4(6)(44) <= grid5(8)(44);
grid4(7)(44) <= grid5(9)(44);
grid4(8)(44) <= grid5(10)(44);
grid4(9)(44) <= grid5(11)(44);

----------------------------- 
-- COLUMN 45
----------------------------- 
-- full adder c45, number 0
45_FA_0: fullAdder
	port map (
		i0 => grid5(0)(45),
		i1 => grid5(1)(45),
		ci => grid5(2)(45),
		s => grid4(3)(45),
		co => grid4(0)(46) );

-- full adder c45, number 1
45_FA_1: fullAdder
	port map (
		i0 => grid5(3)(45),
		i1 => grid5(4)(45),
		ci => grid5(5)(45),
		s => grid4(4)(45),
		co => grid4(1)(46) );

-- half adder c45, number 0
45_HA_0: halfAdder
	port map (
		i0 => grid5(6)(45),
		i1 => grid5(7)(45),
		s => grid4(5)(45),
		co => grid4(2)(46) );

-- move the other elements of the column
grid4(6)(45) <= grid5(8)(45);
grid4(7)(45) <= grid5(9)(45);
grid4(8)(45) <= grid5(10)(45);
grid4(9)(45) <= grid5(11)(45);

