
module iir_filter_DW01_add_9 ( A, B, CI, SUM, CO );
  input [45:0] A;
  input [45:0] B;
  output [45:0] SUM;
  input CI;
  output CO;
  wire   A_21_, A_20_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112;
  assign SUM[21] = A_21_;
  assign A_21_ = A[21];
  assign SUM[20] = A_20_;
  assign A_20_ = A[20];

  XOR2_X1 U2 ( .A(n1), .B(n2), .Z(SUM[45]) );
  XOR2_X1 U3 ( .A(B[45]), .B(A[45]), .Z(n2) );
  OAI21_X1 U4 ( .B1(n3), .B2(n4), .A(n5), .ZN(n1) );
  OAI21_X1 U5 ( .B1(A[44]), .B2(n6), .A(B[44]), .ZN(n5) );
  INV_X1 U6 ( .A(n3), .ZN(n6) );
  INV_X1 U7 ( .A(A[44]), .ZN(n4) );
  AOI21_X1 U8 ( .B1(A[43]), .B2(B[43]), .A(n7), .ZN(n3) );
  INV_X1 U9 ( .A(n8), .ZN(n7) );
  OAI22_X1 U10 ( .A1(n9), .A2(n10), .B1(A[43]), .B2(B[43]), .ZN(n8) );
  AOI21_X1 U11 ( .B1(n11), .B2(n12), .A(n13), .ZN(n9) );
  NAND3_X1 U12 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n12) );
  AOI21_X1 U13 ( .B1(n17), .B2(n16), .A(n18), .ZN(n11) );
  INV_X1 U14 ( .A(n19), .ZN(n18) );
  XOR2_X1 U15 ( .A(n20), .B(n21), .Z(SUM[42]) );
  NOR2_X1 U16 ( .A1(n10), .A2(n13), .ZN(n21) );
  NOR2_X1 U17 ( .A1(B[42]), .A2(A[42]), .ZN(n13) );
  AND2_X1 U18 ( .A1(B[42]), .A2(A[42]), .ZN(n10) );
  OAI21_X1 U19 ( .B1(n22), .B2(n23), .A(n19), .ZN(n20) );
  XOR2_X1 U20 ( .A(n24), .B(n23), .Z(SUM[41]) );
  AOI21_X1 U21 ( .B1(n15), .B2(n14), .A(n17), .ZN(n23) );
  INV_X1 U22 ( .A(n25), .ZN(n15) );
  NAND2_X1 U23 ( .A1(n16), .A2(n19), .ZN(n24) );
  NAND2_X1 U24 ( .A1(B[41]), .A2(A[41]), .ZN(n19) );
  INV_X1 U25 ( .A(n22), .ZN(n16) );
  NOR2_X1 U26 ( .A1(B[41]), .A2(A[41]), .ZN(n22) );
  XOR2_X1 U27 ( .A(n14), .B(n26), .Z(SUM[40]) );
  NOR2_X1 U28 ( .A1(n17), .A2(n25), .ZN(n26) );
  NOR2_X1 U29 ( .A1(B[40]), .A2(A[40]), .ZN(n25) );
  AND2_X1 U30 ( .A1(B[40]), .A2(A[40]), .ZN(n17) );
  OAI21_X1 U31 ( .B1(n27), .B2(n28), .A(n29), .ZN(n14) );
  XOR2_X1 U32 ( .A(n30), .B(n28), .Z(SUM[39]) );
  AOI21_X1 U33 ( .B1(n31), .B2(n32), .A(n33), .ZN(n28) );
  INV_X1 U34 ( .A(n34), .ZN(n31) );
  NAND2_X1 U35 ( .A1(n35), .A2(n29), .ZN(n30) );
  NAND2_X1 U36 ( .A1(B[39]), .A2(A[39]), .ZN(n29) );
  INV_X1 U37 ( .A(n27), .ZN(n35) );
  NOR2_X1 U38 ( .A1(B[39]), .A2(A[39]), .ZN(n27) );
  XOR2_X1 U39 ( .A(n32), .B(n36), .Z(SUM[38]) );
  NOR2_X1 U40 ( .A1(n33), .A2(n34), .ZN(n36) );
  NOR2_X1 U41 ( .A1(B[38]), .A2(A[38]), .ZN(n34) );
  AND2_X1 U42 ( .A1(B[38]), .A2(A[38]), .ZN(n33) );
  OAI21_X1 U43 ( .B1(n37), .B2(n38), .A(n39), .ZN(n32) );
  XOR2_X1 U44 ( .A(n40), .B(n38), .Z(SUM[37]) );
  AOI21_X1 U45 ( .B1(n41), .B2(n42), .A(n43), .ZN(n38) );
  INV_X1 U46 ( .A(n44), .ZN(n41) );
  NAND2_X1 U47 ( .A1(n45), .A2(n39), .ZN(n40) );
  NAND2_X1 U48 ( .A1(B[37]), .A2(A[37]), .ZN(n39) );
  INV_X1 U49 ( .A(n37), .ZN(n45) );
  NOR2_X1 U50 ( .A1(B[37]), .A2(A[37]), .ZN(n37) );
  XOR2_X1 U51 ( .A(n42), .B(n46), .Z(SUM[36]) );
  NOR2_X1 U52 ( .A1(n43), .A2(n44), .ZN(n46) );
  NOR2_X1 U53 ( .A1(B[36]), .A2(A[36]), .ZN(n44) );
  AND2_X1 U54 ( .A1(B[36]), .A2(A[36]), .ZN(n43) );
  OAI21_X1 U55 ( .B1(n47), .B2(n48), .A(n49), .ZN(n42) );
  XOR2_X1 U56 ( .A(n50), .B(n48), .Z(SUM[35]) );
  AOI21_X1 U57 ( .B1(n51), .B2(n52), .A(n53), .ZN(n48) );
  INV_X1 U58 ( .A(n54), .ZN(n51) );
  NAND2_X1 U59 ( .A1(n55), .A2(n49), .ZN(n50) );
  NAND2_X1 U60 ( .A1(B[35]), .A2(A[35]), .ZN(n49) );
  INV_X1 U61 ( .A(n47), .ZN(n55) );
  NOR2_X1 U62 ( .A1(B[35]), .A2(A[35]), .ZN(n47) );
  XOR2_X1 U63 ( .A(n52), .B(n56), .Z(SUM[34]) );
  NOR2_X1 U64 ( .A1(n53), .A2(n54), .ZN(n56) );
  NOR2_X1 U65 ( .A1(B[34]), .A2(A[34]), .ZN(n54) );
  AND2_X1 U66 ( .A1(B[34]), .A2(A[34]), .ZN(n53) );
  OAI21_X1 U67 ( .B1(n57), .B2(n58), .A(n59), .ZN(n52) );
  XOR2_X1 U68 ( .A(n60), .B(n58), .Z(SUM[33]) );
  AOI21_X1 U69 ( .B1(n61), .B2(n62), .A(n63), .ZN(n58) );
  INV_X1 U70 ( .A(n64), .ZN(n61) );
  NAND2_X1 U71 ( .A1(n65), .A2(n59), .ZN(n60) );
  NAND2_X1 U72 ( .A1(B[33]), .A2(A[33]), .ZN(n59) );
  INV_X1 U73 ( .A(n57), .ZN(n65) );
  NOR2_X1 U74 ( .A1(B[33]), .A2(A[33]), .ZN(n57) );
  XOR2_X1 U75 ( .A(n62), .B(n66), .Z(SUM[32]) );
  NOR2_X1 U76 ( .A1(n63), .A2(n64), .ZN(n66) );
  NOR2_X1 U77 ( .A1(B[32]), .A2(A[32]), .ZN(n64) );
  AND2_X1 U78 ( .A1(B[32]), .A2(A[32]), .ZN(n63) );
  OAI21_X1 U79 ( .B1(n67), .B2(n68), .A(n69), .ZN(n62) );
  XOR2_X1 U80 ( .A(n70), .B(n68), .Z(SUM[31]) );
  AOI21_X1 U81 ( .B1(n71), .B2(n72), .A(n73), .ZN(n68) );
  INV_X1 U82 ( .A(n74), .ZN(n71) );
  NAND2_X1 U83 ( .A1(n75), .A2(n69), .ZN(n70) );
  NAND2_X1 U84 ( .A1(B[31]), .A2(A[31]), .ZN(n69) );
  INV_X1 U85 ( .A(n67), .ZN(n75) );
  NOR2_X1 U86 ( .A1(B[31]), .A2(A[31]), .ZN(n67) );
  XOR2_X1 U87 ( .A(n72), .B(n76), .Z(SUM[30]) );
  NOR2_X1 U88 ( .A1(n73), .A2(n74), .ZN(n76) );
  NOR2_X1 U89 ( .A1(B[30]), .A2(A[30]), .ZN(n74) );
  AND2_X1 U90 ( .A1(B[30]), .A2(A[30]), .ZN(n73) );
  OAI21_X1 U91 ( .B1(n77), .B2(n78), .A(n79), .ZN(n72) );
  XOR2_X1 U92 ( .A(n80), .B(n78), .Z(SUM[29]) );
  AOI21_X1 U93 ( .B1(n81), .B2(n82), .A(n83), .ZN(n78) );
  INV_X1 U94 ( .A(n84), .ZN(n81) );
  NAND2_X1 U95 ( .A1(n85), .A2(n79), .ZN(n80) );
  NAND2_X1 U96 ( .A1(B[29]), .A2(A[29]), .ZN(n79) );
  INV_X1 U97 ( .A(n77), .ZN(n85) );
  NOR2_X1 U98 ( .A1(B[29]), .A2(A[29]), .ZN(n77) );
  XOR2_X1 U99 ( .A(n82), .B(n86), .Z(SUM[28]) );
  NOR2_X1 U100 ( .A1(n83), .A2(n84), .ZN(n86) );
  NOR2_X1 U101 ( .A1(B[28]), .A2(A[28]), .ZN(n84) );
  AND2_X1 U102 ( .A1(B[28]), .A2(A[28]), .ZN(n83) );
  OAI21_X1 U103 ( .B1(n87), .B2(n88), .A(n89), .ZN(n82) );
  XOR2_X1 U104 ( .A(n90), .B(n88), .Z(SUM[27]) );
  AOI21_X1 U105 ( .B1(n91), .B2(n92), .A(n93), .ZN(n88) );
  INV_X1 U106 ( .A(n94), .ZN(n92) );
  NAND2_X1 U107 ( .A1(n95), .A2(n89), .ZN(n90) );
  NAND2_X1 U108 ( .A1(B[27]), .A2(A[27]), .ZN(n89) );
  INV_X1 U109 ( .A(n87), .ZN(n95) );
  NOR2_X1 U110 ( .A1(B[27]), .A2(A[27]), .ZN(n87) );
  XOR2_X1 U111 ( .A(n91), .B(n96), .Z(SUM[26]) );
  NOR2_X1 U112 ( .A1(n93), .A2(n94), .ZN(n96) );
  NOR2_X1 U113 ( .A1(B[26]), .A2(A[26]), .ZN(n94) );
  AND2_X1 U114 ( .A1(B[26]), .A2(A[26]), .ZN(n93) );
  OAI21_X1 U115 ( .B1(n97), .B2(n98), .A(n99), .ZN(n91) );
  XOR2_X1 U116 ( .A(n100), .B(n98), .Z(SUM[25]) );
  AOI21_X1 U117 ( .B1(n101), .B2(n102), .A(n103), .ZN(n98) );
  INV_X1 U118 ( .A(n104), .ZN(n101) );
  NAND2_X1 U119 ( .A1(n105), .A2(n99), .ZN(n100) );
  NAND2_X1 U120 ( .A1(B[25]), .A2(A[25]), .ZN(n99) );
  INV_X1 U121 ( .A(n97), .ZN(n105) );
  NOR2_X1 U122 ( .A1(B[25]), .A2(A[25]), .ZN(n97) );
  XOR2_X1 U123 ( .A(n102), .B(n106), .Z(SUM[24]) );
  NOR2_X1 U124 ( .A1(n103), .A2(n104), .ZN(n106) );
  NOR2_X1 U125 ( .A1(B[24]), .A2(A[24]), .ZN(n104) );
  AND2_X1 U126 ( .A1(B[24]), .A2(A[24]), .ZN(n103) );
  OAI21_X1 U127 ( .B1(n107), .B2(n108), .A(n109), .ZN(n102) );
  XOR2_X1 U128 ( .A(n108), .B(n110), .Z(SUM[23]) );
  NAND2_X1 U129 ( .A1(n111), .A2(n109), .ZN(n110) );
  NAND2_X1 U130 ( .A1(B[23]), .A2(A[23]), .ZN(n109) );
  INV_X1 U131 ( .A(n107), .ZN(n111) );
  NOR2_X1 U132 ( .A1(B[23]), .A2(A[23]), .ZN(n107) );
  INV_X1 U133 ( .A(n112), .ZN(SUM[22]) );
  OAI21_X1 U134 ( .B1(B[22]), .B2(A[22]), .A(n108), .ZN(n112) );
  NAND2_X1 U135 ( .A1(B[22]), .A2(A[22]), .ZN(n108) );
endmodule


module iir_filter_DW02_mult_5 ( A, B, TC, PRODUCT );
  input [23:0] A;
  input [23:0] B;
  output [47:0] PRODUCT;
  input TC;
  wire   ab_23__23_, ab_23__22_, ab_23__21_, ab_23__20_, ab_23__19_,
         ab_23__18_, ab_23__17_, ab_23__16_, ab_23__15_, ab_23__14_,
         ab_23__13_, ab_23__12_, ab_23__11_, ab_23__10_, ab_23__9_, ab_23__8_,
         ab_23__7_, ab_23__6_, ab_23__5_, ab_23__4_, ab_23__3_, ab_23__2_,
         ab_23__1_, ab_23__0_, ab_22__23_, ab_22__22_, ab_22__21_, ab_22__20_,
         ab_22__19_, ab_22__18_, ab_22__17_, ab_22__16_, ab_22__15_,
         ab_22__14_, ab_22__13_, ab_22__12_, ab_22__11_, ab_22__10_, ab_22__9_,
         ab_22__8_, ab_22__7_, ab_22__6_, ab_22__5_, ab_22__4_, ab_22__3_,
         ab_22__2_, ab_22__1_, ab_22__0_, ab_21__23_, ab_21__22_, ab_21__21_,
         ab_21__20_, ab_21__19_, ab_21__18_, ab_21__17_, ab_21__16_,
         ab_21__15_, ab_21__14_, ab_21__13_, ab_21__12_, ab_21__11_,
         ab_21__10_, ab_21__9_, ab_21__8_, ab_21__7_, ab_21__6_, ab_21__5_,
         ab_21__4_, ab_21__3_, ab_21__2_, ab_21__1_, ab_21__0_, ab_20__23_,
         ab_20__22_, ab_20__21_, ab_20__20_, ab_20__19_, ab_20__18_,
         ab_20__17_, ab_20__16_, ab_20__15_, ab_20__14_, ab_20__13_,
         ab_20__12_, ab_20__11_, ab_20__10_, ab_20__9_, ab_20__8_, ab_20__7_,
         ab_20__6_, ab_20__5_, ab_20__4_, ab_20__3_, ab_20__2_, ab_20__1_,
         ab_20__0_, ab_19__23_, ab_19__22_, ab_19__21_, ab_19__20_, ab_19__19_,
         ab_19__18_, ab_19__17_, ab_19__16_, ab_19__15_, ab_19__14_,
         ab_19__13_, ab_19__12_, ab_19__11_, ab_19__10_, ab_19__9_, ab_19__8_,
         ab_19__7_, ab_19__6_, ab_19__5_, ab_19__4_, ab_19__3_, ab_19__2_,
         ab_19__1_, ab_19__0_, ab_18__23_, ab_18__22_, ab_18__21_, ab_18__20_,
         ab_18__19_, ab_18__18_, ab_18__17_, ab_18__16_, ab_18__15_,
         ab_18__14_, ab_18__13_, ab_18__12_, ab_18__11_, ab_18__10_, ab_18__9_,
         ab_18__8_, ab_18__7_, ab_18__6_, ab_18__5_, ab_18__4_, ab_18__3_,
         ab_18__2_, ab_18__1_, ab_18__0_, ab_17__23_, ab_17__22_, ab_17__21_,
         ab_17__20_, ab_17__19_, ab_17__18_, ab_17__17_, ab_17__16_,
         ab_17__15_, ab_17__14_, ab_17__13_, ab_17__12_, ab_17__11_,
         ab_17__10_, ab_17__9_, ab_17__8_, ab_17__7_, ab_17__6_, ab_17__5_,
         ab_17__4_, ab_17__3_, ab_17__2_, ab_17__1_, ab_17__0_, ab_16__23_,
         ab_16__22_, ab_16__21_, ab_16__20_, ab_16__19_, ab_16__18_,
         ab_16__17_, ab_16__16_, ab_16__15_, ab_16__14_, ab_16__13_,
         ab_16__12_, ab_16__11_, ab_16__10_, ab_16__9_, ab_16__8_, ab_16__7_,
         ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_, ab_16__1_,
         ab_16__0_, ab_15__23_, ab_15__22_, ab_15__21_, ab_15__20_, ab_15__19_,
         ab_15__18_, ab_15__17_, ab_15__16_, ab_15__15_, ab_15__14_,
         ab_15__13_, ab_15__12_, ab_15__11_, ab_15__10_, ab_15__9_, ab_15__8_,
         ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_, ab_15__3_, ab_15__2_,
         ab_15__1_, ab_15__0_, ab_14__23_, ab_14__22_, ab_14__21_, ab_14__20_,
         ab_14__19_, ab_14__18_, ab_14__17_, ab_14__16_, ab_14__15_,
         ab_14__14_, ab_14__13_, ab_14__12_, ab_14__11_, ab_14__10_, ab_14__9_,
         ab_14__8_, ab_14__7_, ab_14__6_, ab_14__5_, ab_14__4_, ab_14__3_,
         ab_14__2_, ab_14__1_, ab_14__0_, ab_13__23_, ab_13__22_, ab_13__21_,
         ab_13__20_, ab_13__19_, ab_13__18_, ab_13__17_, ab_13__16_,
         ab_13__15_, ab_13__14_, ab_13__13_, ab_13__12_, ab_13__11_,
         ab_13__10_, ab_13__9_, ab_13__8_, ab_13__7_, ab_13__6_, ab_13__5_,
         ab_13__4_, ab_13__3_, ab_13__2_, ab_13__1_, ab_13__0_, ab_12__23_,
         ab_12__22_, ab_12__21_, ab_12__20_, ab_12__19_, ab_12__18_,
         ab_12__17_, ab_12__16_, ab_12__15_, ab_12__14_, ab_12__13_,
         ab_12__12_, ab_12__11_, ab_12__10_, ab_12__9_, ab_12__8_, ab_12__7_,
         ab_12__6_, ab_12__5_, ab_12__4_, ab_12__3_, ab_12__2_, ab_12__1_,
         ab_12__0_, ab_11__23_, ab_11__22_, ab_11__21_, ab_11__20_, ab_11__19_,
         ab_11__18_, ab_11__17_, ab_11__16_, ab_11__15_, ab_11__14_,
         ab_11__13_, ab_11__12_, ab_11__11_, ab_11__10_, ab_11__9_, ab_11__8_,
         ab_11__7_, ab_11__6_, ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_,
         ab_11__1_, ab_11__0_, ab_10__23_, ab_10__22_, ab_10__21_, ab_10__20_,
         ab_10__19_, ab_10__18_, ab_10__17_, ab_10__16_, ab_10__15_,
         ab_10__14_, ab_10__13_, ab_10__12_, ab_10__11_, ab_10__10_, ab_10__9_,
         ab_10__8_, ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_,
         ab_10__2_, ab_10__1_, ab_10__0_, ab_9__23_, ab_9__22_, ab_9__21_,
         ab_9__20_, ab_9__19_, ab_9__18_, ab_9__17_, ab_9__16_, ab_9__15_,
         ab_9__14_, ab_9__13_, ab_9__12_, ab_9__11_, ab_9__10_, ab_9__9_,
         ab_9__8_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_,
         ab_9__1_, ab_9__0_, ab_8__23_, ab_8__22_, ab_8__21_, ab_8__20_,
         ab_8__19_, ab_8__18_, ab_8__17_, ab_8__16_, ab_8__15_, ab_8__14_,
         ab_8__13_, ab_8__12_, ab_8__11_, ab_8__10_, ab_8__9_, ab_8__8_,
         ab_8__7_, ab_8__6_, ab_8__5_, ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_,
         ab_8__0_, ab_7__23_, ab_7__22_, ab_7__21_, ab_7__20_, ab_7__19_,
         ab_7__18_, ab_7__17_, ab_7__16_, ab_7__15_, ab_7__14_, ab_7__13_,
         ab_7__12_, ab_7__11_, ab_7__10_, ab_7__9_, ab_7__8_, ab_7__7_,
         ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_,
         ab_6__23_, ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_, ab_6__18_,
         ab_6__17_, ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_, ab_6__12_,
         ab_6__11_, ab_6__10_, ab_6__9_, ab_6__8_, ab_6__7_, ab_6__6_,
         ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_, ab_5__23_,
         ab_5__22_, ab_5__21_, ab_5__20_, ab_5__19_, ab_5__18_, ab_5__17_,
         ab_5__16_, ab_5__15_, ab_5__14_, ab_5__13_, ab_5__12_, ab_5__11_,
         ab_5__10_, ab_5__9_, ab_5__8_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_,
         ab_5__3_, ab_5__2_, ab_5__1_, ab_5__0_, ab_4__23_, ab_4__22_,
         ab_4__21_, ab_4__20_, ab_4__19_, ab_4__18_, ab_4__17_, ab_4__16_,
         ab_4__15_, ab_4__14_, ab_4__13_, ab_4__12_, ab_4__11_, ab_4__10_,
         ab_4__9_, ab_4__8_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_,
         ab_4__2_, ab_4__1_, ab_4__0_, ab_3__23_, ab_3__22_, ab_3__21_,
         ab_3__20_, ab_3__19_, ab_3__18_, ab_3__17_, ab_3__16_, ab_3__15_,
         ab_3__14_, ab_3__13_, ab_3__12_, ab_3__11_, ab_3__10_, ab_3__9_,
         ab_3__8_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_, ab_3__2_,
         ab_3__1_, ab_3__0_, ab_2__23_, ab_2__22_, ab_2__21_, ab_2__20_,
         ab_2__19_, ab_2__18_, ab_2__17_, ab_2__16_, ab_2__15_, ab_2__14_,
         ab_2__13_, ab_2__12_, ab_2__11_, ab_2__10_, ab_2__9_, ab_2__8_,
         ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_,
         ab_2__0_, ab_1__23_, ab_1__22_, ab_1__21_, ab_1__20_, ab_1__19_,
         ab_1__18_, ab_1__17_, ab_1__16_, ab_1__15_, ab_1__14_, ab_1__13_,
         ab_1__12_, ab_1__11_, ab_1__10_, ab_1__9_, ab_1__8_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_0__23_,
         ab_0__22_, ab_0__21_, ab_0__20_, ab_0__19_, ab_0__18_, ab_0__17_,
         ab_0__16_, ab_0__15_, ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_,
         ab_0__10_, ab_0__9_, ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_23__23_, CARRYB_23__22_, CARRYB_23__21_,
         CARRYB_23__20_, CARRYB_23__19_, CARRYB_23__18_, CARRYB_23__17_,
         CARRYB_23__16_, CARRYB_23__15_, CARRYB_23__14_, CARRYB_23__13_,
         CARRYB_23__12_, CARRYB_23__11_, CARRYB_23__10_, CARRYB_23__9_,
         CARRYB_23__8_, CARRYB_23__7_, CARRYB_23__6_, CARRYB_23__5_,
         CARRYB_23__4_, CARRYB_23__3_, CARRYB_23__2_, CARRYB_23__1_,
         CARRYB_23__0_, CARRYB_22__22_, CARRYB_22__21_, CARRYB_22__20_,
         CARRYB_22__19_, CARRYB_22__18_, CARRYB_22__17_, CARRYB_22__16_,
         CARRYB_22__15_, CARRYB_22__14_, CARRYB_22__13_, CARRYB_22__12_,
         CARRYB_22__11_, CARRYB_22__10_, CARRYB_22__9_, CARRYB_22__8_,
         CARRYB_22__7_, CARRYB_22__6_, CARRYB_22__5_, CARRYB_22__4_,
         CARRYB_22__3_, CARRYB_22__2_, CARRYB_22__1_, CARRYB_22__0_,
         CARRYB_21__22_, CARRYB_21__21_, CARRYB_21__20_, CARRYB_21__19_,
         CARRYB_21__18_, CARRYB_21__17_, CARRYB_21__16_, CARRYB_21__15_,
         CARRYB_21__14_, CARRYB_21__13_, CARRYB_21__12_, CARRYB_21__11_,
         CARRYB_21__10_, CARRYB_21__9_, CARRYB_21__8_, CARRYB_21__7_,
         CARRYB_21__6_, CARRYB_21__5_, CARRYB_21__4_, CARRYB_21__3_,
         CARRYB_21__2_, CARRYB_21__1_, CARRYB_21__0_, CARRYB_20__22_,
         CARRYB_20__21_, CARRYB_20__20_, CARRYB_20__19_, CARRYB_20__18_,
         CARRYB_20__17_, CARRYB_20__16_, CARRYB_20__15_, CARRYB_20__14_,
         CARRYB_20__13_, CARRYB_20__12_, CARRYB_20__11_, CARRYB_20__10_,
         CARRYB_20__9_, CARRYB_20__8_, CARRYB_20__7_, CARRYB_20__6_,
         CARRYB_20__5_, CARRYB_20__4_, CARRYB_20__3_, CARRYB_20__2_,
         CARRYB_20__1_, CARRYB_20__0_, CARRYB_19__22_, CARRYB_19__21_,
         CARRYB_19__20_, CARRYB_19__19_, CARRYB_19__18_, CARRYB_19__17_,
         CARRYB_19__16_, CARRYB_19__15_, CARRYB_19__14_, CARRYB_19__13_,
         CARRYB_19__12_, CARRYB_19__11_, CARRYB_19__10_, CARRYB_19__9_,
         CARRYB_19__8_, CARRYB_19__7_, CARRYB_19__6_, CARRYB_19__5_,
         CARRYB_19__4_, CARRYB_19__3_, CARRYB_19__2_, CARRYB_19__1_,
         CARRYB_19__0_, CARRYB_18__22_, CARRYB_18__21_, CARRYB_18__20_,
         CARRYB_18__19_, CARRYB_18__18_, CARRYB_18__17_, CARRYB_18__16_,
         CARRYB_18__15_, CARRYB_18__14_, CARRYB_18__13_, CARRYB_18__12_,
         CARRYB_18__11_, CARRYB_18__10_, CARRYB_18__9_, CARRYB_18__8_,
         CARRYB_18__7_, CARRYB_18__6_, CARRYB_18__5_, CARRYB_18__4_,
         CARRYB_18__3_, CARRYB_18__2_, CARRYB_18__1_, CARRYB_18__0_,
         CARRYB_17__22_, CARRYB_17__21_, CARRYB_17__20_, CARRYB_17__19_,
         CARRYB_17__18_, CARRYB_17__17_, CARRYB_17__16_, CARRYB_17__15_,
         CARRYB_17__14_, CARRYB_17__13_, CARRYB_17__12_, CARRYB_17__11_,
         CARRYB_17__10_, CARRYB_17__9_, CARRYB_17__8_, CARRYB_17__7_,
         CARRYB_17__6_, CARRYB_17__5_, CARRYB_17__4_, CARRYB_17__3_,
         CARRYB_17__2_, CARRYB_17__1_, CARRYB_17__0_, CARRYB_16__22_,
         CARRYB_16__21_, CARRYB_16__20_, CARRYB_16__19_, CARRYB_16__18_,
         CARRYB_16__17_, CARRYB_16__16_, CARRYB_16__15_, CARRYB_16__14_,
         CARRYB_16__13_, CARRYB_16__12_, CARRYB_16__11_, CARRYB_16__10_,
         CARRYB_16__9_, CARRYB_16__8_, CARRYB_16__7_, CARRYB_16__6_,
         CARRYB_16__5_, CARRYB_16__4_, CARRYB_16__3_, CARRYB_16__2_,
         CARRYB_16__1_, CARRYB_16__0_, CARRYB_15__22_, CARRYB_15__21_,
         CARRYB_15__20_, CARRYB_15__19_, CARRYB_15__18_, CARRYB_15__17_,
         CARRYB_15__16_, CARRYB_15__15_, CARRYB_15__14_, CARRYB_15__13_,
         CARRYB_15__12_, CARRYB_15__11_, CARRYB_15__10_, CARRYB_15__9_,
         CARRYB_15__8_, CARRYB_15__7_, CARRYB_15__6_, CARRYB_15__5_,
         CARRYB_15__4_, CARRYB_15__3_, CARRYB_15__2_, CARRYB_15__1_,
         CARRYB_15__0_, CARRYB_14__22_, CARRYB_14__21_, CARRYB_14__20_,
         CARRYB_14__19_, CARRYB_14__18_, CARRYB_14__17_, CARRYB_14__16_,
         CARRYB_14__15_, CARRYB_14__14_, CARRYB_14__13_, CARRYB_14__12_,
         CARRYB_14__11_, CARRYB_14__10_, CARRYB_14__9_, CARRYB_14__8_,
         CARRYB_14__7_, CARRYB_14__6_, CARRYB_14__5_, CARRYB_14__4_,
         CARRYB_14__3_, CARRYB_14__2_, CARRYB_14__1_, CARRYB_14__0_,
         CARRYB_13__22_, CARRYB_13__21_, CARRYB_13__20_, CARRYB_13__19_,
         CARRYB_13__18_, CARRYB_13__17_, CARRYB_13__16_, CARRYB_13__15_,
         CARRYB_13__14_, CARRYB_13__13_, CARRYB_13__12_, CARRYB_13__11_,
         CARRYB_13__10_, CARRYB_13__9_, CARRYB_13__8_, CARRYB_13__7_,
         CARRYB_13__6_, CARRYB_13__5_, CARRYB_13__4_, CARRYB_13__3_,
         CARRYB_13__2_, CARRYB_13__1_, CARRYB_13__0_, CARRYB_12__22_,
         CARRYB_12__21_, CARRYB_12__20_, CARRYB_12__19_, CARRYB_12__18_,
         CARRYB_12__17_, CARRYB_12__16_, CARRYB_12__15_, CARRYB_12__14_,
         CARRYB_12__13_, CARRYB_12__12_, CARRYB_12__11_, CARRYB_12__10_,
         CARRYB_12__9_, CARRYB_12__8_, CARRYB_12__7_, CARRYB_12__6_,
         CARRYB_12__5_, CARRYB_12__4_, CARRYB_12__3_, CARRYB_12__2_,
         CARRYB_12__1_, CARRYB_12__0_, CARRYB_11__22_, CARRYB_11__21_,
         CARRYB_11__20_, CARRYB_11__19_, CARRYB_11__18_, CARRYB_11__17_,
         CARRYB_11__16_, CARRYB_11__15_, CARRYB_11__14_, CARRYB_11__13_,
         CARRYB_11__12_, CARRYB_11__11_, CARRYB_11__10_, CARRYB_11__9_,
         CARRYB_11__8_, CARRYB_11__7_, CARRYB_11__6_, CARRYB_11__5_,
         CARRYB_11__4_, CARRYB_11__3_, CARRYB_11__2_, CARRYB_11__1_,
         CARRYB_11__0_, CARRYB_10__22_, CARRYB_10__21_, CARRYB_10__20_,
         CARRYB_10__19_, CARRYB_10__18_, CARRYB_10__17_, CARRYB_10__16_,
         CARRYB_10__15_, CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_,
         CARRYB_10__11_, CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_,
         CARRYB_10__7_, CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_,
         CARRYB_10__3_, CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_,
         CARRYB_9__22_, CARRYB_9__21_, CARRYB_9__20_, CARRYB_9__19_,
         CARRYB_9__18_, CARRYB_9__17_, CARRYB_9__16_, CARRYB_9__15_,
         CARRYB_9__14_, CARRYB_9__13_, CARRYB_9__12_, CARRYB_9__11_,
         CARRYB_9__10_, CARRYB_9__9_, CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_,
         CARRYB_9__5_, CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_,
         CARRYB_9__0_, CARRYB_8__22_, CARRYB_8__21_, CARRYB_8__20_,
         CARRYB_8__19_, CARRYB_8__18_, CARRYB_8__17_, CARRYB_8__16_,
         CARRYB_8__15_, CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_,
         CARRYB_8__11_, CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_,
         CARRYB_8__7_, CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_,
         CARRYB_8__2_, CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__22_,
         CARRYB_7__21_, CARRYB_7__20_, CARRYB_7__19_, CARRYB_7__18_,
         CARRYB_7__17_, CARRYB_7__16_, CARRYB_7__15_, CARRYB_7__14_,
         CARRYB_7__13_, CARRYB_7__12_, CARRYB_7__11_, CARRYB_7__10_,
         CARRYB_7__9_, CARRYB_7__8_, CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_,
         CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_,
         CARRYB_6__22_, CARRYB_6__21_, CARRYB_6__20_, CARRYB_6__19_,
         CARRYB_6__18_, CARRYB_6__17_, CARRYB_6__16_, CARRYB_6__15_,
         CARRYB_6__14_, CARRYB_6__13_, CARRYB_6__12_, CARRYB_6__11_,
         CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_, CARRYB_6__7_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__22_, CARRYB_5__21_, CARRYB_5__20_,
         CARRYB_5__19_, CARRYB_5__18_, CARRYB_5__17_, CARRYB_5__16_,
         CARRYB_5__15_, CARRYB_5__14_, CARRYB_5__13_, CARRYB_5__12_,
         CARRYB_5__11_, CARRYB_5__10_, CARRYB_5__9_, CARRYB_5__8_,
         CARRYB_5__7_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__22_,
         CARRYB_4__21_, CARRYB_4__20_, CARRYB_4__19_, CARRYB_4__18_,
         CARRYB_4__17_, CARRYB_4__16_, CARRYB_4__15_, CARRYB_4__14_,
         CARRYB_4__13_, CARRYB_4__12_, CARRYB_4__11_, CARRYB_4__10_,
         CARRYB_4__9_, CARRYB_4__8_, CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__22_, CARRYB_3__21_, CARRYB_3__20_, CARRYB_3__19_,
         CARRYB_3__18_, CARRYB_3__17_, CARRYB_3__16_, CARRYB_3__15_,
         CARRYB_3__14_, CARRYB_3__13_, CARRYB_3__12_, CARRYB_3__11_,
         CARRYB_3__10_, CARRYB_3__9_, CARRYB_3__8_, CARRYB_3__7_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__22_, CARRYB_2__21_, CARRYB_2__20_,
         CARRYB_2__19_, CARRYB_2__18_, CARRYB_2__17_, CARRYB_2__16_,
         CARRYB_2__15_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__22_,
         CARRYB_1__21_, CARRYB_1__20_, CARRYB_1__19_, CARRYB_1__18_,
         CARRYB_1__17_, CARRYB_1__16_, CARRYB_1__15_, CARRYB_1__14_,
         CARRYB_1__13_, CARRYB_1__12_, CARRYB_1__11_, CARRYB_1__10_,
         CARRYB_1__9_, CARRYB_1__8_, CARRYB_1__7_, CARRYB_1__6_, CARRYB_1__5_,
         CARRYB_1__4_, CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_,
         SUMB_23__23_, SUMB_23__22_, SUMB_23__21_, SUMB_23__20_, SUMB_23__19_,
         SUMB_23__18_, SUMB_23__17_, SUMB_23__16_, SUMB_23__15_, SUMB_23__14_,
         SUMB_23__13_, SUMB_23__12_, SUMB_23__11_, SUMB_23__10_, SUMB_23__9_,
         SUMB_23__8_, SUMB_23__7_, SUMB_23__6_, SUMB_23__5_, SUMB_23__4_,
         SUMB_23__3_, SUMB_23__2_, SUMB_23__1_, SUMB_23__0_, SUMB_22__22_,
         SUMB_22__21_, SUMB_22__20_, SUMB_22__19_, SUMB_22__18_, SUMB_22__17_,
         SUMB_22__16_, SUMB_22__15_, SUMB_22__14_, SUMB_22__13_, SUMB_22__12_,
         SUMB_22__11_, SUMB_22__10_, SUMB_22__9_, SUMB_22__8_, SUMB_22__7_,
         SUMB_22__6_, SUMB_22__5_, SUMB_22__4_, SUMB_22__3_, SUMB_22__2_,
         SUMB_22__1_, SUMB_21__22_, SUMB_21__21_, SUMB_21__20_, SUMB_21__19_,
         SUMB_21__18_, SUMB_21__17_, SUMB_21__16_, SUMB_21__15_, SUMB_21__14_,
         SUMB_21__13_, SUMB_21__12_, SUMB_21__11_, SUMB_21__10_, SUMB_21__9_,
         SUMB_21__8_, SUMB_21__7_, SUMB_21__6_, SUMB_21__5_, SUMB_21__4_,
         SUMB_21__3_, SUMB_21__2_, SUMB_21__1_, SUMB_20__22_, SUMB_20__21_,
         SUMB_20__20_, SUMB_20__19_, SUMB_20__18_, SUMB_20__17_, SUMB_20__16_,
         SUMB_20__15_, SUMB_20__14_, SUMB_20__13_, SUMB_20__12_, SUMB_20__11_,
         SUMB_20__10_, SUMB_20__9_, SUMB_20__8_, SUMB_20__7_, SUMB_20__6_,
         SUMB_20__5_, SUMB_20__4_, SUMB_20__3_, SUMB_20__2_, SUMB_20__1_,
         SUMB_19__22_, SUMB_19__21_, SUMB_19__20_, SUMB_19__19_, SUMB_19__18_,
         SUMB_19__17_, SUMB_19__16_, SUMB_19__15_, SUMB_19__14_, SUMB_19__13_,
         SUMB_19__12_, SUMB_19__11_, SUMB_19__10_, SUMB_19__9_, SUMB_19__8_,
         SUMB_19__7_, SUMB_19__6_, SUMB_19__5_, SUMB_19__4_, SUMB_19__3_,
         SUMB_19__2_, SUMB_19__1_, SUMB_18__22_, SUMB_18__21_, SUMB_18__20_,
         SUMB_18__19_, SUMB_18__18_, SUMB_18__17_, SUMB_18__16_, SUMB_18__15_,
         SUMB_18__14_, SUMB_18__13_, SUMB_18__12_, SUMB_18__11_, SUMB_18__10_,
         SUMB_18__9_, SUMB_18__8_, SUMB_18__7_, SUMB_18__6_, SUMB_18__5_,
         SUMB_18__4_, SUMB_18__3_, SUMB_18__2_, SUMB_18__1_, SUMB_17__22_,
         SUMB_17__21_, SUMB_17__20_, SUMB_17__19_, SUMB_17__18_, SUMB_17__17_,
         SUMB_17__16_, SUMB_17__15_, SUMB_17__14_, SUMB_17__13_, SUMB_17__12_,
         SUMB_17__11_, SUMB_17__10_, SUMB_17__9_, SUMB_17__8_, SUMB_17__7_,
         SUMB_17__6_, SUMB_17__5_, SUMB_17__4_, SUMB_17__3_, SUMB_17__2_,
         SUMB_17__1_, SUMB_16__22_, SUMB_16__21_, SUMB_16__20_, SUMB_16__19_,
         SUMB_16__18_, SUMB_16__17_, SUMB_16__16_, SUMB_16__15_, SUMB_16__14_,
         SUMB_16__13_, SUMB_16__12_, SUMB_16__11_, SUMB_16__10_, SUMB_16__9_,
         SUMB_16__8_, SUMB_16__7_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_,
         SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, SUMB_15__22_, SUMB_15__21_,
         SUMB_15__20_, SUMB_15__19_, SUMB_15__18_, SUMB_15__17_, SUMB_15__16_,
         SUMB_15__15_, SUMB_15__14_, SUMB_15__13_, SUMB_15__12_, SUMB_15__11_,
         SUMB_15__10_, SUMB_15__9_, SUMB_15__8_, SUMB_15__7_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_14__22_, SUMB_14__21_, SUMB_14__20_, SUMB_14__19_, SUMB_14__18_,
         SUMB_14__17_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_, SUMB_14__13_,
         SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_, SUMB_14__8_,
         SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_,
         SUMB_14__2_, SUMB_14__1_, SUMB_13__22_, SUMB_13__21_, SUMB_13__20_,
         SUMB_13__19_, SUMB_13__18_, SUMB_13__17_, SUMB_13__16_, SUMB_13__15_,
         SUMB_13__14_, SUMB_13__13_, SUMB_13__12_, SUMB_13__11_, SUMB_13__10_,
         SUMB_13__9_, SUMB_13__8_, SUMB_13__7_, SUMB_13__6_, SUMB_13__5_,
         SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_, SUMB_12__22_,
         SUMB_12__21_, SUMB_12__20_, SUMB_12__19_, SUMB_12__18_, SUMB_12__17_,
         SUMB_12__16_, SUMB_12__15_, SUMB_12__14_, SUMB_12__13_, SUMB_12__12_,
         SUMB_12__11_, SUMB_12__10_, SUMB_12__9_, SUMB_12__8_, SUMB_12__7_,
         SUMB_12__6_, SUMB_12__5_, SUMB_12__4_, SUMB_12__3_, SUMB_12__2_,
         SUMB_12__1_, SUMB_11__22_, SUMB_11__21_, SUMB_11__20_, SUMB_11__19_,
         SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_, SUMB_11__14_,
         SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_, SUMB_11__9_,
         SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_, SUMB_11__4_,
         SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__22_, SUMB_10__21_,
         SUMB_10__20_, SUMB_10__19_, SUMB_10__18_, SUMB_10__17_, SUMB_10__16_,
         SUMB_10__15_, SUMB_10__14_, SUMB_10__13_, SUMB_10__12_, SUMB_10__11_,
         SUMB_10__10_, SUMB_10__9_, SUMB_10__8_, SUMB_10__7_, SUMB_10__6_,
         SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_,
         SUMB_9__22_, SUMB_9__21_, SUMB_9__20_, SUMB_9__19_, SUMB_9__18_,
         SUMB_9__17_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_, SUMB_9__13_,
         SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_, SUMB_9__8_,
         SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_,
         SUMB_9__2_, SUMB_9__1_, SUMB_8__22_, SUMB_8__21_, SUMB_8__20_,
         SUMB_8__19_, SUMB_8__18_, SUMB_8__17_, SUMB_8__16_, SUMB_8__15_,
         SUMB_8__14_, SUMB_8__13_, SUMB_8__12_, SUMB_8__11_, SUMB_8__10_,
         SUMB_8__9_, SUMB_8__8_, SUMB_8__7_, SUMB_8__6_, SUMB_8__5_,
         SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_, SUMB_7__22_,
         SUMB_7__21_, SUMB_7__20_, SUMB_7__19_, SUMB_7__18_, SUMB_7__17_,
         SUMB_7__16_, SUMB_7__15_, SUMB_7__14_, SUMB_7__13_, SUMB_7__12_,
         SUMB_7__11_, SUMB_7__10_, SUMB_7__9_, SUMB_7__8_, SUMB_7__7_,
         SUMB_7__6_, SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_,
         SUMB_7__1_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_, SUMB_6__19_,
         SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_, SUMB_6__14_,
         SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_, SUMB_6__9_,
         SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_,
         SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__22_, SUMB_5__21_,
         SUMB_5__20_, SUMB_5__19_, SUMB_5__18_, SUMB_5__17_, SUMB_5__16_,
         SUMB_5__15_, SUMB_5__14_, SUMB_5__13_, SUMB_5__12_, SUMB_5__11_,
         SUMB_5__10_, SUMB_5__9_, SUMB_5__8_, SUMB_5__7_, SUMB_5__6_,
         SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_,
         SUMB_4__22_, SUMB_4__21_, SUMB_4__20_, SUMB_4__19_, SUMB_4__18_,
         SUMB_4__17_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_, SUMB_4__13_,
         SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_, SUMB_4__8_,
         SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_,
         SUMB_4__2_, SUMB_4__1_, SUMB_3__22_, SUMB_3__21_, SUMB_3__20_,
         SUMB_3__19_, SUMB_3__18_, SUMB_3__17_, SUMB_3__16_, SUMB_3__15_,
         SUMB_3__14_, SUMB_3__13_, SUMB_3__12_, SUMB_3__11_, SUMB_3__10_,
         SUMB_3__9_, SUMB_3__8_, SUMB_3__7_, SUMB_3__6_, SUMB_3__5_,
         SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_, SUMB_2__22_,
         SUMB_2__21_, SUMB_2__20_, SUMB_2__19_, SUMB_2__18_, SUMB_2__17_,
         SUMB_2__16_, SUMB_2__15_, SUMB_2__14_, SUMB_2__13_, SUMB_2__12_,
         SUMB_2__11_, SUMB_2__10_, SUMB_2__9_, SUMB_2__8_, SUMB_2__7_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__22_, SUMB_1__21_, SUMB_1__20_, SUMB_1__19_,
         SUMB_1__18_, SUMB_1__17_, SUMB_1__16_, SUMB_1__15_, SUMB_1__14_,
         SUMB_1__13_, SUMB_1__12_, SUMB_1__11_, SUMB_1__10_, SUMB_1__9_,
         SUMB_1__8_, SUMB_1__7_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_,
         SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, QA, QB, A1_45_, A1_44_, A1_43_,
         A1_42_, A1_41_, A1_40_, A1_39_, A1_38_, A1_37_, A1_36_, A1_35_,
         A1_34_, A1_33_, A1_32_, A1_31_, A1_30_, A1_29_, A1_28_, A1_27_,
         A1_26_, A1_25_, A1_24_, A1_23_, A1_22_, A1_21_, A1_20_, A1_19_,
         A1_18_, A1_17_, A1_16_, A1_15_, A1_14_, A1_13_, A1_12_, A1_11_,
         A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_,
         A1_0_, A2_45_, A2_44_, A2_43_, A2_42_, A2_41_, A2_40_, A2_39_, A2_38_,
         A2_37_, A2_36_, A2_35_, A2_34_, A2_33_, A2_32_, A2_31_, A2_30_,
         A2_29_, A2_28_, A2_27_, A2_26_, A2_25_, A2_24_, A2_23_, A2_22_, n1,
         n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21;

  FA_X1 S14_23_0 ( .A(A[23]), .B(B[23]), .CI(SUMB_23__0_), .CO(A2_22_), .S(
        A1_21_) );
  FA_X1 S4_0 ( .A(ab_23__0_), .B(CARRYB_22__0_), .CI(SUMB_22__1_), .CO(
        CARRYB_23__0_), .S(SUMB_23__0_) );
  FA_X1 S4_1 ( .A(ab_23__1_), .B(CARRYB_22__1_), .CI(SUMB_22__2_), .CO(
        CARRYB_23__1_), .S(SUMB_23__1_) );
  FA_X1 S4_2 ( .A(ab_23__2_), .B(CARRYB_22__2_), .CI(SUMB_22__3_), .CO(
        CARRYB_23__2_), .S(SUMB_23__2_) );
  FA_X1 S4_3 ( .A(ab_23__3_), .B(CARRYB_22__3_), .CI(SUMB_22__4_), .CO(
        CARRYB_23__3_), .S(SUMB_23__3_) );
  FA_X1 S4_4 ( .A(ab_23__4_), .B(CARRYB_22__4_), .CI(SUMB_22__5_), .CO(
        CARRYB_23__4_), .S(SUMB_23__4_) );
  FA_X1 S4_5 ( .A(ab_23__5_), .B(CARRYB_22__5_), .CI(SUMB_22__6_), .CO(
        CARRYB_23__5_), .S(SUMB_23__5_) );
  FA_X1 S4_6 ( .A(ab_23__6_), .B(CARRYB_22__6_), .CI(SUMB_22__7_), .CO(
        CARRYB_23__6_), .S(SUMB_23__6_) );
  FA_X1 S4_7 ( .A(ab_23__7_), .B(CARRYB_22__7_), .CI(SUMB_22__8_), .CO(
        CARRYB_23__7_), .S(SUMB_23__7_) );
  FA_X1 S4_8 ( .A(ab_23__8_), .B(CARRYB_22__8_), .CI(SUMB_22__9_), .CO(
        CARRYB_23__8_), .S(SUMB_23__8_) );
  FA_X1 S4_9 ( .A(ab_23__9_), .B(CARRYB_22__9_), .CI(SUMB_22__10_), .CO(
        CARRYB_23__9_), .S(SUMB_23__9_) );
  FA_X1 S4_10 ( .A(ab_23__10_), .B(CARRYB_22__10_), .CI(SUMB_22__11_), .CO(
        CARRYB_23__10_), .S(SUMB_23__10_) );
  FA_X1 S4_11 ( .A(ab_23__11_), .B(CARRYB_22__11_), .CI(SUMB_22__12_), .CO(
        CARRYB_23__11_), .S(SUMB_23__11_) );
  FA_X1 S4_12 ( .A(ab_23__12_), .B(CARRYB_22__12_), .CI(SUMB_22__13_), .CO(
        CARRYB_23__12_), .S(SUMB_23__12_) );
  FA_X1 S4_13 ( .A(ab_23__13_), .B(CARRYB_22__13_), .CI(SUMB_22__14_), .CO(
        CARRYB_23__13_), .S(SUMB_23__13_) );
  FA_X1 S4_14 ( .A(ab_23__14_), .B(CARRYB_22__14_), .CI(SUMB_22__15_), .CO(
        CARRYB_23__14_), .S(SUMB_23__14_) );
  FA_X1 S4_15 ( .A(ab_23__15_), .B(CARRYB_22__15_), .CI(SUMB_22__16_), .CO(
        CARRYB_23__15_), .S(SUMB_23__15_) );
  FA_X1 S4_16 ( .A(ab_23__16_), .B(CARRYB_22__16_), .CI(SUMB_22__17_), .CO(
        CARRYB_23__16_), .S(SUMB_23__16_) );
  FA_X1 S4_17 ( .A(ab_23__17_), .B(CARRYB_22__17_), .CI(SUMB_22__18_), .CO(
        CARRYB_23__17_), .S(SUMB_23__17_) );
  FA_X1 S4_18 ( .A(ab_23__18_), .B(CARRYB_22__18_), .CI(SUMB_22__19_), .CO(
        CARRYB_23__18_), .S(SUMB_23__18_) );
  FA_X1 S4_19 ( .A(ab_23__19_), .B(CARRYB_22__19_), .CI(SUMB_22__20_), .CO(
        CARRYB_23__19_), .S(SUMB_23__19_) );
  FA_X1 S4_20 ( .A(ab_23__20_), .B(CARRYB_22__20_), .CI(SUMB_22__21_), .CO(
        CARRYB_23__20_), .S(SUMB_23__20_) );
  FA_X1 S4_21 ( .A(ab_23__21_), .B(CARRYB_22__21_), .CI(SUMB_22__22_), .CO(
        CARRYB_23__21_), .S(SUMB_23__21_) );
  FA_X1 S5_22 ( .A(ab_23__22_), .B(CARRYB_22__22_), .CI(ab_22__23_), .CO(
        CARRYB_23__22_), .S(SUMB_23__22_) );
  FA_X1 S14_23 ( .A(n3), .B(n1), .CI(ab_23__23_), .CO(CARRYB_23__23_), .S(
        SUMB_23__23_) );
  FA_X1 S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), .CO(
        CARRYB_22__0_), .S(A1_20_) );
  FA_X1 S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), .CO(
        CARRYB_22__1_), .S(SUMB_22__1_) );
  FA_X1 S2_22_2 ( .A(ab_22__2_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), .CO(
        CARRYB_22__2_), .S(SUMB_22__2_) );
  FA_X1 S2_22_3 ( .A(ab_22__3_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), .CO(
        CARRYB_22__3_), .S(SUMB_22__3_) );
  FA_X1 S2_22_4 ( .A(ab_22__4_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), .CO(
        CARRYB_22__4_), .S(SUMB_22__4_) );
  FA_X1 S2_22_5 ( .A(ab_22__5_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), .CO(
        CARRYB_22__5_), .S(SUMB_22__5_) );
  FA_X1 S2_22_6 ( .A(ab_22__6_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), .CO(
        CARRYB_22__6_), .S(SUMB_22__6_) );
  FA_X1 S2_22_7 ( .A(ab_22__7_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), .CO(
        CARRYB_22__7_), .S(SUMB_22__7_) );
  FA_X1 S2_22_8 ( .A(ab_22__8_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), .CO(
        CARRYB_22__8_), .S(SUMB_22__8_) );
  FA_X1 S2_22_9 ( .A(ab_22__9_), .B(CARRYB_21__9_), .CI(SUMB_21__10_), .CO(
        CARRYB_22__9_), .S(SUMB_22__9_) );
  FA_X1 S2_22_10 ( .A(ab_22__10_), .B(CARRYB_21__10_), .CI(SUMB_21__11_), .CO(
        CARRYB_22__10_), .S(SUMB_22__10_) );
  FA_X1 S2_22_11 ( .A(ab_22__11_), .B(CARRYB_21__11_), .CI(SUMB_21__12_), .CO(
        CARRYB_22__11_), .S(SUMB_22__11_) );
  FA_X1 S2_22_12 ( .A(ab_22__12_), .B(CARRYB_21__12_), .CI(SUMB_21__13_), .CO(
        CARRYB_22__12_), .S(SUMB_22__12_) );
  FA_X1 S2_22_13 ( .A(ab_22__13_), .B(CARRYB_21__13_), .CI(SUMB_21__14_), .CO(
        CARRYB_22__13_), .S(SUMB_22__13_) );
  FA_X1 S2_22_14 ( .A(ab_22__14_), .B(CARRYB_21__14_), .CI(SUMB_21__15_), .CO(
        CARRYB_22__14_), .S(SUMB_22__14_) );
  FA_X1 S2_22_15 ( .A(ab_22__15_), .B(CARRYB_21__15_), .CI(SUMB_21__16_), .CO(
        CARRYB_22__15_), .S(SUMB_22__15_) );
  FA_X1 S2_22_16 ( .A(ab_22__16_), .B(CARRYB_21__16_), .CI(SUMB_21__17_), .CO(
        CARRYB_22__16_), .S(SUMB_22__16_) );
  FA_X1 S2_22_17 ( .A(ab_22__17_), .B(CARRYB_21__17_), .CI(SUMB_21__18_), .CO(
        CARRYB_22__17_), .S(SUMB_22__17_) );
  FA_X1 S2_22_18 ( .A(ab_22__18_), .B(CARRYB_21__18_), .CI(SUMB_21__19_), .CO(
        CARRYB_22__18_), .S(SUMB_22__18_) );
  FA_X1 S2_22_19 ( .A(ab_22__19_), .B(CARRYB_21__19_), .CI(SUMB_21__20_), .CO(
        CARRYB_22__19_), .S(SUMB_22__19_) );
  FA_X1 S2_22_20 ( .A(ab_22__20_), .B(CARRYB_21__20_), .CI(SUMB_21__21_), .CO(
        CARRYB_22__20_), .S(SUMB_22__20_) );
  FA_X1 S2_22_21 ( .A(ab_22__21_), .B(CARRYB_21__21_), .CI(SUMB_21__22_), .CO(
        CARRYB_22__21_), .S(SUMB_22__21_) );
  FA_X1 S3_22_22 ( .A(ab_22__22_), .B(CARRYB_21__22_), .CI(ab_21__23_), .CO(
        CARRYB_22__22_), .S(SUMB_22__22_) );
  FA_X1 S1_21_0 ( .A(ab_21__0_), .B(CARRYB_20__0_), .CI(SUMB_20__1_), .CO(
        CARRYB_21__0_), .S(A1_19_) );
  FA_X1 S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), .CO(
        CARRYB_21__1_), .S(SUMB_21__1_) );
  FA_X1 S2_21_2 ( .A(ab_21__2_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), .CO(
        CARRYB_21__2_), .S(SUMB_21__2_) );
  FA_X1 S2_21_3 ( .A(ab_21__3_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), .CO(
        CARRYB_21__3_), .S(SUMB_21__3_) );
  FA_X1 S2_21_4 ( .A(ab_21__4_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), .CO(
        CARRYB_21__4_), .S(SUMB_21__4_) );
  FA_X1 S2_21_5 ( .A(ab_21__5_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), .CO(
        CARRYB_21__5_), .S(SUMB_21__5_) );
  FA_X1 S2_21_6 ( .A(ab_21__6_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), .CO(
        CARRYB_21__6_), .S(SUMB_21__6_) );
  FA_X1 S2_21_7 ( .A(ab_21__7_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), .CO(
        CARRYB_21__7_), .S(SUMB_21__7_) );
  FA_X1 S2_21_8 ( .A(ab_21__8_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), .CO(
        CARRYB_21__8_), .S(SUMB_21__8_) );
  FA_X1 S2_21_9 ( .A(ab_21__9_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), .CO(
        CARRYB_21__9_), .S(SUMB_21__9_) );
  FA_X1 S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .CI(SUMB_20__11_), .CO(
        CARRYB_21__10_), .S(SUMB_21__10_) );
  FA_X1 S2_21_11 ( .A(ab_21__11_), .B(CARRYB_20__11_), .CI(SUMB_20__12_), .CO(
        CARRYB_21__11_), .S(SUMB_21__11_) );
  FA_X1 S2_21_12 ( .A(ab_21__12_), .B(CARRYB_20__12_), .CI(SUMB_20__13_), .CO(
        CARRYB_21__12_), .S(SUMB_21__12_) );
  FA_X1 S2_21_13 ( .A(ab_21__13_), .B(CARRYB_20__13_), .CI(SUMB_20__14_), .CO(
        CARRYB_21__13_), .S(SUMB_21__13_) );
  FA_X1 S2_21_14 ( .A(ab_21__14_), .B(CARRYB_20__14_), .CI(SUMB_20__15_), .CO(
        CARRYB_21__14_), .S(SUMB_21__14_) );
  FA_X1 S2_21_15 ( .A(ab_21__15_), .B(CARRYB_20__15_), .CI(SUMB_20__16_), .CO(
        CARRYB_21__15_), .S(SUMB_21__15_) );
  FA_X1 S2_21_16 ( .A(ab_21__16_), .B(CARRYB_20__16_), .CI(SUMB_20__17_), .CO(
        CARRYB_21__16_), .S(SUMB_21__16_) );
  FA_X1 S2_21_17 ( .A(ab_21__17_), .B(CARRYB_20__17_), .CI(SUMB_20__18_), .CO(
        CARRYB_21__17_), .S(SUMB_21__17_) );
  FA_X1 S2_21_18 ( .A(ab_21__18_), .B(CARRYB_20__18_), .CI(SUMB_20__19_), .CO(
        CARRYB_21__18_), .S(SUMB_21__18_) );
  FA_X1 S2_21_19 ( .A(ab_21__19_), .B(CARRYB_20__19_), .CI(SUMB_20__20_), .CO(
        CARRYB_21__19_), .S(SUMB_21__19_) );
  FA_X1 S2_21_20 ( .A(ab_21__20_), .B(CARRYB_20__20_), .CI(SUMB_20__21_), .CO(
        CARRYB_21__20_), .S(SUMB_21__20_) );
  FA_X1 S2_21_21 ( .A(ab_21__21_), .B(CARRYB_20__21_), .CI(SUMB_20__22_), .CO(
        CARRYB_21__21_), .S(SUMB_21__21_) );
  FA_X1 S3_21_22 ( .A(ab_21__22_), .B(CARRYB_20__22_), .CI(ab_20__23_), .CO(
        CARRYB_21__22_), .S(SUMB_21__22_) );
  FA_X1 S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), .CO(
        CARRYB_20__0_), .S(A1_18_) );
  FA_X1 S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), .CO(
        CARRYB_20__1_), .S(SUMB_20__1_) );
  FA_X1 S2_20_2 ( .A(ab_20__2_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), .CO(
        CARRYB_20__2_), .S(SUMB_20__2_) );
  FA_X1 S2_20_3 ( .A(ab_20__3_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), .CO(
        CARRYB_20__3_), .S(SUMB_20__3_) );
  FA_X1 S2_20_4 ( .A(ab_20__4_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), .CO(
        CARRYB_20__4_), .S(SUMB_20__4_) );
  FA_X1 S2_20_5 ( .A(ab_20__5_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), .CO(
        CARRYB_20__5_), .S(SUMB_20__5_) );
  FA_X1 S2_20_6 ( .A(ab_20__6_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), .CO(
        CARRYB_20__6_), .S(SUMB_20__6_) );
  FA_X1 S2_20_7 ( .A(ab_20__7_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), .CO(
        CARRYB_20__7_), .S(SUMB_20__7_) );
  FA_X1 S2_20_8 ( .A(ab_20__8_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), .CO(
        CARRYB_20__8_), .S(SUMB_20__8_) );
  FA_X1 S2_20_9 ( .A(ab_20__9_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), .CO(
        CARRYB_20__9_), .S(SUMB_20__9_) );
  FA_X1 S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), .CO(
        CARRYB_20__10_), .S(SUMB_20__10_) );
  FA_X1 S2_20_11 ( .A(ab_20__11_), .B(CARRYB_19__11_), .CI(SUMB_19__12_), .CO(
        CARRYB_20__11_), .S(SUMB_20__11_) );
  FA_X1 S2_20_12 ( .A(ab_20__12_), .B(CARRYB_19__12_), .CI(SUMB_19__13_), .CO(
        CARRYB_20__12_), .S(SUMB_20__12_) );
  FA_X1 S2_20_13 ( .A(ab_20__13_), .B(CARRYB_19__13_), .CI(SUMB_19__14_), .CO(
        CARRYB_20__13_), .S(SUMB_20__13_) );
  FA_X1 S2_20_14 ( .A(ab_20__14_), .B(CARRYB_19__14_), .CI(SUMB_19__15_), .CO(
        CARRYB_20__14_), .S(SUMB_20__14_) );
  FA_X1 S2_20_15 ( .A(ab_20__15_), .B(CARRYB_19__15_), .CI(SUMB_19__16_), .CO(
        CARRYB_20__15_), .S(SUMB_20__15_) );
  FA_X1 S2_20_16 ( .A(ab_20__16_), .B(CARRYB_19__16_), .CI(SUMB_19__17_), .CO(
        CARRYB_20__16_), .S(SUMB_20__16_) );
  FA_X1 S2_20_17 ( .A(ab_20__17_), .B(CARRYB_19__17_), .CI(SUMB_19__18_), .CO(
        CARRYB_20__17_), .S(SUMB_20__17_) );
  FA_X1 S2_20_18 ( .A(ab_20__18_), .B(CARRYB_19__18_), .CI(SUMB_19__19_), .CO(
        CARRYB_20__18_), .S(SUMB_20__18_) );
  FA_X1 S2_20_19 ( .A(ab_20__19_), .B(CARRYB_19__19_), .CI(SUMB_19__20_), .CO(
        CARRYB_20__19_), .S(SUMB_20__19_) );
  FA_X1 S2_20_20 ( .A(ab_20__20_), .B(CARRYB_19__20_), .CI(SUMB_19__21_), .CO(
        CARRYB_20__20_), .S(SUMB_20__20_) );
  FA_X1 S2_20_21 ( .A(ab_20__21_), .B(CARRYB_19__21_), .CI(SUMB_19__22_), .CO(
        CARRYB_20__21_), .S(SUMB_20__21_) );
  FA_X1 S3_20_22 ( .A(ab_20__22_), .B(CARRYB_19__22_), .CI(ab_19__23_), .CO(
        CARRYB_20__22_), .S(SUMB_20__22_) );
  FA_X1 S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), .CO(
        CARRYB_19__0_), .S(A1_17_) );
  FA_X1 S2_19_1 ( .A(ab_19__1_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), .CO(
        CARRYB_19__1_), .S(SUMB_19__1_) );
  FA_X1 S2_19_2 ( .A(ab_19__2_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), .CO(
        CARRYB_19__2_), .S(SUMB_19__2_) );
  FA_X1 S2_19_3 ( .A(ab_19__3_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), .CO(
        CARRYB_19__3_), .S(SUMB_19__3_) );
  FA_X1 S2_19_4 ( .A(ab_19__4_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), .CO(
        CARRYB_19__4_), .S(SUMB_19__4_) );
  FA_X1 S2_19_5 ( .A(ab_19__5_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), .CO(
        CARRYB_19__5_), .S(SUMB_19__5_) );
  FA_X1 S2_19_6 ( .A(ab_19__6_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), .CO(
        CARRYB_19__6_), .S(SUMB_19__6_) );
  FA_X1 S2_19_7 ( .A(ab_19__7_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), .CO(
        CARRYB_19__7_), .S(SUMB_19__7_) );
  FA_X1 S2_19_8 ( .A(ab_19__8_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), .CO(
        CARRYB_19__8_), .S(SUMB_19__8_) );
  FA_X1 S2_19_9 ( .A(ab_19__9_), .B(CARRYB_18__9_), .CI(SUMB_18__10_), .CO(
        CARRYB_19__9_), .S(SUMB_19__9_) );
  FA_X1 S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), .CO(
        CARRYB_19__10_), .S(SUMB_19__10_) );
  FA_X1 S2_19_11 ( .A(ab_19__11_), .B(CARRYB_18__11_), .CI(SUMB_18__12_), .CO(
        CARRYB_19__11_), .S(SUMB_19__11_) );
  FA_X1 S2_19_12 ( .A(ab_19__12_), .B(CARRYB_18__12_), .CI(SUMB_18__13_), .CO(
        CARRYB_19__12_), .S(SUMB_19__12_) );
  FA_X1 S2_19_13 ( .A(ab_19__13_), .B(CARRYB_18__13_), .CI(SUMB_18__14_), .CO(
        CARRYB_19__13_), .S(SUMB_19__13_) );
  FA_X1 S2_19_14 ( .A(ab_19__14_), .B(CARRYB_18__14_), .CI(SUMB_18__15_), .CO(
        CARRYB_19__14_), .S(SUMB_19__14_) );
  FA_X1 S2_19_15 ( .A(ab_19__15_), .B(CARRYB_18__15_), .CI(SUMB_18__16_), .CO(
        CARRYB_19__15_), .S(SUMB_19__15_) );
  FA_X1 S2_19_16 ( .A(ab_19__16_), .B(CARRYB_18__16_), .CI(SUMB_18__17_), .CO(
        CARRYB_19__16_), .S(SUMB_19__16_) );
  FA_X1 S2_19_17 ( .A(ab_19__17_), .B(CARRYB_18__17_), .CI(SUMB_18__18_), .CO(
        CARRYB_19__17_), .S(SUMB_19__17_) );
  FA_X1 S2_19_18 ( .A(ab_19__18_), .B(CARRYB_18__18_), .CI(SUMB_18__19_), .CO(
        CARRYB_19__18_), .S(SUMB_19__18_) );
  FA_X1 S2_19_19 ( .A(ab_19__19_), .B(CARRYB_18__19_), .CI(SUMB_18__20_), .CO(
        CARRYB_19__19_), .S(SUMB_19__19_) );
  FA_X1 S2_19_20 ( .A(ab_19__20_), .B(CARRYB_18__20_), .CI(SUMB_18__21_), .CO(
        CARRYB_19__20_), .S(SUMB_19__20_) );
  FA_X1 S2_19_21 ( .A(ab_19__21_), .B(CARRYB_18__21_), .CI(SUMB_18__22_), .CO(
        CARRYB_19__21_), .S(SUMB_19__21_) );
  FA_X1 S3_19_22 ( .A(ab_19__22_), .B(CARRYB_18__22_), .CI(ab_18__23_), .CO(
        CARRYB_19__22_), .S(SUMB_19__22_) );
  FA_X1 S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), .CO(
        CARRYB_18__0_), .S(A1_16_) );
  FA_X1 S2_18_1 ( .A(ab_18__1_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), .CO(
        CARRYB_18__1_), .S(SUMB_18__1_) );
  FA_X1 S2_18_2 ( .A(ab_18__2_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), .CO(
        CARRYB_18__2_), .S(SUMB_18__2_) );
  FA_X1 S2_18_3 ( .A(ab_18__3_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), .CO(
        CARRYB_18__3_), .S(SUMB_18__3_) );
  FA_X1 S2_18_4 ( .A(ab_18__4_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), .CO(
        CARRYB_18__4_), .S(SUMB_18__4_) );
  FA_X1 S2_18_5 ( .A(ab_18__5_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), .CO(
        CARRYB_18__5_), .S(SUMB_18__5_) );
  FA_X1 S2_18_6 ( .A(ab_18__6_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), .CO(
        CARRYB_18__6_), .S(SUMB_18__6_) );
  FA_X1 S2_18_7 ( .A(ab_18__7_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), .CO(
        CARRYB_18__7_), .S(SUMB_18__7_) );
  FA_X1 S2_18_8 ( .A(ab_18__8_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), .CO(
        CARRYB_18__8_), .S(SUMB_18__8_) );
  FA_X1 S2_18_9 ( .A(ab_18__9_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), .CO(
        CARRYB_18__9_), .S(SUMB_18__9_) );
  FA_X1 S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), .CO(
        CARRYB_18__10_), .S(SUMB_18__10_) );
  FA_X1 S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), .CO(
        CARRYB_18__11_), .S(SUMB_18__11_) );
  FA_X1 S2_18_12 ( .A(ab_18__12_), .B(CARRYB_17__12_), .CI(SUMB_17__13_), .CO(
        CARRYB_18__12_), .S(SUMB_18__12_) );
  FA_X1 S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .CI(SUMB_17__14_), .CO(
        CARRYB_18__13_), .S(SUMB_18__13_) );
  FA_X1 S2_18_14 ( .A(ab_18__14_), .B(CARRYB_17__14_), .CI(SUMB_17__15_), .CO(
        CARRYB_18__14_), .S(SUMB_18__14_) );
  FA_X1 S2_18_15 ( .A(ab_18__15_), .B(CARRYB_17__15_), .CI(SUMB_17__16_), .CO(
        CARRYB_18__15_), .S(SUMB_18__15_) );
  FA_X1 S2_18_16 ( .A(ab_18__16_), .B(CARRYB_17__16_), .CI(SUMB_17__17_), .CO(
        CARRYB_18__16_), .S(SUMB_18__16_) );
  FA_X1 S2_18_17 ( .A(ab_18__17_), .B(CARRYB_17__17_), .CI(SUMB_17__18_), .CO(
        CARRYB_18__17_), .S(SUMB_18__17_) );
  FA_X1 S2_18_18 ( .A(ab_18__18_), .B(CARRYB_17__18_), .CI(SUMB_17__19_), .CO(
        CARRYB_18__18_), .S(SUMB_18__18_) );
  FA_X1 S2_18_19 ( .A(ab_18__19_), .B(CARRYB_17__19_), .CI(SUMB_17__20_), .CO(
        CARRYB_18__19_), .S(SUMB_18__19_) );
  FA_X1 S2_18_20 ( .A(ab_18__20_), .B(CARRYB_17__20_), .CI(SUMB_17__21_), .CO(
        CARRYB_18__20_), .S(SUMB_18__20_) );
  FA_X1 S2_18_21 ( .A(ab_18__21_), .B(CARRYB_17__21_), .CI(SUMB_17__22_), .CO(
        CARRYB_18__21_), .S(SUMB_18__21_) );
  FA_X1 S3_18_22 ( .A(ab_18__22_), .B(CARRYB_17__22_), .CI(ab_17__23_), .CO(
        CARRYB_18__22_), .S(SUMB_18__22_) );
  FA_X1 S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), .CO(
        CARRYB_17__0_), .S(A1_15_) );
  FA_X1 S2_17_1 ( .A(ab_17__1_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), .CO(
        CARRYB_17__1_), .S(SUMB_17__1_) );
  FA_X1 S2_17_2 ( .A(ab_17__2_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), .CO(
        CARRYB_17__2_), .S(SUMB_17__2_) );
  FA_X1 S2_17_3 ( .A(ab_17__3_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), .CO(
        CARRYB_17__3_), .S(SUMB_17__3_) );
  FA_X1 S2_17_4 ( .A(ab_17__4_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), .CO(
        CARRYB_17__4_), .S(SUMB_17__4_) );
  FA_X1 S2_17_5 ( .A(ab_17__5_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), .CO(
        CARRYB_17__5_), .S(SUMB_17__5_) );
  FA_X1 S2_17_6 ( .A(ab_17__6_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), .CO(
        CARRYB_17__6_), .S(SUMB_17__6_) );
  FA_X1 S2_17_7 ( .A(ab_17__7_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), .CO(
        CARRYB_17__7_), .S(SUMB_17__7_) );
  FA_X1 S2_17_8 ( .A(ab_17__8_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), .CO(
        CARRYB_17__8_), .S(SUMB_17__8_) );
  FA_X1 S2_17_9 ( .A(ab_17__9_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), .CO(
        CARRYB_17__9_), .S(SUMB_17__9_) );
  FA_X1 S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), .CO(
        CARRYB_17__10_), .S(SUMB_17__10_) );
  FA_X1 S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), .CO(
        CARRYB_17__11_), .S(SUMB_17__11_) );
  FA_X1 S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), .CO(
        CARRYB_17__12_), .S(SUMB_17__12_) );
  FA_X1 S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), .CO(
        CARRYB_17__13_), .S(SUMB_17__13_) );
  FA_X1 S2_17_14 ( .A(ab_17__14_), .B(CARRYB_16__14_), .CI(SUMB_16__15_), .CO(
        CARRYB_17__14_), .S(SUMB_17__14_) );
  FA_X1 S2_17_15 ( .A(ab_17__15_), .B(CARRYB_16__15_), .CI(SUMB_16__16_), .CO(
        CARRYB_17__15_), .S(SUMB_17__15_) );
  FA_X1 S2_17_16 ( .A(ab_17__16_), .B(CARRYB_16__16_), .CI(SUMB_16__17_), .CO(
        CARRYB_17__16_), .S(SUMB_17__16_) );
  FA_X1 S2_17_17 ( .A(ab_17__17_), .B(CARRYB_16__17_), .CI(SUMB_16__18_), .CO(
        CARRYB_17__17_), .S(SUMB_17__17_) );
  FA_X1 S2_17_18 ( .A(ab_17__18_), .B(CARRYB_16__18_), .CI(SUMB_16__19_), .CO(
        CARRYB_17__18_), .S(SUMB_17__18_) );
  FA_X1 S2_17_19 ( .A(ab_17__19_), .B(CARRYB_16__19_), .CI(SUMB_16__20_), .CO(
        CARRYB_17__19_), .S(SUMB_17__19_) );
  FA_X1 S2_17_20 ( .A(ab_17__20_), .B(CARRYB_16__20_), .CI(SUMB_16__21_), .CO(
        CARRYB_17__20_), .S(SUMB_17__20_) );
  FA_X1 S2_17_21 ( .A(ab_17__21_), .B(CARRYB_16__21_), .CI(SUMB_16__22_), .CO(
        CARRYB_17__21_), .S(SUMB_17__21_) );
  FA_X1 S3_17_22 ( .A(ab_17__22_), .B(CARRYB_16__22_), .CI(ab_16__23_), .CO(
        CARRYB_17__22_), .S(SUMB_17__22_) );
  FA_X1 S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(A1_14_) );
  FA_X1 S2_16_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  FA_X1 S2_16_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  FA_X1 S2_16_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  FA_X1 S2_16_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  FA_X1 S2_16_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  FA_X1 S2_16_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  FA_X1 S2_16_7 ( .A(ab_16__7_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), .CO(
        CARRYB_16__7_), .S(SUMB_16__7_) );
  FA_X1 S2_16_8 ( .A(ab_16__8_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), .CO(
        CARRYB_16__8_), .S(SUMB_16__8_) );
  FA_X1 S2_16_9 ( .A(ab_16__9_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), .CO(
        CARRYB_16__9_), .S(SUMB_16__9_) );
  FA_X1 S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), .CO(
        CARRYB_16__10_), .S(SUMB_16__10_) );
  FA_X1 S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), .CO(
        CARRYB_16__11_), .S(SUMB_16__11_) );
  FA_X1 S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), .CO(
        CARRYB_16__12_), .S(SUMB_16__12_) );
  FA_X1 S2_16_13 ( .A(ab_16__13_), .B(CARRYB_15__13_), .CI(SUMB_15__14_), .CO(
        CARRYB_16__13_), .S(SUMB_16__13_) );
  FA_X1 S2_16_14 ( .A(ab_16__14_), .B(CARRYB_15__14_), .CI(SUMB_15__15_), .CO(
        CARRYB_16__14_), .S(SUMB_16__14_) );
  FA_X1 S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .CI(SUMB_15__16_), .CO(
        CARRYB_16__15_), .S(SUMB_16__15_) );
  FA_X1 S2_16_16 ( .A(ab_16__16_), .B(CARRYB_15__16_), .CI(SUMB_15__17_), .CO(
        CARRYB_16__16_), .S(SUMB_16__16_) );
  FA_X1 S2_16_17 ( .A(ab_16__17_), .B(CARRYB_15__17_), .CI(SUMB_15__18_), .CO(
        CARRYB_16__17_), .S(SUMB_16__17_) );
  FA_X1 S2_16_18 ( .A(ab_16__18_), .B(CARRYB_15__18_), .CI(SUMB_15__19_), .CO(
        CARRYB_16__18_), .S(SUMB_16__18_) );
  FA_X1 S2_16_19 ( .A(ab_16__19_), .B(CARRYB_15__19_), .CI(SUMB_15__20_), .CO(
        CARRYB_16__19_), .S(SUMB_16__19_) );
  FA_X1 S2_16_20 ( .A(ab_16__20_), .B(CARRYB_15__20_), .CI(SUMB_15__21_), .CO(
        CARRYB_16__20_), .S(SUMB_16__20_) );
  FA_X1 S2_16_21 ( .A(ab_16__21_), .B(CARRYB_15__21_), .CI(SUMB_15__22_), .CO(
        CARRYB_16__21_), .S(SUMB_16__21_) );
  FA_X1 S3_16_22 ( .A(ab_16__22_), .B(CARRYB_15__22_), .CI(ab_15__23_), .CO(
        CARRYB_16__22_), .S(SUMB_16__22_) );
  FA_X1 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  FA_X1 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  FA_X1 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  FA_X1 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  FA_X1 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  FA_X1 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  FA_X1 S2_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  FA_X1 S2_15_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), .CO(
        CARRYB_15__7_), .S(SUMB_15__7_) );
  FA_X1 S2_15_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), .CO(
        CARRYB_15__8_), .S(SUMB_15__8_) );
  FA_X1 S2_15_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), .CO(
        CARRYB_15__9_), .S(SUMB_15__9_) );
  FA_X1 S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), .CO(
        CARRYB_15__10_), .S(SUMB_15__10_) );
  FA_X1 S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), .CO(
        CARRYB_15__11_), .S(SUMB_15__11_) );
  FA_X1 S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), .CO(
        CARRYB_15__12_), .S(SUMB_15__12_) );
  FA_X1 S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), .CO(
        CARRYB_15__13_), .S(SUMB_15__13_) );
  FA_X1 S2_15_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), .CO(
        CARRYB_15__14_), .S(SUMB_15__14_) );
  FA_X1 S2_15_15 ( .A(ab_15__15_), .B(CARRYB_14__15_), .CI(SUMB_14__16_), .CO(
        CARRYB_15__15_), .S(SUMB_15__15_) );
  FA_X1 S2_15_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .CI(SUMB_14__17_), .CO(
        CARRYB_15__16_), .S(SUMB_15__16_) );
  FA_X1 S2_15_17 ( .A(ab_15__17_), .B(CARRYB_14__17_), .CI(SUMB_14__18_), .CO(
        CARRYB_15__17_), .S(SUMB_15__17_) );
  FA_X1 S2_15_18 ( .A(ab_15__18_), .B(CARRYB_14__18_), .CI(SUMB_14__19_), .CO(
        CARRYB_15__18_), .S(SUMB_15__18_) );
  FA_X1 S2_15_19 ( .A(ab_15__19_), .B(CARRYB_14__19_), .CI(SUMB_14__20_), .CO(
        CARRYB_15__19_), .S(SUMB_15__19_) );
  FA_X1 S2_15_20 ( .A(ab_15__20_), .B(CARRYB_14__20_), .CI(SUMB_14__21_), .CO(
        CARRYB_15__20_), .S(SUMB_15__20_) );
  FA_X1 S2_15_21 ( .A(ab_15__21_), .B(CARRYB_14__21_), .CI(SUMB_14__22_), .CO(
        CARRYB_15__21_), .S(SUMB_15__21_) );
  FA_X1 S3_15_22 ( .A(ab_15__22_), .B(CARRYB_14__22_), .CI(ab_14__23_), .CO(
        CARRYB_15__22_), .S(SUMB_15__22_) );
  FA_X1 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  FA_X1 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  FA_X1 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  FA_X1 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  FA_X1 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  FA_X1 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  FA_X1 S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  FA_X1 S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), .CO(
        CARRYB_14__7_), .S(SUMB_14__7_) );
  FA_X1 S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), .CO(
        CARRYB_14__8_), .S(SUMB_14__8_) );
  FA_X1 S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), .CO(
        CARRYB_14__9_), .S(SUMB_14__9_) );
  FA_X1 S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), .CO(
        CARRYB_14__10_), .S(SUMB_14__10_) );
  FA_X1 S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), .CO(
        CARRYB_14__11_), .S(SUMB_14__11_) );
  FA_X1 S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), .CO(
        CARRYB_14__12_), .S(SUMB_14__12_) );
  FA_X1 S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), .CO(
        CARRYB_14__13_), .S(SUMB_14__13_) );
  FA_X1 S2_14_14 ( .A(ab_14__14_), .B(CARRYB_13__14_), .CI(SUMB_13__15_), .CO(
        CARRYB_14__14_), .S(SUMB_14__14_) );
  FA_X1 S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), .CO(
        CARRYB_14__15_), .S(SUMB_14__15_) );
  FA_X1 S2_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), .CO(
        CARRYB_14__16_), .S(SUMB_14__16_) );
  FA_X1 S2_14_17 ( .A(ab_14__17_), .B(CARRYB_13__17_), .CI(SUMB_13__18_), .CO(
        CARRYB_14__17_), .S(SUMB_14__17_) );
  FA_X1 S2_14_18 ( .A(ab_14__18_), .B(CARRYB_13__18_), .CI(SUMB_13__19_), .CO(
        CARRYB_14__18_), .S(SUMB_14__18_) );
  FA_X1 S2_14_19 ( .A(ab_14__19_), .B(CARRYB_13__19_), .CI(SUMB_13__20_), .CO(
        CARRYB_14__19_), .S(SUMB_14__19_) );
  FA_X1 S2_14_20 ( .A(ab_14__20_), .B(CARRYB_13__20_), .CI(SUMB_13__21_), .CO(
        CARRYB_14__20_), .S(SUMB_14__20_) );
  FA_X1 S2_14_21 ( .A(ab_14__21_), .B(CARRYB_13__21_), .CI(SUMB_13__22_), .CO(
        CARRYB_14__21_), .S(SUMB_14__21_) );
  FA_X1 S3_14_22 ( .A(ab_14__22_), .B(CARRYB_13__22_), .CI(ab_13__23_), .CO(
        CARRYB_14__22_), .S(SUMB_14__22_) );
  FA_X1 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  FA_X1 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  FA_X1 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  FA_X1 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  FA_X1 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  FA_X1 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  FA_X1 S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  FA_X1 S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), .CO(
        CARRYB_13__7_), .S(SUMB_13__7_) );
  FA_X1 S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), .CO(
        CARRYB_13__8_), .S(SUMB_13__8_) );
  FA_X1 S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), .CO(
        CARRYB_13__9_), .S(SUMB_13__9_) );
  FA_X1 S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), .CO(
        CARRYB_13__10_), .S(SUMB_13__10_) );
  FA_X1 S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), .CO(
        CARRYB_13__11_), .S(SUMB_13__11_) );
  FA_X1 S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), .CO(
        CARRYB_13__12_), .S(SUMB_13__12_) );
  FA_X1 S2_13_13 ( .A(ab_13__13_), .B(CARRYB_12__13_), .CI(SUMB_12__14_), .CO(
        CARRYB_13__13_), .S(SUMB_13__13_) );
  FA_X1 S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), .CO(
        CARRYB_13__14_), .S(SUMB_13__14_) );
  FA_X1 S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), .CO(
        CARRYB_13__15_), .S(SUMB_13__15_) );
  FA_X1 S2_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), .CO(
        CARRYB_13__16_), .S(SUMB_13__16_) );
  FA_X1 S2_13_17 ( .A(ab_13__17_), .B(CARRYB_12__17_), .CI(SUMB_12__18_), .CO(
        CARRYB_13__17_), .S(SUMB_13__17_) );
  FA_X1 S2_13_18 ( .A(ab_13__18_), .B(CARRYB_12__18_), .CI(SUMB_12__19_), .CO(
        CARRYB_13__18_), .S(SUMB_13__18_) );
  FA_X1 S2_13_19 ( .A(ab_13__19_), .B(CARRYB_12__19_), .CI(SUMB_12__20_), .CO(
        CARRYB_13__19_), .S(SUMB_13__19_) );
  FA_X1 S2_13_20 ( .A(ab_13__20_), .B(CARRYB_12__20_), .CI(SUMB_12__21_), .CO(
        CARRYB_13__20_), .S(SUMB_13__20_) );
  FA_X1 S2_13_21 ( .A(ab_13__21_), .B(CARRYB_12__21_), .CI(SUMB_12__22_), .CO(
        CARRYB_13__21_), .S(SUMB_13__21_) );
  FA_X1 S3_13_22 ( .A(ab_13__22_), .B(CARRYB_12__22_), .CI(ab_12__23_), .CO(
        CARRYB_13__22_), .S(SUMB_13__22_) );
  FA_X1 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  FA_X1 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  FA_X1 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  FA_X1 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  FA_X1 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  FA_X1 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  FA_X1 S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  FA_X1 S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), .CO(
        CARRYB_12__7_), .S(SUMB_12__7_) );
  FA_X1 S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), .CO(
        CARRYB_12__8_), .S(SUMB_12__8_) );
  FA_X1 S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), .CO(
        CARRYB_12__9_), .S(SUMB_12__9_) );
  FA_X1 S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), .CO(
        CARRYB_12__10_), .S(SUMB_12__10_) );
  FA_X1 S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), .CO(
        CARRYB_12__11_), .S(SUMB_12__11_) );
  FA_X1 S2_12_12 ( .A(ab_12__12_), .B(CARRYB_11__12_), .CI(SUMB_11__13_), .CO(
        CARRYB_12__12_), .S(SUMB_12__12_) );
  FA_X1 S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), .CO(
        CARRYB_12__13_), .S(SUMB_12__13_) );
  FA_X1 S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), .CO(
        CARRYB_12__14_), .S(SUMB_12__14_) );
  FA_X1 S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), .CO(
        CARRYB_12__15_), .S(SUMB_12__15_) );
  FA_X1 S2_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), .CO(
        CARRYB_12__16_), .S(SUMB_12__16_) );
  FA_X1 S2_12_17 ( .A(ab_12__17_), .B(CARRYB_11__17_), .CI(SUMB_11__18_), .CO(
        CARRYB_12__17_), .S(SUMB_12__17_) );
  FA_X1 S2_12_18 ( .A(ab_12__18_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), .CO(
        CARRYB_12__18_), .S(SUMB_12__18_) );
  FA_X1 S2_12_19 ( .A(ab_12__19_), .B(CARRYB_11__19_), .CI(SUMB_11__20_), .CO(
        CARRYB_12__19_), .S(SUMB_12__19_) );
  FA_X1 S2_12_20 ( .A(ab_12__20_), .B(CARRYB_11__20_), .CI(SUMB_11__21_), .CO(
        CARRYB_12__20_), .S(SUMB_12__20_) );
  FA_X1 S2_12_21 ( .A(ab_12__21_), .B(CARRYB_11__21_), .CI(SUMB_11__22_), .CO(
        CARRYB_12__21_), .S(SUMB_12__21_) );
  FA_X1 S3_12_22 ( .A(ab_12__22_), .B(CARRYB_11__22_), .CI(ab_11__23_), .CO(
        CARRYB_12__22_), .S(SUMB_12__22_) );
  FA_X1 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  FA_X1 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  FA_X1 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  FA_X1 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  FA_X1 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  FA_X1 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  FA_X1 S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  FA_X1 S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), .CO(
        CARRYB_11__7_), .S(SUMB_11__7_) );
  FA_X1 S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), .CO(
        CARRYB_11__8_), .S(SUMB_11__8_) );
  FA_X1 S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), .CO(
        CARRYB_11__9_), .S(SUMB_11__9_) );
  FA_X1 S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), .CO(
        CARRYB_11__10_), .S(SUMB_11__10_) );
  FA_X1 S2_11_11 ( .A(ab_11__11_), .B(CARRYB_10__11_), .CI(SUMB_10__12_), .CO(
        CARRYB_11__11_), .S(SUMB_11__11_) );
  FA_X1 S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), .CO(
        CARRYB_11__12_), .S(SUMB_11__12_) );
  FA_X1 S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), .CO(
        CARRYB_11__13_), .S(SUMB_11__13_) );
  FA_X1 S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), .CO(
        CARRYB_11__14_), .S(SUMB_11__14_) );
  FA_X1 S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), .CO(
        CARRYB_11__15_), .S(SUMB_11__15_) );
  FA_X1 S2_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(SUMB_10__17_), .CO(
        CARRYB_11__16_), .S(SUMB_11__16_) );
  FA_X1 S2_11_17 ( .A(ab_11__17_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), .CO(
        CARRYB_11__17_), .S(SUMB_11__17_) );
  FA_X1 S2_11_18 ( .A(ab_11__18_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), .CO(
        CARRYB_11__18_), .S(SUMB_11__18_) );
  FA_X1 S2_11_19 ( .A(ab_11__19_), .B(CARRYB_10__19_), .CI(SUMB_10__20_), .CO(
        CARRYB_11__19_), .S(SUMB_11__19_) );
  FA_X1 S2_11_20 ( .A(ab_11__20_), .B(CARRYB_10__20_), .CI(SUMB_10__21_), .CO(
        CARRYB_11__20_), .S(SUMB_11__20_) );
  FA_X1 S2_11_21 ( .A(ab_11__21_), .B(CARRYB_10__21_), .CI(SUMB_10__22_), .CO(
        CARRYB_11__21_), .S(SUMB_11__21_) );
  FA_X1 S3_11_22 ( .A(ab_11__22_), .B(CARRYB_10__22_), .CI(ab_10__23_), .CO(
        CARRYB_11__22_), .S(SUMB_11__22_) );
  FA_X1 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  FA_X1 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  FA_X1 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  FA_X1 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  FA_X1 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  FA_X1 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  FA_X1 S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  FA_X1 S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  FA_X1 S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  FA_X1 S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  FA_X1 S2_10_10 ( .A(ab_10__10_), .B(CARRYB_9__10_), .CI(SUMB_9__11_), .CO(
        CARRYB_10__10_), .S(SUMB_10__10_) );
  FA_X1 S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), .CO(
        CARRYB_10__11_), .S(SUMB_10__11_) );
  FA_X1 S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), .CO(
        CARRYB_10__12_), .S(SUMB_10__12_) );
  FA_X1 S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), .CO(
        CARRYB_10__13_), .S(SUMB_10__13_) );
  FA_X1 S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), .CO(
        CARRYB_10__14_), .S(SUMB_10__14_) );
  FA_X1 S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), .CO(
        CARRYB_10__15_), .S(SUMB_10__15_) );
  FA_X1 S2_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), .CO(
        CARRYB_10__16_), .S(SUMB_10__16_) );
  FA_X1 S2_10_17 ( .A(ab_10__17_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), .CO(
        CARRYB_10__17_), .S(SUMB_10__17_) );
  FA_X1 S2_10_18 ( .A(ab_10__18_), .B(CARRYB_9__18_), .CI(SUMB_9__19_), .CO(
        CARRYB_10__18_), .S(SUMB_10__18_) );
  FA_X1 S2_10_19 ( .A(ab_10__19_), .B(CARRYB_9__19_), .CI(SUMB_9__20_), .CO(
        CARRYB_10__19_), .S(SUMB_10__19_) );
  FA_X1 S2_10_20 ( .A(ab_10__20_), .B(CARRYB_9__20_), .CI(SUMB_9__21_), .CO(
        CARRYB_10__20_), .S(SUMB_10__20_) );
  FA_X1 S2_10_21 ( .A(ab_10__21_), .B(CARRYB_9__21_), .CI(SUMB_9__22_), .CO(
        CARRYB_10__21_), .S(SUMB_10__21_) );
  FA_X1 S3_10_22 ( .A(ab_10__22_), .B(CARRYB_9__22_), .CI(ab_9__23_), .CO(
        CARRYB_10__22_), .S(SUMB_10__22_) );
  FA_X1 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  FA_X1 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  FA_X1 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  FA_X1 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  FA_X1 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  FA_X1 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  FA_X1 S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  FA_X1 S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  FA_X1 S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  FA_X1 S2_9_9 ( .A(ab_9__9_), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  FA_X1 S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), .CO(
        CARRYB_9__10_), .S(SUMB_9__10_) );
  FA_X1 S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), .CO(
        CARRYB_9__11_), .S(SUMB_9__11_) );
  FA_X1 S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), .CO(
        CARRYB_9__12_), .S(SUMB_9__12_) );
  FA_X1 S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), .CO(
        CARRYB_9__13_), .S(SUMB_9__13_) );
  FA_X1 S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), .CO(
        CARRYB_9__14_), .S(SUMB_9__14_) );
  FA_X1 S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), .CO(
        CARRYB_9__15_), .S(SUMB_9__15_) );
  FA_X1 S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), .CO(
        CARRYB_9__16_), .S(SUMB_9__16_) );
  FA_X1 S2_9_17 ( .A(ab_9__17_), .B(CARRYB_8__17_), .CI(SUMB_8__18_), .CO(
        CARRYB_9__17_), .S(SUMB_9__17_) );
  FA_X1 S2_9_18 ( .A(ab_9__18_), .B(CARRYB_8__18_), .CI(SUMB_8__19_), .CO(
        CARRYB_9__18_), .S(SUMB_9__18_) );
  FA_X1 S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), .CO(
        CARRYB_9__19_), .S(SUMB_9__19_) );
  FA_X1 S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(SUMB_8__21_), .CO(
        CARRYB_9__20_), .S(SUMB_9__20_) );
  FA_X1 S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), .CO(
        CARRYB_9__21_), .S(SUMB_9__21_) );
  FA_X1 S3_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .CI(ab_8__23_), .CO(
        CARRYB_9__22_), .S(SUMB_9__22_) );
  FA_X1 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  FA_X1 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  FA_X1 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  FA_X1 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  FA_X1 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  FA_X1 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  FA_X1 S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  FA_X1 S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  FA_X1 S2_8_8 ( .A(ab_8__8_), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  FA_X1 S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  FA_X1 S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), .CO(
        CARRYB_8__10_), .S(SUMB_8__10_) );
  FA_X1 S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), .CO(
        CARRYB_8__11_), .S(SUMB_8__11_) );
  FA_X1 S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), .CO(
        CARRYB_8__12_), .S(SUMB_8__12_) );
  FA_X1 S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), .CO(
        CARRYB_8__13_), .S(SUMB_8__13_) );
  FA_X1 S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), .CO(
        CARRYB_8__14_), .S(SUMB_8__14_) );
  FA_X1 S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), .CO(
        CARRYB_8__15_), .S(SUMB_8__15_) );
  FA_X1 S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), .CO(
        CARRYB_8__16_), .S(SUMB_8__16_) );
  FA_X1 S2_8_17 ( .A(ab_8__17_), .B(CARRYB_7__17_), .CI(SUMB_7__18_), .CO(
        CARRYB_8__17_), .S(SUMB_8__17_) );
  FA_X1 S2_8_18 ( .A(ab_8__18_), .B(CARRYB_7__18_), .CI(SUMB_7__19_), .CO(
        CARRYB_8__18_), .S(SUMB_8__18_) );
  FA_X1 S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), .CO(
        CARRYB_8__19_), .S(SUMB_8__19_) );
  FA_X1 S2_8_20 ( .A(ab_8__20_), .B(CARRYB_7__20_), .CI(SUMB_7__21_), .CO(
        CARRYB_8__20_), .S(SUMB_8__20_) );
  FA_X1 S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), .CO(
        CARRYB_8__21_), .S(SUMB_8__21_) );
  FA_X1 S3_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(ab_7__23_), .CO(
        CARRYB_8__22_), .S(SUMB_8__22_) );
  FA_X1 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(A1_5_) );
  FA_X1 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S2_7_7 ( .A(ab_7__7_), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  FA_X1 S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  FA_X1 S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  FA_X1 S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), .CO(
        CARRYB_7__10_), .S(SUMB_7__10_) );
  FA_X1 S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), .CO(
        CARRYB_7__11_), .S(SUMB_7__11_) );
  FA_X1 S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), .CO(
        CARRYB_7__12_), .S(SUMB_7__12_) );
  FA_X1 S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), .CO(
        CARRYB_7__13_), .S(SUMB_7__13_) );
  FA_X1 S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), .CO(
        CARRYB_7__14_), .S(SUMB_7__14_) );
  FA_X1 S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), .CO(
        CARRYB_7__15_), .S(SUMB_7__15_) );
  FA_X1 S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), .CO(
        CARRYB_7__16_), .S(SUMB_7__16_) );
  FA_X1 S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), .CO(
        CARRYB_7__17_), .S(SUMB_7__17_) );
  FA_X1 S2_7_18 ( .A(ab_7__18_), .B(CARRYB_6__18_), .CI(SUMB_6__19_), .CO(
        CARRYB_7__18_), .S(SUMB_7__18_) );
  FA_X1 S2_7_19 ( .A(ab_7__19_), .B(CARRYB_6__19_), .CI(SUMB_6__20_), .CO(
        CARRYB_7__19_), .S(SUMB_7__19_) );
  FA_X1 S2_7_20 ( .A(ab_7__20_), .B(CARRYB_6__20_), .CI(SUMB_6__21_), .CO(
        CARRYB_7__20_), .S(SUMB_7__20_) );
  FA_X1 S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), .CO(
        CARRYB_7__21_), .S(SUMB_7__21_) );
  FA_X1 S3_7_22 ( .A(ab_7__22_), .B(CARRYB_6__22_), .CI(ab_6__23_), .CO(
        CARRYB_7__22_), .S(SUMB_7__22_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S2_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  FA_X1 S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  FA_X1 S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  FA_X1 S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), .CO(
        CARRYB_6__10_), .S(SUMB_6__10_) );
  FA_X1 S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), .CO(
        CARRYB_6__11_), .S(SUMB_6__11_) );
  FA_X1 S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), .CO(
        CARRYB_6__12_), .S(SUMB_6__12_) );
  FA_X1 S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), .CO(
        CARRYB_6__13_), .S(SUMB_6__13_) );
  FA_X1 S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), .CO(
        CARRYB_6__14_), .S(SUMB_6__14_) );
  FA_X1 S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), .CO(
        CARRYB_6__15_), .S(SUMB_6__15_) );
  FA_X1 S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), .CO(
        CARRYB_6__16_), .S(SUMB_6__16_) );
  FA_X1 S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), .CO(
        CARRYB_6__17_), .S(SUMB_6__17_) );
  FA_X1 S2_6_18 ( .A(ab_6__18_), .B(CARRYB_5__18_), .CI(SUMB_5__19_), .CO(
        CARRYB_6__18_), .S(SUMB_6__18_) );
  FA_X1 S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), .CO(
        CARRYB_6__19_), .S(SUMB_6__19_) );
  FA_X1 S2_6_20 ( .A(ab_6__20_), .B(CARRYB_5__20_), .CI(SUMB_5__21_), .CO(
        CARRYB_6__20_), .S(SUMB_6__20_) );
  FA_X1 S2_6_21 ( .A(ab_6__21_), .B(CARRYB_5__21_), .CI(SUMB_5__22_), .CO(
        CARRYB_6__21_), .S(SUMB_6__21_) );
  FA_X1 S3_6_22 ( .A(ab_6__22_), .B(CARRYB_5__22_), .CI(ab_5__23_), .CO(
        CARRYB_6__22_), .S(SUMB_6__22_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  FA_X1 S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  FA_X1 S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  FA_X1 S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), .CO(
        CARRYB_5__10_), .S(SUMB_5__10_) );
  FA_X1 S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), .CO(
        CARRYB_5__11_), .S(SUMB_5__11_) );
  FA_X1 S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), .CO(
        CARRYB_5__12_), .S(SUMB_5__12_) );
  FA_X1 S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), .CO(
        CARRYB_5__13_), .S(SUMB_5__13_) );
  FA_X1 S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), .CO(
        CARRYB_5__14_), .S(SUMB_5__14_) );
  FA_X1 S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), .CO(
        CARRYB_5__15_), .S(SUMB_5__15_) );
  FA_X1 S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), .CO(
        CARRYB_5__16_), .S(SUMB_5__16_) );
  FA_X1 S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), .CO(
        CARRYB_5__17_), .S(SUMB_5__17_) );
  FA_X1 S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), .CO(
        CARRYB_5__18_), .S(SUMB_5__18_) );
  FA_X1 S2_5_19 ( .A(ab_5__19_), .B(CARRYB_4__19_), .CI(SUMB_4__20_), .CO(
        CARRYB_5__19_), .S(SUMB_5__19_) );
  FA_X1 S2_5_20 ( .A(ab_5__20_), .B(CARRYB_4__20_), .CI(SUMB_4__21_), .CO(
        CARRYB_5__20_), .S(SUMB_5__20_) );
  FA_X1 S2_5_21 ( .A(ab_5__21_), .B(CARRYB_4__21_), .CI(SUMB_4__22_), .CO(
        CARRYB_5__21_), .S(SUMB_5__21_) );
  FA_X1 S3_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(ab_4__23_), .CO(
        CARRYB_5__22_), .S(SUMB_5__22_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  FA_X1 S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  FA_X1 S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  FA_X1 S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), .CO(
        CARRYB_4__10_), .S(SUMB_4__10_) );
  FA_X1 S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), .CO(
        CARRYB_4__11_), .S(SUMB_4__11_) );
  FA_X1 S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), .CO(
        CARRYB_4__12_), .S(SUMB_4__12_) );
  FA_X1 S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), .CO(
        CARRYB_4__13_), .S(SUMB_4__13_) );
  FA_X1 S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), .CO(
        CARRYB_4__14_), .S(SUMB_4__14_) );
  FA_X1 S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), .CO(
        CARRYB_4__15_), .S(SUMB_4__15_) );
  FA_X1 S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), .CO(
        CARRYB_4__16_), .S(SUMB_4__16_) );
  FA_X1 S2_4_17 ( .A(ab_4__17_), .B(CARRYB_3__17_), .CI(SUMB_3__18_), .CO(
        CARRYB_4__17_), .S(SUMB_4__17_) );
  FA_X1 S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), .CO(
        CARRYB_4__18_), .S(SUMB_4__18_) );
  FA_X1 S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), .CO(
        CARRYB_4__19_), .S(SUMB_4__19_) );
  FA_X1 S2_4_20 ( .A(ab_4__20_), .B(CARRYB_3__20_), .CI(SUMB_3__21_), .CO(
        CARRYB_4__20_), .S(SUMB_4__20_) );
  FA_X1 S2_4_21 ( .A(ab_4__21_), .B(CARRYB_3__21_), .CI(SUMB_3__22_), .CO(
        CARRYB_4__21_), .S(SUMB_4__21_) );
  FA_X1 S3_4_22 ( .A(ab_4__22_), .B(CARRYB_3__22_), .CI(ab_3__23_), .CO(
        CARRYB_4__22_), .S(SUMB_4__22_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  FA_X1 S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  FA_X1 S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  FA_X1 S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), .CO(
        CARRYB_3__10_), .S(SUMB_3__10_) );
  FA_X1 S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), .CO(
        CARRYB_3__11_), .S(SUMB_3__11_) );
  FA_X1 S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), .CO(
        CARRYB_3__12_), .S(SUMB_3__12_) );
  FA_X1 S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), .CO(
        CARRYB_3__13_), .S(SUMB_3__13_) );
  FA_X1 S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), .CO(
        CARRYB_3__14_), .S(SUMB_3__14_) );
  FA_X1 S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), .CO(
        CARRYB_3__15_), .S(SUMB_3__15_) );
  FA_X1 S2_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(SUMB_2__17_), .CO(
        CARRYB_3__16_), .S(SUMB_3__16_) );
  FA_X1 S2_3_17 ( .A(ab_3__17_), .B(CARRYB_2__17_), .CI(SUMB_2__18_), .CO(
        CARRYB_3__17_), .S(SUMB_3__17_) );
  FA_X1 S2_3_18 ( .A(ab_3__18_), .B(CARRYB_2__18_), .CI(SUMB_2__19_), .CO(
        CARRYB_3__18_), .S(SUMB_3__18_) );
  FA_X1 S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), .CO(
        CARRYB_3__19_), .S(SUMB_3__19_) );
  FA_X1 S2_3_20 ( .A(ab_3__20_), .B(CARRYB_2__20_), .CI(SUMB_2__21_), .CO(
        CARRYB_3__20_), .S(SUMB_3__20_) );
  FA_X1 S2_3_21 ( .A(ab_3__21_), .B(CARRYB_2__21_), .CI(SUMB_2__22_), .CO(
        CARRYB_3__21_), .S(SUMB_3__21_) );
  FA_X1 S3_3_22 ( .A(ab_3__22_), .B(CARRYB_2__22_), .CI(ab_2__23_), .CO(
        CARRYB_3__22_), .S(SUMB_3__22_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S2_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(SUMB_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  FA_X1 S2_2_7 ( .A(ab_2__7_), .B(CARRYB_1__7_), .CI(SUMB_1__8_), .CO(
        CARRYB_2__7_), .S(SUMB_2__7_) );
  FA_X1 S2_2_8 ( .A(ab_2__8_), .B(CARRYB_1__8_), .CI(SUMB_1__9_), .CO(
        CARRYB_2__8_), .S(SUMB_2__8_) );
  FA_X1 S2_2_9 ( .A(ab_2__9_), .B(CARRYB_1__9_), .CI(SUMB_1__10_), .CO(
        CARRYB_2__9_), .S(SUMB_2__9_) );
  FA_X1 S2_2_10 ( .A(ab_2__10_), .B(CARRYB_1__10_), .CI(SUMB_1__11_), .CO(
        CARRYB_2__10_), .S(SUMB_2__10_) );
  FA_X1 S2_2_11 ( .A(ab_2__11_), .B(CARRYB_1__11_), .CI(SUMB_1__12_), .CO(
        CARRYB_2__11_), .S(SUMB_2__11_) );
  FA_X1 S2_2_12 ( .A(ab_2__12_), .B(CARRYB_1__12_), .CI(SUMB_1__13_), .CO(
        CARRYB_2__12_), .S(SUMB_2__12_) );
  FA_X1 S2_2_13 ( .A(ab_2__13_), .B(CARRYB_1__13_), .CI(SUMB_1__14_), .CO(
        CARRYB_2__13_), .S(SUMB_2__13_) );
  FA_X1 S2_2_14 ( .A(ab_2__14_), .B(CARRYB_1__14_), .CI(SUMB_1__15_), .CO(
        CARRYB_2__14_), .S(SUMB_2__14_) );
  FA_X1 S2_2_15 ( .A(ab_2__15_), .B(CARRYB_1__15_), .CI(SUMB_1__16_), .CO(
        CARRYB_2__15_), .S(SUMB_2__15_) );
  FA_X1 S2_2_16 ( .A(ab_2__16_), .B(CARRYB_1__16_), .CI(SUMB_1__17_), .CO(
        CARRYB_2__16_), .S(SUMB_2__16_) );
  FA_X1 S2_2_17 ( .A(ab_2__17_), .B(CARRYB_1__17_), .CI(SUMB_1__18_), .CO(
        CARRYB_2__17_), .S(SUMB_2__17_) );
  FA_X1 S2_2_18 ( .A(ab_2__18_), .B(CARRYB_1__18_), .CI(SUMB_1__19_), .CO(
        CARRYB_2__18_), .S(SUMB_2__18_) );
  FA_X1 S2_2_19 ( .A(ab_2__19_), .B(CARRYB_1__19_), .CI(SUMB_1__20_), .CO(
        CARRYB_2__19_), .S(SUMB_2__19_) );
  FA_X1 S2_2_20 ( .A(ab_2__20_), .B(CARRYB_1__20_), .CI(SUMB_1__21_), .CO(
        CARRYB_2__20_), .S(SUMB_2__20_) );
  FA_X1 S2_2_21 ( .A(ab_2__21_), .B(CARRYB_1__21_), .CI(SUMB_1__22_), .CO(
        CARRYB_2__21_), .S(SUMB_2__21_) );
  FA_X1 S3_2_22 ( .A(ab_2__22_), .B(CARRYB_1__22_), .CI(ab_1__23_), .CO(
        CARRYB_2__22_), .S(SUMB_2__22_) );
  iir_filter_DW01_add_9 FS_1 ( .A({A1_45_, A1_44_, A1_43_, A1_42_, A1_41_, 
        A1_40_, A1_39_, A1_38_, A1_37_, A1_36_, A1_35_, A1_34_, A1_33_, A1_32_, 
        A1_31_, A1_30_, A1_29_, A1_28_, A1_27_, A1_26_, A1_25_, A1_24_, A1_23_, 
        A1_22_, A1_21_, A1_20_, A1_19_, A1_18_, A1_17_, A1_16_, A1_15_, A1_14_, 
        A1_13_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, A1_5_, 
        A1_4_, A1_3_, A1_2_, A1_1_, A1_0_}), .B({A2_45_, A2_44_, A2_43_, 
        A2_42_, A2_41_, A2_40_, A2_39_, A2_38_, A2_37_, A2_36_, A2_35_, A2_34_, 
        A2_33_, A2_32_, A2_31_, A2_30_, A2_29_, A2_28_, A2_27_, A2_26_, A2_25_, 
        A2_24_, A2_23_, A2_22_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({PRODUCT[47], SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, PRODUCT[44:22], SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21}) );
  BUF_X1 U2 ( .A(QB), .Z(n1) );
  BUF_X1 U3 ( .A(QB), .Z(n2) );
  BUF_X1 U4 ( .A(QA), .Z(n3) );
  BUF_X1 U5 ( .A(QA), .Z(n4) );
  INV_X1 U6 ( .A(B[22]), .ZN(n15) );
  INV_X1 U7 ( .A(B[21]), .ZN(n16) );
  INV_X1 U8 ( .A(B[20]), .ZN(n17) );
  INV_X1 U9 ( .A(B[19]), .ZN(n19) );
  INV_X1 U10 ( .A(B[18]), .ZN(n20) );
  INV_X1 U11 ( .A(B[17]), .ZN(n21) );
  INV_X1 U12 ( .A(B[16]), .ZN(n22) );
  INV_X1 U13 ( .A(B[15]), .ZN(n23) );
  INV_X1 U14 ( .A(B[14]), .ZN(n24) );
  INV_X1 U15 ( .A(B[13]), .ZN(n25) );
  INV_X1 U16 ( .A(B[12]), .ZN(n26) );
  INV_X1 U17 ( .A(B[11]), .ZN(n27) );
  INV_X1 U18 ( .A(B[10]), .ZN(n28) );
  INV_X1 U19 ( .A(B[9]), .ZN(n7) );
  INV_X1 U20 ( .A(B[8]), .ZN(n8) );
  INV_X1 U21 ( .A(B[7]), .ZN(n9) );
  INV_X1 U22 ( .A(B[6]), .ZN(n10) );
  INV_X1 U23 ( .A(B[5]), .ZN(n11) );
  INV_X1 U24 ( .A(B[4]), .ZN(n12) );
  INV_X1 U25 ( .A(B[3]), .ZN(n13) );
  INV_X1 U26 ( .A(B[2]), .ZN(n14) );
  INV_X1 U27 ( .A(A[2]), .ZN(n36) );
  INV_X1 U28 ( .A(A[3]), .ZN(n35) );
  INV_X1 U29 ( .A(A[4]), .ZN(n34) );
  INV_X1 U30 ( .A(A[5]), .ZN(n33) );
  INV_X1 U31 ( .A(A[6]), .ZN(n32) );
  INV_X1 U32 ( .A(B[1]), .ZN(n18) );
  INV_X1 U33 ( .A(A[1]), .ZN(n40) );
  INV_X1 U34 ( .A(B[0]), .ZN(n29) );
  INV_X1 U35 ( .A(A[0]), .ZN(n51) );
  INV_X1 U36 ( .A(A[7]), .ZN(n31) );
  INV_X1 U37 ( .A(A[8]), .ZN(n30) );
  INV_X1 U38 ( .A(A[10]), .ZN(n50) );
  INV_X1 U39 ( .A(A[11]), .ZN(n49) );
  INV_X1 U40 ( .A(A[12]), .ZN(n48) );
  INV_X1 U41 ( .A(A[13]), .ZN(n47) );
  INV_X1 U42 ( .A(A[14]), .ZN(n46) );
  INV_X1 U43 ( .A(A[9]), .ZN(n6) );
  INV_X1 U44 ( .A(A[22]), .ZN(n37) );
  INV_X1 U45 ( .A(A[15]), .ZN(n45) );
  INV_X1 U46 ( .A(A[16]), .ZN(n44) );
  INV_X1 U47 ( .A(A[17]), .ZN(n43) );
  INV_X1 U48 ( .A(A[18]), .ZN(n42) );
  INV_X1 U49 ( .A(A[19]), .ZN(n41) );
  INV_X1 U50 ( .A(A[20]), .ZN(n39) );
  INV_X1 U51 ( .A(A[21]), .ZN(n38) );
  AND2_X1 U52 ( .A1(SUMB_23__23_), .A2(CARRYB_23__22_), .ZN(A2_45_) );
  XOR2_X1 U53 ( .A(CARRYB_23__22_), .B(SUMB_23__23_), .Z(A1_44_) );
  AND2_X1 U54 ( .A1(SUMB_23__22_), .A2(CARRYB_23__21_), .ZN(A2_44_) );
  XOR2_X1 U55 ( .A(CARRYB_23__21_), .B(SUMB_23__22_), .Z(A1_43_) );
  AND2_X1 U56 ( .A1(SUMB_23__21_), .A2(CARRYB_23__20_), .ZN(A2_43_) );
  XOR2_X1 U57 ( .A(CARRYB_23__20_), .B(SUMB_23__21_), .Z(A1_42_) );
  AND2_X1 U58 ( .A1(SUMB_23__20_), .A2(CARRYB_23__19_), .ZN(A2_42_) );
  XOR2_X1 U59 ( .A(CARRYB_23__19_), .B(SUMB_23__20_), .Z(A1_41_) );
  AND2_X1 U60 ( .A1(SUMB_23__19_), .A2(CARRYB_23__18_), .ZN(A2_41_) );
  XOR2_X1 U61 ( .A(CARRYB_23__18_), .B(SUMB_23__19_), .Z(A1_40_) );
  AND2_X1 U62 ( .A1(SUMB_23__18_), .A2(CARRYB_23__17_), .ZN(A2_40_) );
  XOR2_X1 U63 ( .A(CARRYB_23__17_), .B(SUMB_23__18_), .Z(A1_39_) );
  AND2_X1 U64 ( .A1(SUMB_23__17_), .A2(CARRYB_23__16_), .ZN(A2_39_) );
  XOR2_X1 U65 ( .A(CARRYB_23__16_), .B(SUMB_23__17_), .Z(A1_38_) );
  AND2_X1 U66 ( .A1(SUMB_23__16_), .A2(CARRYB_23__15_), .ZN(A2_38_) );
  XOR2_X1 U67 ( .A(CARRYB_23__15_), .B(SUMB_23__16_), .Z(A1_37_) );
  AND2_X1 U68 ( .A1(SUMB_23__15_), .A2(CARRYB_23__14_), .ZN(A2_37_) );
  XOR2_X1 U69 ( .A(CARRYB_23__14_), .B(SUMB_23__15_), .Z(A1_36_) );
  AND2_X1 U70 ( .A1(SUMB_23__14_), .A2(CARRYB_23__13_), .ZN(A2_36_) );
  XOR2_X1 U71 ( .A(CARRYB_23__13_), .B(SUMB_23__14_), .Z(A1_35_) );
  AND2_X1 U72 ( .A1(SUMB_23__13_), .A2(CARRYB_23__12_), .ZN(A2_35_) );
  XOR2_X1 U73 ( .A(CARRYB_23__12_), .B(SUMB_23__13_), .Z(A1_34_) );
  AND2_X1 U74 ( .A1(SUMB_23__12_), .A2(CARRYB_23__11_), .ZN(A2_34_) );
  XOR2_X1 U75 ( .A(CARRYB_23__11_), .B(SUMB_23__12_), .Z(A1_33_) );
  AND2_X1 U76 ( .A1(SUMB_23__11_), .A2(CARRYB_23__10_), .ZN(A2_33_) );
  XOR2_X1 U77 ( .A(CARRYB_23__10_), .B(SUMB_23__11_), .Z(A1_32_) );
  AND2_X1 U78 ( .A1(SUMB_23__10_), .A2(CARRYB_23__9_), .ZN(A2_32_) );
  XOR2_X1 U79 ( .A(CARRYB_23__9_), .B(SUMB_23__10_), .Z(A1_31_) );
  AND2_X1 U80 ( .A1(SUMB_23__9_), .A2(CARRYB_23__8_), .ZN(A2_31_) );
  XOR2_X1 U81 ( .A(CARRYB_23__8_), .B(SUMB_23__9_), .Z(A1_30_) );
  AND2_X1 U82 ( .A1(SUMB_23__8_), .A2(CARRYB_23__7_), .ZN(A2_30_) );
  XOR2_X1 U83 ( .A(CARRYB_23__7_), .B(SUMB_23__8_), .Z(A1_29_) );
  AND2_X1 U84 ( .A1(SUMB_23__7_), .A2(CARRYB_23__6_), .ZN(A2_29_) );
  XOR2_X1 U85 ( .A(CARRYB_23__6_), .B(SUMB_23__7_), .Z(A1_28_) );
  AND2_X1 U86 ( .A1(SUMB_23__6_), .A2(CARRYB_23__5_), .ZN(A2_28_) );
  XOR2_X1 U87 ( .A(CARRYB_23__5_), .B(SUMB_23__6_), .Z(A1_27_) );
  AND2_X1 U88 ( .A1(SUMB_23__5_), .A2(CARRYB_23__4_), .ZN(A2_27_) );
  XOR2_X1 U89 ( .A(CARRYB_23__4_), .B(SUMB_23__5_), .Z(A1_26_) );
  AND2_X1 U90 ( .A1(SUMB_23__4_), .A2(CARRYB_23__3_), .ZN(A2_26_) );
  XOR2_X1 U91 ( .A(CARRYB_23__3_), .B(SUMB_23__4_), .Z(A1_25_) );
  AND2_X1 U92 ( .A1(SUMB_23__3_), .A2(CARRYB_23__2_), .ZN(A2_25_) );
  XOR2_X1 U93 ( .A(CARRYB_23__2_), .B(SUMB_23__3_), .Z(A1_24_) );
  AND2_X1 U94 ( .A1(SUMB_23__2_), .A2(CARRYB_23__1_), .ZN(A2_24_) );
  XOR2_X1 U95 ( .A(CARRYB_23__1_), .B(SUMB_23__2_), .Z(A1_23_) );
  AND2_X1 U96 ( .A1(SUMB_23__1_), .A2(CARRYB_23__0_), .ZN(A2_23_) );
  XOR2_X1 U97 ( .A(CARRYB_23__0_), .B(SUMB_23__1_), .Z(A1_22_) );
  AND2_X1 U98 ( .A1(ab_1__22_), .A2(ab_0__23_), .ZN(CARRYB_1__22_) );
  XOR2_X1 U99 ( .A(ab_1__22_), .B(ab_0__23_), .Z(SUMB_1__22_) );
  AND2_X1 U100 ( .A1(ab_1__21_), .A2(ab_0__22_), .ZN(CARRYB_1__21_) );
  XOR2_X1 U101 ( .A(ab_1__21_), .B(ab_0__22_), .Z(SUMB_1__21_) );
  AND2_X1 U102 ( .A1(ab_1__20_), .A2(ab_0__21_), .ZN(CARRYB_1__20_) );
  XOR2_X1 U103 ( .A(ab_1__20_), .B(ab_0__21_), .Z(SUMB_1__20_) );
  AND2_X1 U104 ( .A1(ab_1__19_), .A2(ab_0__20_), .ZN(CARRYB_1__19_) );
  XOR2_X1 U105 ( .A(ab_1__19_), .B(ab_0__20_), .Z(SUMB_1__19_) );
  AND2_X1 U106 ( .A1(ab_1__18_), .A2(ab_0__19_), .ZN(CARRYB_1__18_) );
  XOR2_X1 U107 ( .A(ab_1__18_), .B(ab_0__19_), .Z(SUMB_1__18_) );
  AND2_X1 U108 ( .A1(ab_1__17_), .A2(ab_0__18_), .ZN(CARRYB_1__17_) );
  XOR2_X1 U109 ( .A(ab_1__17_), .B(ab_0__18_), .Z(SUMB_1__17_) );
  AND2_X1 U110 ( .A1(ab_1__16_), .A2(ab_0__17_), .ZN(CARRYB_1__16_) );
  XOR2_X1 U111 ( .A(ab_1__16_), .B(ab_0__17_), .Z(SUMB_1__16_) );
  AND2_X1 U112 ( .A1(ab_1__15_), .A2(ab_0__16_), .ZN(CARRYB_1__15_) );
  XOR2_X1 U113 ( .A(ab_1__15_), .B(ab_0__16_), .Z(SUMB_1__15_) );
  AND2_X1 U114 ( .A1(ab_1__14_), .A2(ab_0__15_), .ZN(CARRYB_1__14_) );
  XOR2_X1 U115 ( .A(ab_1__14_), .B(ab_0__15_), .Z(SUMB_1__14_) );
  AND2_X1 U116 ( .A1(ab_1__13_), .A2(ab_0__14_), .ZN(CARRYB_1__13_) );
  XOR2_X1 U117 ( .A(ab_1__13_), .B(ab_0__14_), .Z(SUMB_1__13_) );
  AND2_X1 U118 ( .A1(ab_1__12_), .A2(ab_0__13_), .ZN(CARRYB_1__12_) );
  XOR2_X1 U119 ( .A(ab_1__12_), .B(ab_0__13_), .Z(SUMB_1__12_) );
  AND2_X1 U120 ( .A1(ab_1__11_), .A2(ab_0__12_), .ZN(CARRYB_1__11_) );
  XOR2_X1 U121 ( .A(ab_1__11_), .B(ab_0__12_), .Z(SUMB_1__11_) );
  AND2_X1 U122 ( .A1(ab_1__10_), .A2(ab_0__11_), .ZN(CARRYB_1__10_) );
  XOR2_X1 U123 ( .A(ab_1__10_), .B(ab_0__11_), .Z(SUMB_1__10_) );
  AND2_X1 U124 ( .A1(ab_1__9_), .A2(ab_0__10_), .ZN(CARRYB_1__9_) );
  XOR2_X1 U125 ( .A(ab_1__9_), .B(ab_0__10_), .Z(SUMB_1__9_) );
  AND2_X1 U126 ( .A1(ab_1__8_), .A2(ab_0__9_), .ZN(CARRYB_1__8_) );
  XOR2_X1 U127 ( .A(ab_1__8_), .B(ab_0__9_), .Z(SUMB_1__8_) );
  AND2_X1 U128 ( .A1(ab_1__7_), .A2(ab_0__8_), .ZN(CARRYB_1__7_) );
  XOR2_X1 U129 ( .A(ab_1__7_), .B(ab_0__8_), .Z(SUMB_1__7_) );
  AND2_X1 U130 ( .A1(ab_1__6_), .A2(ab_0__7_), .ZN(CARRYB_1__6_) );
  XOR2_X1 U131 ( .A(ab_1__6_), .B(ab_0__7_), .Z(SUMB_1__6_) );
  AND2_X1 U132 ( .A1(ab_1__5_), .A2(ab_0__6_), .ZN(CARRYB_1__5_) );
  XOR2_X1 U133 ( .A(ab_1__5_), .B(ab_0__6_), .Z(SUMB_1__5_) );
  AND2_X1 U134 ( .A1(ab_1__4_), .A2(ab_0__5_), .ZN(CARRYB_1__4_) );
  XOR2_X1 U135 ( .A(ab_1__4_), .B(ab_0__5_), .Z(SUMB_1__4_) );
  AND2_X1 U136 ( .A1(ab_1__3_), .A2(ab_0__4_), .ZN(CARRYB_1__3_) );
  XOR2_X1 U137 ( .A(ab_1__3_), .B(ab_0__4_), .Z(SUMB_1__3_) );
  AND2_X1 U138 ( .A1(ab_1__2_), .A2(ab_0__3_), .ZN(CARRYB_1__2_) );
  XOR2_X1 U139 ( .A(ab_1__2_), .B(ab_0__3_), .Z(SUMB_1__2_) );
  AND2_X1 U140 ( .A1(ab_1__1_), .A2(ab_0__2_), .ZN(CARRYB_1__1_) );
  XOR2_X1 U141 ( .A(ab_1__1_), .B(ab_0__2_), .Z(SUMB_1__1_) );
  NOR2_X1 U142 ( .A1(n6), .A2(n7), .ZN(ab_9__9_) );
  NOR2_X1 U143 ( .A1(n6), .A2(n8), .ZN(ab_9__8_) );
  NOR2_X1 U144 ( .A1(n6), .A2(n9), .ZN(ab_9__7_) );
  NOR2_X1 U145 ( .A1(n6), .A2(n10), .ZN(ab_9__6_) );
  NOR2_X1 U146 ( .A1(n6), .A2(n11), .ZN(ab_9__5_) );
  NOR2_X1 U147 ( .A1(n6), .A2(n12), .ZN(ab_9__4_) );
  NOR2_X1 U148 ( .A1(n6), .A2(n13), .ZN(ab_9__3_) );
  NOR2_X1 U149 ( .A1(n6), .A2(n14), .ZN(ab_9__2_) );
  NOR2_X1 U150 ( .A1(A[9]), .A2(n1), .ZN(ab_9__23_) );
  NOR2_X1 U151 ( .A1(n6), .A2(n15), .ZN(ab_9__22_) );
  NOR2_X1 U152 ( .A1(n6), .A2(n16), .ZN(ab_9__21_) );
  NOR2_X1 U153 ( .A1(n6), .A2(n17), .ZN(ab_9__20_) );
  NOR2_X1 U154 ( .A1(n6), .A2(n18), .ZN(ab_9__1_) );
  NOR2_X1 U155 ( .A1(n6), .A2(n19), .ZN(ab_9__19_) );
  NOR2_X1 U156 ( .A1(n6), .A2(n20), .ZN(ab_9__18_) );
  NOR2_X1 U157 ( .A1(n6), .A2(n21), .ZN(ab_9__17_) );
  NOR2_X1 U158 ( .A1(n6), .A2(n22), .ZN(ab_9__16_) );
  NOR2_X1 U159 ( .A1(n6), .A2(n23), .ZN(ab_9__15_) );
  NOR2_X1 U160 ( .A1(n6), .A2(n24), .ZN(ab_9__14_) );
  NOR2_X1 U161 ( .A1(n6), .A2(n25), .ZN(ab_9__13_) );
  NOR2_X1 U162 ( .A1(n6), .A2(n26), .ZN(ab_9__12_) );
  NOR2_X1 U163 ( .A1(n6), .A2(n27), .ZN(ab_9__11_) );
  NOR2_X1 U164 ( .A1(n6), .A2(n28), .ZN(ab_9__10_) );
  NOR2_X1 U165 ( .A1(n6), .A2(n29), .ZN(ab_9__0_) );
  NOR2_X1 U166 ( .A1(n7), .A2(n30), .ZN(ab_8__9_) );
  NOR2_X1 U167 ( .A1(n8), .A2(n30), .ZN(ab_8__8_) );
  NOR2_X1 U168 ( .A1(n9), .A2(n30), .ZN(ab_8__7_) );
  NOR2_X1 U169 ( .A1(n10), .A2(n30), .ZN(ab_8__6_) );
  NOR2_X1 U170 ( .A1(n11), .A2(n30), .ZN(ab_8__5_) );
  NOR2_X1 U171 ( .A1(n12), .A2(n30), .ZN(ab_8__4_) );
  NOR2_X1 U172 ( .A1(n13), .A2(n30), .ZN(ab_8__3_) );
  NOR2_X1 U173 ( .A1(n14), .A2(n30), .ZN(ab_8__2_) );
  NOR2_X1 U174 ( .A1(A[8]), .A2(n1), .ZN(ab_8__23_) );
  NOR2_X1 U175 ( .A1(n15), .A2(n30), .ZN(ab_8__22_) );
  NOR2_X1 U176 ( .A1(n16), .A2(n30), .ZN(ab_8__21_) );
  NOR2_X1 U177 ( .A1(n17), .A2(n30), .ZN(ab_8__20_) );
  NOR2_X1 U178 ( .A1(n18), .A2(n30), .ZN(ab_8__1_) );
  NOR2_X1 U179 ( .A1(n19), .A2(n30), .ZN(ab_8__19_) );
  NOR2_X1 U180 ( .A1(n20), .A2(n30), .ZN(ab_8__18_) );
  NOR2_X1 U181 ( .A1(n21), .A2(n30), .ZN(ab_8__17_) );
  NOR2_X1 U182 ( .A1(n22), .A2(n30), .ZN(ab_8__16_) );
  NOR2_X1 U183 ( .A1(n23), .A2(n30), .ZN(ab_8__15_) );
  NOR2_X1 U184 ( .A1(n24), .A2(n30), .ZN(ab_8__14_) );
  NOR2_X1 U185 ( .A1(n25), .A2(n30), .ZN(ab_8__13_) );
  NOR2_X1 U186 ( .A1(n26), .A2(n30), .ZN(ab_8__12_) );
  NOR2_X1 U187 ( .A1(n27), .A2(n30), .ZN(ab_8__11_) );
  NOR2_X1 U188 ( .A1(n28), .A2(n30), .ZN(ab_8__10_) );
  NOR2_X1 U189 ( .A1(n29), .A2(n30), .ZN(ab_8__0_) );
  NOR2_X1 U190 ( .A1(n7), .A2(n31), .ZN(ab_7__9_) );
  NOR2_X1 U191 ( .A1(n8), .A2(n31), .ZN(ab_7__8_) );
  NOR2_X1 U192 ( .A1(n9), .A2(n31), .ZN(ab_7__7_) );
  NOR2_X1 U193 ( .A1(n10), .A2(n31), .ZN(ab_7__6_) );
  NOR2_X1 U194 ( .A1(n11), .A2(n31), .ZN(ab_7__5_) );
  NOR2_X1 U195 ( .A1(n12), .A2(n31), .ZN(ab_7__4_) );
  NOR2_X1 U196 ( .A1(n13), .A2(n31), .ZN(ab_7__3_) );
  NOR2_X1 U197 ( .A1(n14), .A2(n31), .ZN(ab_7__2_) );
  NOR2_X1 U198 ( .A1(A[7]), .A2(n1), .ZN(ab_7__23_) );
  NOR2_X1 U199 ( .A1(n15), .A2(n31), .ZN(ab_7__22_) );
  NOR2_X1 U200 ( .A1(n16), .A2(n31), .ZN(ab_7__21_) );
  NOR2_X1 U201 ( .A1(n17), .A2(n31), .ZN(ab_7__20_) );
  NOR2_X1 U202 ( .A1(n18), .A2(n31), .ZN(ab_7__1_) );
  NOR2_X1 U203 ( .A1(n19), .A2(n31), .ZN(ab_7__19_) );
  NOR2_X1 U204 ( .A1(n20), .A2(n31), .ZN(ab_7__18_) );
  NOR2_X1 U205 ( .A1(n21), .A2(n31), .ZN(ab_7__17_) );
  NOR2_X1 U206 ( .A1(n22), .A2(n31), .ZN(ab_7__16_) );
  NOR2_X1 U207 ( .A1(n23), .A2(n31), .ZN(ab_7__15_) );
  NOR2_X1 U208 ( .A1(n24), .A2(n31), .ZN(ab_7__14_) );
  NOR2_X1 U209 ( .A1(n25), .A2(n31), .ZN(ab_7__13_) );
  NOR2_X1 U210 ( .A1(n26), .A2(n31), .ZN(ab_7__12_) );
  NOR2_X1 U211 ( .A1(n27), .A2(n31), .ZN(ab_7__11_) );
  NOR2_X1 U212 ( .A1(n28), .A2(n31), .ZN(ab_7__10_) );
  NOR2_X1 U213 ( .A1(n29), .A2(n31), .ZN(ab_7__0_) );
  NOR2_X1 U214 ( .A1(n7), .A2(n32), .ZN(ab_6__9_) );
  NOR2_X1 U215 ( .A1(n8), .A2(n32), .ZN(ab_6__8_) );
  NOR2_X1 U216 ( .A1(n9), .A2(n32), .ZN(ab_6__7_) );
  NOR2_X1 U217 ( .A1(n10), .A2(n32), .ZN(ab_6__6_) );
  NOR2_X1 U218 ( .A1(n11), .A2(n32), .ZN(ab_6__5_) );
  NOR2_X1 U219 ( .A1(n12), .A2(n32), .ZN(ab_6__4_) );
  NOR2_X1 U220 ( .A1(n13), .A2(n32), .ZN(ab_6__3_) );
  NOR2_X1 U221 ( .A1(n14), .A2(n32), .ZN(ab_6__2_) );
  NOR2_X1 U222 ( .A1(A[6]), .A2(n1), .ZN(ab_6__23_) );
  NOR2_X1 U223 ( .A1(n15), .A2(n32), .ZN(ab_6__22_) );
  NOR2_X1 U224 ( .A1(n16), .A2(n32), .ZN(ab_6__21_) );
  NOR2_X1 U225 ( .A1(n17), .A2(n32), .ZN(ab_6__20_) );
  NOR2_X1 U226 ( .A1(n18), .A2(n32), .ZN(ab_6__1_) );
  NOR2_X1 U227 ( .A1(n19), .A2(n32), .ZN(ab_6__19_) );
  NOR2_X1 U228 ( .A1(n20), .A2(n32), .ZN(ab_6__18_) );
  NOR2_X1 U229 ( .A1(n21), .A2(n32), .ZN(ab_6__17_) );
  NOR2_X1 U230 ( .A1(n22), .A2(n32), .ZN(ab_6__16_) );
  NOR2_X1 U231 ( .A1(n23), .A2(n32), .ZN(ab_6__15_) );
  NOR2_X1 U232 ( .A1(n24), .A2(n32), .ZN(ab_6__14_) );
  NOR2_X1 U233 ( .A1(n25), .A2(n32), .ZN(ab_6__13_) );
  NOR2_X1 U234 ( .A1(n26), .A2(n32), .ZN(ab_6__12_) );
  NOR2_X1 U235 ( .A1(n27), .A2(n32), .ZN(ab_6__11_) );
  NOR2_X1 U236 ( .A1(n28), .A2(n32), .ZN(ab_6__10_) );
  NOR2_X1 U237 ( .A1(n29), .A2(n32), .ZN(ab_6__0_) );
  NOR2_X1 U238 ( .A1(n7), .A2(n33), .ZN(ab_5__9_) );
  NOR2_X1 U239 ( .A1(n8), .A2(n33), .ZN(ab_5__8_) );
  NOR2_X1 U240 ( .A1(n9), .A2(n33), .ZN(ab_5__7_) );
  NOR2_X1 U241 ( .A1(n10), .A2(n33), .ZN(ab_5__6_) );
  NOR2_X1 U242 ( .A1(n11), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U243 ( .A1(n12), .A2(n33), .ZN(ab_5__4_) );
  NOR2_X1 U244 ( .A1(n13), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U245 ( .A1(n14), .A2(n33), .ZN(ab_5__2_) );
  NOR2_X1 U246 ( .A1(A[5]), .A2(n1), .ZN(ab_5__23_) );
  NOR2_X1 U247 ( .A1(n15), .A2(n33), .ZN(ab_5__22_) );
  NOR2_X1 U248 ( .A1(n16), .A2(n33), .ZN(ab_5__21_) );
  NOR2_X1 U249 ( .A1(n17), .A2(n33), .ZN(ab_5__20_) );
  NOR2_X1 U250 ( .A1(n18), .A2(n33), .ZN(ab_5__1_) );
  NOR2_X1 U251 ( .A1(n19), .A2(n33), .ZN(ab_5__19_) );
  NOR2_X1 U252 ( .A1(n20), .A2(n33), .ZN(ab_5__18_) );
  NOR2_X1 U253 ( .A1(n21), .A2(n33), .ZN(ab_5__17_) );
  NOR2_X1 U254 ( .A1(n22), .A2(n33), .ZN(ab_5__16_) );
  NOR2_X1 U255 ( .A1(n23), .A2(n33), .ZN(ab_5__15_) );
  NOR2_X1 U256 ( .A1(n24), .A2(n33), .ZN(ab_5__14_) );
  NOR2_X1 U257 ( .A1(n25), .A2(n33), .ZN(ab_5__13_) );
  NOR2_X1 U258 ( .A1(n26), .A2(n33), .ZN(ab_5__12_) );
  NOR2_X1 U259 ( .A1(n27), .A2(n33), .ZN(ab_5__11_) );
  NOR2_X1 U260 ( .A1(n28), .A2(n33), .ZN(ab_5__10_) );
  NOR2_X1 U261 ( .A1(n29), .A2(n33), .ZN(ab_5__0_) );
  NOR2_X1 U262 ( .A1(n7), .A2(n34), .ZN(ab_4__9_) );
  NOR2_X1 U263 ( .A1(n8), .A2(n34), .ZN(ab_4__8_) );
  NOR2_X1 U264 ( .A1(n9), .A2(n34), .ZN(ab_4__7_) );
  NOR2_X1 U265 ( .A1(n10), .A2(n34), .ZN(ab_4__6_) );
  NOR2_X1 U266 ( .A1(n11), .A2(n34), .ZN(ab_4__5_) );
  NOR2_X1 U267 ( .A1(n12), .A2(n34), .ZN(ab_4__4_) );
  NOR2_X1 U268 ( .A1(n13), .A2(n34), .ZN(ab_4__3_) );
  NOR2_X1 U269 ( .A1(n14), .A2(n34), .ZN(ab_4__2_) );
  NOR2_X1 U270 ( .A1(A[4]), .A2(n1), .ZN(ab_4__23_) );
  NOR2_X1 U271 ( .A1(n15), .A2(n34), .ZN(ab_4__22_) );
  NOR2_X1 U272 ( .A1(n16), .A2(n34), .ZN(ab_4__21_) );
  NOR2_X1 U273 ( .A1(n17), .A2(n34), .ZN(ab_4__20_) );
  NOR2_X1 U274 ( .A1(n18), .A2(n34), .ZN(ab_4__1_) );
  NOR2_X1 U275 ( .A1(n19), .A2(n34), .ZN(ab_4__19_) );
  NOR2_X1 U276 ( .A1(n20), .A2(n34), .ZN(ab_4__18_) );
  NOR2_X1 U277 ( .A1(n21), .A2(n34), .ZN(ab_4__17_) );
  NOR2_X1 U278 ( .A1(n22), .A2(n34), .ZN(ab_4__16_) );
  NOR2_X1 U279 ( .A1(n23), .A2(n34), .ZN(ab_4__15_) );
  NOR2_X1 U280 ( .A1(n24), .A2(n34), .ZN(ab_4__14_) );
  NOR2_X1 U281 ( .A1(n25), .A2(n34), .ZN(ab_4__13_) );
  NOR2_X1 U282 ( .A1(n26), .A2(n34), .ZN(ab_4__12_) );
  NOR2_X1 U283 ( .A1(n27), .A2(n34), .ZN(ab_4__11_) );
  NOR2_X1 U284 ( .A1(n28), .A2(n34), .ZN(ab_4__10_) );
  NOR2_X1 U285 ( .A1(n29), .A2(n34), .ZN(ab_4__0_) );
  NOR2_X1 U286 ( .A1(n7), .A2(n35), .ZN(ab_3__9_) );
  NOR2_X1 U287 ( .A1(n8), .A2(n35), .ZN(ab_3__8_) );
  NOR2_X1 U288 ( .A1(n9), .A2(n35), .ZN(ab_3__7_) );
  NOR2_X1 U289 ( .A1(n10), .A2(n35), .ZN(ab_3__6_) );
  NOR2_X1 U290 ( .A1(n11), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U291 ( .A1(n12), .A2(n35), .ZN(ab_3__4_) );
  NOR2_X1 U292 ( .A1(n13), .A2(n35), .ZN(ab_3__3_) );
  NOR2_X1 U293 ( .A1(n14), .A2(n35), .ZN(ab_3__2_) );
  NOR2_X1 U294 ( .A1(A[3]), .A2(n1), .ZN(ab_3__23_) );
  NOR2_X1 U295 ( .A1(n15), .A2(n35), .ZN(ab_3__22_) );
  NOR2_X1 U296 ( .A1(n16), .A2(n35), .ZN(ab_3__21_) );
  NOR2_X1 U297 ( .A1(n17), .A2(n35), .ZN(ab_3__20_) );
  NOR2_X1 U298 ( .A1(n18), .A2(n35), .ZN(ab_3__1_) );
  NOR2_X1 U299 ( .A1(n19), .A2(n35), .ZN(ab_3__19_) );
  NOR2_X1 U300 ( .A1(n20), .A2(n35), .ZN(ab_3__18_) );
  NOR2_X1 U301 ( .A1(n21), .A2(n35), .ZN(ab_3__17_) );
  NOR2_X1 U302 ( .A1(n22), .A2(n35), .ZN(ab_3__16_) );
  NOR2_X1 U303 ( .A1(n23), .A2(n35), .ZN(ab_3__15_) );
  NOR2_X1 U304 ( .A1(n24), .A2(n35), .ZN(ab_3__14_) );
  NOR2_X1 U305 ( .A1(n25), .A2(n35), .ZN(ab_3__13_) );
  NOR2_X1 U306 ( .A1(n26), .A2(n35), .ZN(ab_3__12_) );
  NOR2_X1 U307 ( .A1(n27), .A2(n35), .ZN(ab_3__11_) );
  NOR2_X1 U308 ( .A1(n28), .A2(n35), .ZN(ab_3__10_) );
  NOR2_X1 U309 ( .A1(n29), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U310 ( .A1(n7), .A2(n36), .ZN(ab_2__9_) );
  NOR2_X1 U311 ( .A1(n8), .A2(n36), .ZN(ab_2__8_) );
  NOR2_X1 U312 ( .A1(n9), .A2(n36), .ZN(ab_2__7_) );
  NOR2_X1 U313 ( .A1(n10), .A2(n36), .ZN(ab_2__6_) );
  NOR2_X1 U314 ( .A1(n11), .A2(n36), .ZN(ab_2__5_) );
  NOR2_X1 U315 ( .A1(n12), .A2(n36), .ZN(ab_2__4_) );
  NOR2_X1 U316 ( .A1(n13), .A2(n36), .ZN(ab_2__3_) );
  NOR2_X1 U317 ( .A1(n14), .A2(n36), .ZN(ab_2__2_) );
  NOR2_X1 U318 ( .A1(A[2]), .A2(n1), .ZN(ab_2__23_) );
  NOR2_X1 U319 ( .A1(n15), .A2(n36), .ZN(ab_2__22_) );
  NOR2_X1 U320 ( .A1(n16), .A2(n36), .ZN(ab_2__21_) );
  NOR2_X1 U321 ( .A1(n17), .A2(n36), .ZN(ab_2__20_) );
  NOR2_X1 U322 ( .A1(n18), .A2(n36), .ZN(ab_2__1_) );
  NOR2_X1 U323 ( .A1(n19), .A2(n36), .ZN(ab_2__19_) );
  NOR2_X1 U324 ( .A1(n20), .A2(n36), .ZN(ab_2__18_) );
  NOR2_X1 U325 ( .A1(n21), .A2(n36), .ZN(ab_2__17_) );
  NOR2_X1 U326 ( .A1(n22), .A2(n36), .ZN(ab_2__16_) );
  NOR2_X1 U327 ( .A1(n23), .A2(n36), .ZN(ab_2__15_) );
  NOR2_X1 U328 ( .A1(n24), .A2(n36), .ZN(ab_2__14_) );
  NOR2_X1 U329 ( .A1(n25), .A2(n36), .ZN(ab_2__13_) );
  NOR2_X1 U330 ( .A1(n26), .A2(n36), .ZN(ab_2__12_) );
  NOR2_X1 U331 ( .A1(n27), .A2(n36), .ZN(ab_2__11_) );
  NOR2_X1 U332 ( .A1(n28), .A2(n36), .ZN(ab_2__10_) );
  NOR2_X1 U333 ( .A1(n29), .A2(n36), .ZN(ab_2__0_) );
  NOR2_X1 U334 ( .A1(B[9]), .A2(n4), .ZN(ab_23__9_) );
  NOR2_X1 U335 ( .A1(B[8]), .A2(n4), .ZN(ab_23__8_) );
  NOR2_X1 U336 ( .A1(B[7]), .A2(n4), .ZN(ab_23__7_) );
  NOR2_X1 U337 ( .A1(B[6]), .A2(n4), .ZN(ab_23__6_) );
  NOR2_X1 U338 ( .A1(B[5]), .A2(n3), .ZN(ab_23__5_) );
  NOR2_X1 U339 ( .A1(B[4]), .A2(n3), .ZN(ab_23__4_) );
  NOR2_X1 U340 ( .A1(B[3]), .A2(n3), .ZN(ab_23__3_) );
  NOR2_X1 U341 ( .A1(B[2]), .A2(n3), .ZN(ab_23__2_) );
  NOR2_X1 U342 ( .A1(n1), .A2(n3), .ZN(ab_23__23_) );
  NOR2_X1 U343 ( .A1(B[22]), .A2(n3), .ZN(ab_23__22_) );
  NOR2_X1 U344 ( .A1(B[21]), .A2(n3), .ZN(ab_23__21_) );
  NOR2_X1 U345 ( .A1(B[20]), .A2(n3), .ZN(ab_23__20_) );
  NOR2_X1 U346 ( .A1(B[1]), .A2(n3), .ZN(ab_23__1_) );
  NOR2_X1 U347 ( .A1(B[19]), .A2(n3), .ZN(ab_23__19_) );
  NOR2_X1 U348 ( .A1(B[18]), .A2(n3), .ZN(ab_23__18_) );
  NOR2_X1 U349 ( .A1(B[17]), .A2(n3), .ZN(ab_23__17_) );
  NOR2_X1 U350 ( .A1(B[16]), .A2(n3), .ZN(ab_23__16_) );
  NOR2_X1 U351 ( .A1(B[15]), .A2(n3), .ZN(ab_23__15_) );
  NOR2_X1 U352 ( .A1(B[14]), .A2(n3), .ZN(ab_23__14_) );
  NOR2_X1 U353 ( .A1(B[13]), .A2(n3), .ZN(ab_23__13_) );
  NOR2_X1 U354 ( .A1(B[12]), .A2(n3), .ZN(ab_23__12_) );
  NOR2_X1 U355 ( .A1(B[11]), .A2(n3), .ZN(ab_23__11_) );
  NOR2_X1 U356 ( .A1(B[10]), .A2(n3), .ZN(ab_23__10_) );
  NOR2_X1 U357 ( .A1(B[0]), .A2(n3), .ZN(ab_23__0_) );
  NOR2_X1 U358 ( .A1(n7), .A2(n37), .ZN(ab_22__9_) );
  NOR2_X1 U359 ( .A1(n8), .A2(n37), .ZN(ab_22__8_) );
  NOR2_X1 U360 ( .A1(n9), .A2(n37), .ZN(ab_22__7_) );
  NOR2_X1 U361 ( .A1(n10), .A2(n37), .ZN(ab_22__6_) );
  NOR2_X1 U362 ( .A1(n11), .A2(n37), .ZN(ab_22__5_) );
  NOR2_X1 U363 ( .A1(n12), .A2(n37), .ZN(ab_22__4_) );
  NOR2_X1 U364 ( .A1(n13), .A2(n37), .ZN(ab_22__3_) );
  NOR2_X1 U365 ( .A1(n14), .A2(n37), .ZN(ab_22__2_) );
  NOR2_X1 U366 ( .A1(A[22]), .A2(n1), .ZN(ab_22__23_) );
  NOR2_X1 U367 ( .A1(n15), .A2(n37), .ZN(ab_22__22_) );
  NOR2_X1 U368 ( .A1(n16), .A2(n37), .ZN(ab_22__21_) );
  NOR2_X1 U369 ( .A1(n17), .A2(n37), .ZN(ab_22__20_) );
  NOR2_X1 U370 ( .A1(n18), .A2(n37), .ZN(ab_22__1_) );
  NOR2_X1 U371 ( .A1(n19), .A2(n37), .ZN(ab_22__19_) );
  NOR2_X1 U372 ( .A1(n20), .A2(n37), .ZN(ab_22__18_) );
  NOR2_X1 U373 ( .A1(n21), .A2(n37), .ZN(ab_22__17_) );
  NOR2_X1 U374 ( .A1(n22), .A2(n37), .ZN(ab_22__16_) );
  NOR2_X1 U375 ( .A1(n23), .A2(n37), .ZN(ab_22__15_) );
  NOR2_X1 U376 ( .A1(n24), .A2(n37), .ZN(ab_22__14_) );
  NOR2_X1 U377 ( .A1(n25), .A2(n37), .ZN(ab_22__13_) );
  NOR2_X1 U378 ( .A1(n26), .A2(n37), .ZN(ab_22__12_) );
  NOR2_X1 U379 ( .A1(n27), .A2(n37), .ZN(ab_22__11_) );
  NOR2_X1 U380 ( .A1(n28), .A2(n37), .ZN(ab_22__10_) );
  NOR2_X1 U381 ( .A1(n29), .A2(n37), .ZN(ab_22__0_) );
  NOR2_X1 U382 ( .A1(n7), .A2(n38), .ZN(ab_21__9_) );
  NOR2_X1 U383 ( .A1(n8), .A2(n38), .ZN(ab_21__8_) );
  NOR2_X1 U384 ( .A1(n9), .A2(n38), .ZN(ab_21__7_) );
  NOR2_X1 U385 ( .A1(n10), .A2(n38), .ZN(ab_21__6_) );
  NOR2_X1 U386 ( .A1(n11), .A2(n38), .ZN(ab_21__5_) );
  NOR2_X1 U387 ( .A1(n12), .A2(n38), .ZN(ab_21__4_) );
  NOR2_X1 U388 ( .A1(n13), .A2(n38), .ZN(ab_21__3_) );
  NOR2_X1 U389 ( .A1(n14), .A2(n38), .ZN(ab_21__2_) );
  NOR2_X1 U390 ( .A1(A[21]), .A2(n1), .ZN(ab_21__23_) );
  NOR2_X1 U391 ( .A1(n15), .A2(n38), .ZN(ab_21__22_) );
  NOR2_X1 U392 ( .A1(n16), .A2(n38), .ZN(ab_21__21_) );
  NOR2_X1 U393 ( .A1(n17), .A2(n38), .ZN(ab_21__20_) );
  NOR2_X1 U394 ( .A1(n18), .A2(n38), .ZN(ab_21__1_) );
  NOR2_X1 U395 ( .A1(n19), .A2(n38), .ZN(ab_21__19_) );
  NOR2_X1 U396 ( .A1(n20), .A2(n38), .ZN(ab_21__18_) );
  NOR2_X1 U397 ( .A1(n21), .A2(n38), .ZN(ab_21__17_) );
  NOR2_X1 U398 ( .A1(n22), .A2(n38), .ZN(ab_21__16_) );
  NOR2_X1 U399 ( .A1(n23), .A2(n38), .ZN(ab_21__15_) );
  NOR2_X1 U400 ( .A1(n24), .A2(n38), .ZN(ab_21__14_) );
  NOR2_X1 U401 ( .A1(n25), .A2(n38), .ZN(ab_21__13_) );
  NOR2_X1 U402 ( .A1(n26), .A2(n38), .ZN(ab_21__12_) );
  NOR2_X1 U403 ( .A1(n27), .A2(n38), .ZN(ab_21__11_) );
  NOR2_X1 U404 ( .A1(n28), .A2(n38), .ZN(ab_21__10_) );
  NOR2_X1 U405 ( .A1(n29), .A2(n38), .ZN(ab_21__0_) );
  NOR2_X1 U406 ( .A1(n7), .A2(n39), .ZN(ab_20__9_) );
  NOR2_X1 U407 ( .A1(n8), .A2(n39), .ZN(ab_20__8_) );
  NOR2_X1 U408 ( .A1(n9), .A2(n39), .ZN(ab_20__7_) );
  NOR2_X1 U409 ( .A1(n10), .A2(n39), .ZN(ab_20__6_) );
  NOR2_X1 U410 ( .A1(n11), .A2(n39), .ZN(ab_20__5_) );
  NOR2_X1 U411 ( .A1(n12), .A2(n39), .ZN(ab_20__4_) );
  NOR2_X1 U412 ( .A1(n13), .A2(n39), .ZN(ab_20__3_) );
  NOR2_X1 U413 ( .A1(n14), .A2(n39), .ZN(ab_20__2_) );
  NOR2_X1 U414 ( .A1(A[20]), .A2(n1), .ZN(ab_20__23_) );
  NOR2_X1 U415 ( .A1(n15), .A2(n39), .ZN(ab_20__22_) );
  NOR2_X1 U416 ( .A1(n16), .A2(n39), .ZN(ab_20__21_) );
  NOR2_X1 U417 ( .A1(n17), .A2(n39), .ZN(ab_20__20_) );
  NOR2_X1 U418 ( .A1(n18), .A2(n39), .ZN(ab_20__1_) );
  NOR2_X1 U419 ( .A1(n19), .A2(n39), .ZN(ab_20__19_) );
  NOR2_X1 U420 ( .A1(n20), .A2(n39), .ZN(ab_20__18_) );
  NOR2_X1 U421 ( .A1(n21), .A2(n39), .ZN(ab_20__17_) );
  NOR2_X1 U422 ( .A1(n22), .A2(n39), .ZN(ab_20__16_) );
  NOR2_X1 U423 ( .A1(n23), .A2(n39), .ZN(ab_20__15_) );
  NOR2_X1 U424 ( .A1(n24), .A2(n39), .ZN(ab_20__14_) );
  NOR2_X1 U425 ( .A1(n25), .A2(n39), .ZN(ab_20__13_) );
  NOR2_X1 U426 ( .A1(n26), .A2(n39), .ZN(ab_20__12_) );
  NOR2_X1 U427 ( .A1(n27), .A2(n39), .ZN(ab_20__11_) );
  NOR2_X1 U428 ( .A1(n28), .A2(n39), .ZN(ab_20__10_) );
  NOR2_X1 U429 ( .A1(n29), .A2(n39), .ZN(ab_20__0_) );
  NOR2_X1 U430 ( .A1(n7), .A2(n40), .ZN(ab_1__9_) );
  NOR2_X1 U431 ( .A1(n8), .A2(n40), .ZN(ab_1__8_) );
  NOR2_X1 U432 ( .A1(n9), .A2(n40), .ZN(ab_1__7_) );
  NOR2_X1 U433 ( .A1(n10), .A2(n40), .ZN(ab_1__6_) );
  NOR2_X1 U434 ( .A1(n11), .A2(n40), .ZN(ab_1__5_) );
  NOR2_X1 U435 ( .A1(n12), .A2(n40), .ZN(ab_1__4_) );
  NOR2_X1 U436 ( .A1(n13), .A2(n40), .ZN(ab_1__3_) );
  NOR2_X1 U437 ( .A1(n14), .A2(n40), .ZN(ab_1__2_) );
  NOR2_X1 U438 ( .A1(A[1]), .A2(n1), .ZN(ab_1__23_) );
  NOR2_X1 U439 ( .A1(n15), .A2(n40), .ZN(ab_1__22_) );
  NOR2_X1 U440 ( .A1(n16), .A2(n40), .ZN(ab_1__21_) );
  NOR2_X1 U441 ( .A1(n17), .A2(n40), .ZN(ab_1__20_) );
  NOR2_X1 U442 ( .A1(n19), .A2(n40), .ZN(ab_1__19_) );
  NOR2_X1 U443 ( .A1(n20), .A2(n40), .ZN(ab_1__18_) );
  NOR2_X1 U444 ( .A1(n21), .A2(n40), .ZN(ab_1__17_) );
  NOR2_X1 U445 ( .A1(n22), .A2(n40), .ZN(ab_1__16_) );
  NOR2_X1 U446 ( .A1(n23), .A2(n40), .ZN(ab_1__15_) );
  NOR2_X1 U447 ( .A1(n24), .A2(n40), .ZN(ab_1__14_) );
  NOR2_X1 U448 ( .A1(n25), .A2(n40), .ZN(ab_1__13_) );
  NOR2_X1 U449 ( .A1(n26), .A2(n40), .ZN(ab_1__12_) );
  NOR2_X1 U450 ( .A1(n27), .A2(n40), .ZN(ab_1__11_) );
  NOR2_X1 U451 ( .A1(n28), .A2(n40), .ZN(ab_1__10_) );
  NOR2_X1 U452 ( .A1(n7), .A2(n41), .ZN(ab_19__9_) );
  NOR2_X1 U453 ( .A1(n8), .A2(n41), .ZN(ab_19__8_) );
  NOR2_X1 U454 ( .A1(n9), .A2(n41), .ZN(ab_19__7_) );
  NOR2_X1 U455 ( .A1(n10), .A2(n41), .ZN(ab_19__6_) );
  NOR2_X1 U456 ( .A1(n11), .A2(n41), .ZN(ab_19__5_) );
  NOR2_X1 U457 ( .A1(n12), .A2(n41), .ZN(ab_19__4_) );
  NOR2_X1 U458 ( .A1(n13), .A2(n41), .ZN(ab_19__3_) );
  NOR2_X1 U459 ( .A1(n14), .A2(n41), .ZN(ab_19__2_) );
  NOR2_X1 U460 ( .A1(A[19]), .A2(n1), .ZN(ab_19__23_) );
  NOR2_X1 U461 ( .A1(n15), .A2(n41), .ZN(ab_19__22_) );
  NOR2_X1 U462 ( .A1(n16), .A2(n41), .ZN(ab_19__21_) );
  NOR2_X1 U463 ( .A1(n17), .A2(n41), .ZN(ab_19__20_) );
  NOR2_X1 U464 ( .A1(n18), .A2(n41), .ZN(ab_19__1_) );
  NOR2_X1 U465 ( .A1(n19), .A2(n41), .ZN(ab_19__19_) );
  NOR2_X1 U466 ( .A1(n20), .A2(n41), .ZN(ab_19__18_) );
  NOR2_X1 U467 ( .A1(n21), .A2(n41), .ZN(ab_19__17_) );
  NOR2_X1 U468 ( .A1(n22), .A2(n41), .ZN(ab_19__16_) );
  NOR2_X1 U469 ( .A1(n23), .A2(n41), .ZN(ab_19__15_) );
  NOR2_X1 U470 ( .A1(n24), .A2(n41), .ZN(ab_19__14_) );
  NOR2_X1 U471 ( .A1(n25), .A2(n41), .ZN(ab_19__13_) );
  NOR2_X1 U472 ( .A1(n26), .A2(n41), .ZN(ab_19__12_) );
  NOR2_X1 U473 ( .A1(n27), .A2(n41), .ZN(ab_19__11_) );
  NOR2_X1 U474 ( .A1(n28), .A2(n41), .ZN(ab_19__10_) );
  NOR2_X1 U475 ( .A1(n29), .A2(n41), .ZN(ab_19__0_) );
  NOR2_X1 U476 ( .A1(n7), .A2(n42), .ZN(ab_18__9_) );
  NOR2_X1 U477 ( .A1(n8), .A2(n42), .ZN(ab_18__8_) );
  NOR2_X1 U478 ( .A1(n9), .A2(n42), .ZN(ab_18__7_) );
  NOR2_X1 U479 ( .A1(n10), .A2(n42), .ZN(ab_18__6_) );
  NOR2_X1 U480 ( .A1(n11), .A2(n42), .ZN(ab_18__5_) );
  NOR2_X1 U481 ( .A1(n12), .A2(n42), .ZN(ab_18__4_) );
  NOR2_X1 U482 ( .A1(n13), .A2(n42), .ZN(ab_18__3_) );
  NOR2_X1 U483 ( .A1(n14), .A2(n42), .ZN(ab_18__2_) );
  NOR2_X1 U484 ( .A1(A[18]), .A2(n1), .ZN(ab_18__23_) );
  NOR2_X1 U485 ( .A1(n15), .A2(n42), .ZN(ab_18__22_) );
  NOR2_X1 U486 ( .A1(n16), .A2(n42), .ZN(ab_18__21_) );
  NOR2_X1 U487 ( .A1(n17), .A2(n42), .ZN(ab_18__20_) );
  NOR2_X1 U488 ( .A1(n18), .A2(n42), .ZN(ab_18__1_) );
  NOR2_X1 U489 ( .A1(n19), .A2(n42), .ZN(ab_18__19_) );
  NOR2_X1 U490 ( .A1(n20), .A2(n42), .ZN(ab_18__18_) );
  NOR2_X1 U491 ( .A1(n21), .A2(n42), .ZN(ab_18__17_) );
  NOR2_X1 U492 ( .A1(n22), .A2(n42), .ZN(ab_18__16_) );
  NOR2_X1 U493 ( .A1(n23), .A2(n42), .ZN(ab_18__15_) );
  NOR2_X1 U494 ( .A1(n24), .A2(n42), .ZN(ab_18__14_) );
  NOR2_X1 U495 ( .A1(n25), .A2(n42), .ZN(ab_18__13_) );
  NOR2_X1 U496 ( .A1(n26), .A2(n42), .ZN(ab_18__12_) );
  NOR2_X1 U497 ( .A1(n27), .A2(n42), .ZN(ab_18__11_) );
  NOR2_X1 U498 ( .A1(n28), .A2(n42), .ZN(ab_18__10_) );
  NOR2_X1 U499 ( .A1(n29), .A2(n42), .ZN(ab_18__0_) );
  NOR2_X1 U500 ( .A1(n7), .A2(n43), .ZN(ab_17__9_) );
  NOR2_X1 U501 ( .A1(n8), .A2(n43), .ZN(ab_17__8_) );
  NOR2_X1 U502 ( .A1(n9), .A2(n43), .ZN(ab_17__7_) );
  NOR2_X1 U503 ( .A1(n10), .A2(n43), .ZN(ab_17__6_) );
  NOR2_X1 U504 ( .A1(n11), .A2(n43), .ZN(ab_17__5_) );
  NOR2_X1 U505 ( .A1(n12), .A2(n43), .ZN(ab_17__4_) );
  NOR2_X1 U506 ( .A1(n13), .A2(n43), .ZN(ab_17__3_) );
  NOR2_X1 U507 ( .A1(n14), .A2(n43), .ZN(ab_17__2_) );
  NOR2_X1 U508 ( .A1(A[17]), .A2(n1), .ZN(ab_17__23_) );
  NOR2_X1 U509 ( .A1(n15), .A2(n43), .ZN(ab_17__22_) );
  NOR2_X1 U510 ( .A1(n16), .A2(n43), .ZN(ab_17__21_) );
  NOR2_X1 U511 ( .A1(n17), .A2(n43), .ZN(ab_17__20_) );
  NOR2_X1 U512 ( .A1(n18), .A2(n43), .ZN(ab_17__1_) );
  NOR2_X1 U513 ( .A1(n19), .A2(n43), .ZN(ab_17__19_) );
  NOR2_X1 U514 ( .A1(n20), .A2(n43), .ZN(ab_17__18_) );
  NOR2_X1 U515 ( .A1(n21), .A2(n43), .ZN(ab_17__17_) );
  NOR2_X1 U516 ( .A1(n22), .A2(n43), .ZN(ab_17__16_) );
  NOR2_X1 U517 ( .A1(n23), .A2(n43), .ZN(ab_17__15_) );
  NOR2_X1 U518 ( .A1(n24), .A2(n43), .ZN(ab_17__14_) );
  NOR2_X1 U519 ( .A1(n25), .A2(n43), .ZN(ab_17__13_) );
  NOR2_X1 U520 ( .A1(n26), .A2(n43), .ZN(ab_17__12_) );
  NOR2_X1 U521 ( .A1(n27), .A2(n43), .ZN(ab_17__11_) );
  NOR2_X1 U522 ( .A1(n28), .A2(n43), .ZN(ab_17__10_) );
  NOR2_X1 U523 ( .A1(n29), .A2(n43), .ZN(ab_17__0_) );
  NOR2_X1 U524 ( .A1(n7), .A2(n44), .ZN(ab_16__9_) );
  NOR2_X1 U525 ( .A1(n8), .A2(n44), .ZN(ab_16__8_) );
  NOR2_X1 U526 ( .A1(n9), .A2(n44), .ZN(ab_16__7_) );
  NOR2_X1 U527 ( .A1(n10), .A2(n44), .ZN(ab_16__6_) );
  NOR2_X1 U528 ( .A1(n11), .A2(n44), .ZN(ab_16__5_) );
  NOR2_X1 U529 ( .A1(n12), .A2(n44), .ZN(ab_16__4_) );
  NOR2_X1 U530 ( .A1(n13), .A2(n44), .ZN(ab_16__3_) );
  NOR2_X1 U531 ( .A1(n14), .A2(n44), .ZN(ab_16__2_) );
  NOR2_X1 U532 ( .A1(A[16]), .A2(n1), .ZN(ab_16__23_) );
  NOR2_X1 U533 ( .A1(n15), .A2(n44), .ZN(ab_16__22_) );
  NOR2_X1 U534 ( .A1(n16), .A2(n44), .ZN(ab_16__21_) );
  NOR2_X1 U535 ( .A1(n17), .A2(n44), .ZN(ab_16__20_) );
  NOR2_X1 U536 ( .A1(n18), .A2(n44), .ZN(ab_16__1_) );
  NOR2_X1 U537 ( .A1(n19), .A2(n44), .ZN(ab_16__19_) );
  NOR2_X1 U538 ( .A1(n20), .A2(n44), .ZN(ab_16__18_) );
  NOR2_X1 U539 ( .A1(n21), .A2(n44), .ZN(ab_16__17_) );
  NOR2_X1 U540 ( .A1(n22), .A2(n44), .ZN(ab_16__16_) );
  NOR2_X1 U541 ( .A1(n23), .A2(n44), .ZN(ab_16__15_) );
  NOR2_X1 U542 ( .A1(n24), .A2(n44), .ZN(ab_16__14_) );
  NOR2_X1 U543 ( .A1(n25), .A2(n44), .ZN(ab_16__13_) );
  NOR2_X1 U544 ( .A1(n26), .A2(n44), .ZN(ab_16__12_) );
  NOR2_X1 U545 ( .A1(n27), .A2(n44), .ZN(ab_16__11_) );
  NOR2_X1 U546 ( .A1(n28), .A2(n44), .ZN(ab_16__10_) );
  NOR2_X1 U547 ( .A1(n29), .A2(n44), .ZN(ab_16__0_) );
  NOR2_X1 U548 ( .A1(n7), .A2(n45), .ZN(ab_15__9_) );
  NOR2_X1 U549 ( .A1(n8), .A2(n45), .ZN(ab_15__8_) );
  NOR2_X1 U550 ( .A1(n9), .A2(n45), .ZN(ab_15__7_) );
  NOR2_X1 U551 ( .A1(n10), .A2(n45), .ZN(ab_15__6_) );
  NOR2_X1 U552 ( .A1(n11), .A2(n45), .ZN(ab_15__5_) );
  NOR2_X1 U553 ( .A1(n12), .A2(n45), .ZN(ab_15__4_) );
  NOR2_X1 U554 ( .A1(n13), .A2(n45), .ZN(ab_15__3_) );
  NOR2_X1 U555 ( .A1(n14), .A2(n45), .ZN(ab_15__2_) );
  NOR2_X1 U556 ( .A1(A[15]), .A2(n1), .ZN(ab_15__23_) );
  NOR2_X1 U557 ( .A1(n15), .A2(n45), .ZN(ab_15__22_) );
  NOR2_X1 U558 ( .A1(n16), .A2(n45), .ZN(ab_15__21_) );
  NOR2_X1 U559 ( .A1(n17), .A2(n45), .ZN(ab_15__20_) );
  NOR2_X1 U560 ( .A1(n18), .A2(n45), .ZN(ab_15__1_) );
  NOR2_X1 U561 ( .A1(n19), .A2(n45), .ZN(ab_15__19_) );
  NOR2_X1 U562 ( .A1(n20), .A2(n45), .ZN(ab_15__18_) );
  NOR2_X1 U563 ( .A1(n21), .A2(n45), .ZN(ab_15__17_) );
  NOR2_X1 U564 ( .A1(n22), .A2(n45), .ZN(ab_15__16_) );
  NOR2_X1 U565 ( .A1(n23), .A2(n45), .ZN(ab_15__15_) );
  NOR2_X1 U566 ( .A1(n24), .A2(n45), .ZN(ab_15__14_) );
  NOR2_X1 U567 ( .A1(n25), .A2(n45), .ZN(ab_15__13_) );
  NOR2_X1 U568 ( .A1(n26), .A2(n45), .ZN(ab_15__12_) );
  NOR2_X1 U569 ( .A1(n27), .A2(n45), .ZN(ab_15__11_) );
  NOR2_X1 U570 ( .A1(n28), .A2(n45), .ZN(ab_15__10_) );
  NOR2_X1 U571 ( .A1(n29), .A2(n45), .ZN(ab_15__0_) );
  NOR2_X1 U572 ( .A1(n7), .A2(n46), .ZN(ab_14__9_) );
  NOR2_X1 U573 ( .A1(n8), .A2(n46), .ZN(ab_14__8_) );
  NOR2_X1 U574 ( .A1(n9), .A2(n46), .ZN(ab_14__7_) );
  NOR2_X1 U575 ( .A1(n10), .A2(n46), .ZN(ab_14__6_) );
  NOR2_X1 U576 ( .A1(n11), .A2(n46), .ZN(ab_14__5_) );
  NOR2_X1 U577 ( .A1(n12), .A2(n46), .ZN(ab_14__4_) );
  NOR2_X1 U578 ( .A1(n13), .A2(n46), .ZN(ab_14__3_) );
  NOR2_X1 U579 ( .A1(n14), .A2(n46), .ZN(ab_14__2_) );
  NOR2_X1 U580 ( .A1(A[14]), .A2(n2), .ZN(ab_14__23_) );
  NOR2_X1 U581 ( .A1(n15), .A2(n46), .ZN(ab_14__22_) );
  NOR2_X1 U582 ( .A1(n16), .A2(n46), .ZN(ab_14__21_) );
  NOR2_X1 U583 ( .A1(n17), .A2(n46), .ZN(ab_14__20_) );
  NOR2_X1 U584 ( .A1(n18), .A2(n46), .ZN(ab_14__1_) );
  NOR2_X1 U585 ( .A1(n19), .A2(n46), .ZN(ab_14__19_) );
  NOR2_X1 U586 ( .A1(n20), .A2(n46), .ZN(ab_14__18_) );
  NOR2_X1 U587 ( .A1(n21), .A2(n46), .ZN(ab_14__17_) );
  NOR2_X1 U588 ( .A1(n22), .A2(n46), .ZN(ab_14__16_) );
  NOR2_X1 U589 ( .A1(n23), .A2(n46), .ZN(ab_14__15_) );
  NOR2_X1 U590 ( .A1(n24), .A2(n46), .ZN(ab_14__14_) );
  NOR2_X1 U591 ( .A1(n25), .A2(n46), .ZN(ab_14__13_) );
  NOR2_X1 U592 ( .A1(n26), .A2(n46), .ZN(ab_14__12_) );
  NOR2_X1 U593 ( .A1(n27), .A2(n46), .ZN(ab_14__11_) );
  NOR2_X1 U594 ( .A1(n28), .A2(n46), .ZN(ab_14__10_) );
  NOR2_X1 U595 ( .A1(n29), .A2(n46), .ZN(ab_14__0_) );
  NOR2_X1 U596 ( .A1(n7), .A2(n47), .ZN(ab_13__9_) );
  NOR2_X1 U597 ( .A1(n8), .A2(n47), .ZN(ab_13__8_) );
  NOR2_X1 U598 ( .A1(n9), .A2(n47), .ZN(ab_13__7_) );
  NOR2_X1 U599 ( .A1(n10), .A2(n47), .ZN(ab_13__6_) );
  NOR2_X1 U600 ( .A1(n11), .A2(n47), .ZN(ab_13__5_) );
  NOR2_X1 U601 ( .A1(n12), .A2(n47), .ZN(ab_13__4_) );
  NOR2_X1 U602 ( .A1(n13), .A2(n47), .ZN(ab_13__3_) );
  NOR2_X1 U603 ( .A1(n14), .A2(n47), .ZN(ab_13__2_) );
  NOR2_X1 U604 ( .A1(A[13]), .A2(n2), .ZN(ab_13__23_) );
  NOR2_X1 U605 ( .A1(n15), .A2(n47), .ZN(ab_13__22_) );
  NOR2_X1 U606 ( .A1(n16), .A2(n47), .ZN(ab_13__21_) );
  NOR2_X1 U607 ( .A1(n17), .A2(n47), .ZN(ab_13__20_) );
  NOR2_X1 U608 ( .A1(n18), .A2(n47), .ZN(ab_13__1_) );
  NOR2_X1 U609 ( .A1(n19), .A2(n47), .ZN(ab_13__19_) );
  NOR2_X1 U610 ( .A1(n20), .A2(n47), .ZN(ab_13__18_) );
  NOR2_X1 U611 ( .A1(n21), .A2(n47), .ZN(ab_13__17_) );
  NOR2_X1 U612 ( .A1(n22), .A2(n47), .ZN(ab_13__16_) );
  NOR2_X1 U613 ( .A1(n23), .A2(n47), .ZN(ab_13__15_) );
  NOR2_X1 U614 ( .A1(n24), .A2(n47), .ZN(ab_13__14_) );
  NOR2_X1 U615 ( .A1(n25), .A2(n47), .ZN(ab_13__13_) );
  NOR2_X1 U616 ( .A1(n26), .A2(n47), .ZN(ab_13__12_) );
  NOR2_X1 U617 ( .A1(n27), .A2(n47), .ZN(ab_13__11_) );
  NOR2_X1 U618 ( .A1(n28), .A2(n47), .ZN(ab_13__10_) );
  NOR2_X1 U619 ( .A1(n29), .A2(n47), .ZN(ab_13__0_) );
  NOR2_X1 U620 ( .A1(n7), .A2(n48), .ZN(ab_12__9_) );
  NOR2_X1 U621 ( .A1(n8), .A2(n48), .ZN(ab_12__8_) );
  NOR2_X1 U622 ( .A1(n9), .A2(n48), .ZN(ab_12__7_) );
  NOR2_X1 U623 ( .A1(n10), .A2(n48), .ZN(ab_12__6_) );
  NOR2_X1 U624 ( .A1(n11), .A2(n48), .ZN(ab_12__5_) );
  NOR2_X1 U625 ( .A1(n12), .A2(n48), .ZN(ab_12__4_) );
  NOR2_X1 U626 ( .A1(n13), .A2(n48), .ZN(ab_12__3_) );
  NOR2_X1 U627 ( .A1(n14), .A2(n48), .ZN(ab_12__2_) );
  NOR2_X1 U628 ( .A1(A[12]), .A2(n2), .ZN(ab_12__23_) );
  NOR2_X1 U629 ( .A1(n15), .A2(n48), .ZN(ab_12__22_) );
  NOR2_X1 U630 ( .A1(n16), .A2(n48), .ZN(ab_12__21_) );
  NOR2_X1 U631 ( .A1(n17), .A2(n48), .ZN(ab_12__20_) );
  NOR2_X1 U632 ( .A1(n18), .A2(n48), .ZN(ab_12__1_) );
  NOR2_X1 U633 ( .A1(n19), .A2(n48), .ZN(ab_12__19_) );
  NOR2_X1 U634 ( .A1(n20), .A2(n48), .ZN(ab_12__18_) );
  NOR2_X1 U635 ( .A1(n21), .A2(n48), .ZN(ab_12__17_) );
  NOR2_X1 U636 ( .A1(n22), .A2(n48), .ZN(ab_12__16_) );
  NOR2_X1 U637 ( .A1(n23), .A2(n48), .ZN(ab_12__15_) );
  NOR2_X1 U638 ( .A1(n24), .A2(n48), .ZN(ab_12__14_) );
  NOR2_X1 U639 ( .A1(n25), .A2(n48), .ZN(ab_12__13_) );
  NOR2_X1 U640 ( .A1(n26), .A2(n48), .ZN(ab_12__12_) );
  NOR2_X1 U641 ( .A1(n27), .A2(n48), .ZN(ab_12__11_) );
  NOR2_X1 U642 ( .A1(n28), .A2(n48), .ZN(ab_12__10_) );
  NOR2_X1 U643 ( .A1(n29), .A2(n48), .ZN(ab_12__0_) );
  NOR2_X1 U644 ( .A1(n7), .A2(n49), .ZN(ab_11__9_) );
  NOR2_X1 U645 ( .A1(n8), .A2(n49), .ZN(ab_11__8_) );
  NOR2_X1 U646 ( .A1(n9), .A2(n49), .ZN(ab_11__7_) );
  NOR2_X1 U647 ( .A1(n10), .A2(n49), .ZN(ab_11__6_) );
  NOR2_X1 U648 ( .A1(n11), .A2(n49), .ZN(ab_11__5_) );
  NOR2_X1 U649 ( .A1(n12), .A2(n49), .ZN(ab_11__4_) );
  NOR2_X1 U650 ( .A1(n13), .A2(n49), .ZN(ab_11__3_) );
  NOR2_X1 U651 ( .A1(n14), .A2(n49), .ZN(ab_11__2_) );
  NOR2_X1 U652 ( .A1(A[11]), .A2(n2), .ZN(ab_11__23_) );
  NOR2_X1 U653 ( .A1(n15), .A2(n49), .ZN(ab_11__22_) );
  NOR2_X1 U654 ( .A1(n16), .A2(n49), .ZN(ab_11__21_) );
  NOR2_X1 U655 ( .A1(n17), .A2(n49), .ZN(ab_11__20_) );
  NOR2_X1 U656 ( .A1(n18), .A2(n49), .ZN(ab_11__1_) );
  NOR2_X1 U657 ( .A1(n19), .A2(n49), .ZN(ab_11__19_) );
  NOR2_X1 U658 ( .A1(n20), .A2(n49), .ZN(ab_11__18_) );
  NOR2_X1 U659 ( .A1(n21), .A2(n49), .ZN(ab_11__17_) );
  NOR2_X1 U660 ( .A1(n22), .A2(n49), .ZN(ab_11__16_) );
  NOR2_X1 U661 ( .A1(n23), .A2(n49), .ZN(ab_11__15_) );
  NOR2_X1 U662 ( .A1(n24), .A2(n49), .ZN(ab_11__14_) );
  NOR2_X1 U663 ( .A1(n25), .A2(n49), .ZN(ab_11__13_) );
  NOR2_X1 U664 ( .A1(n26), .A2(n49), .ZN(ab_11__12_) );
  NOR2_X1 U665 ( .A1(n27), .A2(n49), .ZN(ab_11__11_) );
  NOR2_X1 U666 ( .A1(n28), .A2(n49), .ZN(ab_11__10_) );
  NOR2_X1 U667 ( .A1(n29), .A2(n49), .ZN(ab_11__0_) );
  NOR2_X1 U668 ( .A1(n7), .A2(n50), .ZN(ab_10__9_) );
  NOR2_X1 U669 ( .A1(n8), .A2(n50), .ZN(ab_10__8_) );
  NOR2_X1 U670 ( .A1(n9), .A2(n50), .ZN(ab_10__7_) );
  NOR2_X1 U671 ( .A1(n10), .A2(n50), .ZN(ab_10__6_) );
  NOR2_X1 U672 ( .A1(n11), .A2(n50), .ZN(ab_10__5_) );
  NOR2_X1 U673 ( .A1(n12), .A2(n50), .ZN(ab_10__4_) );
  NOR2_X1 U674 ( .A1(n13), .A2(n50), .ZN(ab_10__3_) );
  NOR2_X1 U675 ( .A1(n14), .A2(n50), .ZN(ab_10__2_) );
  NOR2_X1 U676 ( .A1(A[10]), .A2(n2), .ZN(ab_10__23_) );
  NOR2_X1 U677 ( .A1(n15), .A2(n50), .ZN(ab_10__22_) );
  NOR2_X1 U678 ( .A1(n16), .A2(n50), .ZN(ab_10__21_) );
  NOR2_X1 U679 ( .A1(n17), .A2(n50), .ZN(ab_10__20_) );
  NOR2_X1 U680 ( .A1(n18), .A2(n50), .ZN(ab_10__1_) );
  NOR2_X1 U681 ( .A1(n19), .A2(n50), .ZN(ab_10__19_) );
  NOR2_X1 U682 ( .A1(n20), .A2(n50), .ZN(ab_10__18_) );
  NOR2_X1 U683 ( .A1(n21), .A2(n50), .ZN(ab_10__17_) );
  NOR2_X1 U684 ( .A1(n22), .A2(n50), .ZN(ab_10__16_) );
  NOR2_X1 U685 ( .A1(n23), .A2(n50), .ZN(ab_10__15_) );
  NOR2_X1 U686 ( .A1(n24), .A2(n50), .ZN(ab_10__14_) );
  NOR2_X1 U687 ( .A1(n25), .A2(n50), .ZN(ab_10__13_) );
  NOR2_X1 U688 ( .A1(n26), .A2(n50), .ZN(ab_10__12_) );
  NOR2_X1 U689 ( .A1(n27), .A2(n50), .ZN(ab_10__11_) );
  NOR2_X1 U690 ( .A1(n28), .A2(n50), .ZN(ab_10__10_) );
  NOR2_X1 U691 ( .A1(n29), .A2(n50), .ZN(ab_10__0_) );
  NOR2_X1 U692 ( .A1(n7), .A2(n51), .ZN(ab_0__9_) );
  NOR2_X1 U693 ( .A1(n8), .A2(n51), .ZN(ab_0__8_) );
  NOR2_X1 U694 ( .A1(n9), .A2(n51), .ZN(ab_0__7_) );
  NOR2_X1 U695 ( .A1(n10), .A2(n51), .ZN(ab_0__6_) );
  NOR2_X1 U696 ( .A1(n11), .A2(n51), .ZN(ab_0__5_) );
  NOR2_X1 U697 ( .A1(n12), .A2(n51), .ZN(ab_0__4_) );
  NOR2_X1 U698 ( .A1(n13), .A2(n51), .ZN(ab_0__3_) );
  NOR2_X1 U699 ( .A1(n14), .A2(n51), .ZN(ab_0__2_) );
  NOR2_X1 U700 ( .A1(A[0]), .A2(n1), .ZN(ab_0__23_) );
  NOR2_X1 U701 ( .A1(n15), .A2(n51), .ZN(ab_0__22_) );
  NOR2_X1 U702 ( .A1(n16), .A2(n51), .ZN(ab_0__21_) );
  NOR2_X1 U703 ( .A1(n17), .A2(n51), .ZN(ab_0__20_) );
  NOR2_X1 U704 ( .A1(n19), .A2(n51), .ZN(ab_0__19_) );
  NOR2_X1 U705 ( .A1(n20), .A2(n51), .ZN(ab_0__18_) );
  NOR2_X1 U706 ( .A1(n21), .A2(n51), .ZN(ab_0__17_) );
  NOR2_X1 U707 ( .A1(n22), .A2(n51), .ZN(ab_0__16_) );
  NOR2_X1 U708 ( .A1(n23), .A2(n51), .ZN(ab_0__15_) );
  NOR2_X1 U709 ( .A1(n24), .A2(n51), .ZN(ab_0__14_) );
  NOR2_X1 U710 ( .A1(n25), .A2(n51), .ZN(ab_0__13_) );
  NOR2_X1 U711 ( .A1(n26), .A2(n51), .ZN(ab_0__12_) );
  NOR2_X1 U712 ( .A1(n27), .A2(n51), .ZN(ab_0__11_) );
  NOR2_X1 U713 ( .A1(n28), .A2(n51), .ZN(ab_0__10_) );
  INV_X1 U714 ( .A(B[23]), .ZN(QB) );
  INV_X1 U715 ( .A(A[23]), .ZN(QA) );
  AND3_X1 U716 ( .A1(ab_1__1_), .A2(B[0]), .A3(A[0]), .ZN(CARRYB_1__0_) );
  NOR2_X1 U717 ( .A1(n40), .A2(n18), .ZN(ab_1__1_) );
  INV_X1 U719 ( .A(CARRYB_23__23_), .ZN(A1_45_) );
endmodule


module iir_filter_DW01_add_8 ( A, B, CI, SUM, CO );
  input [45:0] A;
  input [45:0] B;
  output [45:0] SUM;
  input CI;
  output CO;
  wire   A_21_, A_20_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112;
  assign SUM[21] = A_21_;
  assign A_21_ = A[21];
  assign SUM[20] = A_20_;
  assign A_20_ = A[20];

  XOR2_X1 U2 ( .A(n1), .B(n2), .Z(SUM[45]) );
  XOR2_X1 U3 ( .A(B[45]), .B(A[45]), .Z(n2) );
  OAI21_X1 U4 ( .B1(n3), .B2(n4), .A(n5), .ZN(n1) );
  OAI21_X1 U5 ( .B1(A[44]), .B2(n6), .A(B[44]), .ZN(n5) );
  INV_X1 U6 ( .A(n3), .ZN(n6) );
  INV_X1 U7 ( .A(A[44]), .ZN(n4) );
  AOI21_X1 U8 ( .B1(A[43]), .B2(B[43]), .A(n7), .ZN(n3) );
  INV_X1 U9 ( .A(n8), .ZN(n7) );
  OAI22_X1 U10 ( .A1(n9), .A2(n10), .B1(A[43]), .B2(B[43]), .ZN(n8) );
  AOI21_X1 U11 ( .B1(n11), .B2(n12), .A(n13), .ZN(n9) );
  NAND3_X1 U12 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n12) );
  AOI21_X1 U13 ( .B1(n17), .B2(n16), .A(n18), .ZN(n11) );
  INV_X1 U14 ( .A(n19), .ZN(n18) );
  XOR2_X1 U15 ( .A(n20), .B(n21), .Z(SUM[42]) );
  NOR2_X1 U16 ( .A1(n10), .A2(n13), .ZN(n21) );
  NOR2_X1 U17 ( .A1(B[42]), .A2(A[42]), .ZN(n13) );
  AND2_X1 U18 ( .A1(B[42]), .A2(A[42]), .ZN(n10) );
  OAI21_X1 U19 ( .B1(n22), .B2(n23), .A(n19), .ZN(n20) );
  XOR2_X1 U20 ( .A(n24), .B(n23), .Z(SUM[41]) );
  AOI21_X1 U21 ( .B1(n15), .B2(n14), .A(n17), .ZN(n23) );
  INV_X1 U22 ( .A(n25), .ZN(n15) );
  NAND2_X1 U23 ( .A1(n16), .A2(n19), .ZN(n24) );
  NAND2_X1 U24 ( .A1(B[41]), .A2(A[41]), .ZN(n19) );
  INV_X1 U25 ( .A(n22), .ZN(n16) );
  NOR2_X1 U26 ( .A1(B[41]), .A2(A[41]), .ZN(n22) );
  XOR2_X1 U27 ( .A(n14), .B(n26), .Z(SUM[40]) );
  NOR2_X1 U28 ( .A1(n17), .A2(n25), .ZN(n26) );
  NOR2_X1 U29 ( .A1(B[40]), .A2(A[40]), .ZN(n25) );
  AND2_X1 U30 ( .A1(B[40]), .A2(A[40]), .ZN(n17) );
  OAI21_X1 U31 ( .B1(n27), .B2(n28), .A(n29), .ZN(n14) );
  XOR2_X1 U32 ( .A(n30), .B(n28), .Z(SUM[39]) );
  AOI21_X1 U33 ( .B1(n31), .B2(n32), .A(n33), .ZN(n28) );
  INV_X1 U34 ( .A(n34), .ZN(n31) );
  NAND2_X1 U35 ( .A1(n35), .A2(n29), .ZN(n30) );
  NAND2_X1 U36 ( .A1(B[39]), .A2(A[39]), .ZN(n29) );
  INV_X1 U37 ( .A(n27), .ZN(n35) );
  NOR2_X1 U38 ( .A1(B[39]), .A2(A[39]), .ZN(n27) );
  XOR2_X1 U39 ( .A(n32), .B(n36), .Z(SUM[38]) );
  NOR2_X1 U40 ( .A1(n33), .A2(n34), .ZN(n36) );
  NOR2_X1 U41 ( .A1(B[38]), .A2(A[38]), .ZN(n34) );
  AND2_X1 U42 ( .A1(B[38]), .A2(A[38]), .ZN(n33) );
  OAI21_X1 U43 ( .B1(n37), .B2(n38), .A(n39), .ZN(n32) );
  XOR2_X1 U44 ( .A(n40), .B(n38), .Z(SUM[37]) );
  AOI21_X1 U45 ( .B1(n41), .B2(n42), .A(n43), .ZN(n38) );
  INV_X1 U46 ( .A(n44), .ZN(n41) );
  NAND2_X1 U47 ( .A1(n45), .A2(n39), .ZN(n40) );
  NAND2_X1 U48 ( .A1(B[37]), .A2(A[37]), .ZN(n39) );
  INV_X1 U49 ( .A(n37), .ZN(n45) );
  NOR2_X1 U50 ( .A1(B[37]), .A2(A[37]), .ZN(n37) );
  XOR2_X1 U51 ( .A(n42), .B(n46), .Z(SUM[36]) );
  NOR2_X1 U52 ( .A1(n43), .A2(n44), .ZN(n46) );
  NOR2_X1 U53 ( .A1(B[36]), .A2(A[36]), .ZN(n44) );
  AND2_X1 U54 ( .A1(B[36]), .A2(A[36]), .ZN(n43) );
  OAI21_X1 U55 ( .B1(n47), .B2(n48), .A(n49), .ZN(n42) );
  XOR2_X1 U56 ( .A(n50), .B(n48), .Z(SUM[35]) );
  AOI21_X1 U57 ( .B1(n51), .B2(n52), .A(n53), .ZN(n48) );
  INV_X1 U58 ( .A(n54), .ZN(n51) );
  NAND2_X1 U59 ( .A1(n55), .A2(n49), .ZN(n50) );
  NAND2_X1 U60 ( .A1(B[35]), .A2(A[35]), .ZN(n49) );
  INV_X1 U61 ( .A(n47), .ZN(n55) );
  NOR2_X1 U62 ( .A1(B[35]), .A2(A[35]), .ZN(n47) );
  XOR2_X1 U63 ( .A(n52), .B(n56), .Z(SUM[34]) );
  NOR2_X1 U64 ( .A1(n53), .A2(n54), .ZN(n56) );
  NOR2_X1 U65 ( .A1(B[34]), .A2(A[34]), .ZN(n54) );
  AND2_X1 U66 ( .A1(B[34]), .A2(A[34]), .ZN(n53) );
  OAI21_X1 U67 ( .B1(n57), .B2(n58), .A(n59), .ZN(n52) );
  XOR2_X1 U68 ( .A(n60), .B(n58), .Z(SUM[33]) );
  AOI21_X1 U69 ( .B1(n61), .B2(n62), .A(n63), .ZN(n58) );
  INV_X1 U70 ( .A(n64), .ZN(n61) );
  NAND2_X1 U71 ( .A1(n65), .A2(n59), .ZN(n60) );
  NAND2_X1 U72 ( .A1(B[33]), .A2(A[33]), .ZN(n59) );
  INV_X1 U73 ( .A(n57), .ZN(n65) );
  NOR2_X1 U74 ( .A1(B[33]), .A2(A[33]), .ZN(n57) );
  XOR2_X1 U75 ( .A(n62), .B(n66), .Z(SUM[32]) );
  NOR2_X1 U76 ( .A1(n63), .A2(n64), .ZN(n66) );
  NOR2_X1 U77 ( .A1(B[32]), .A2(A[32]), .ZN(n64) );
  AND2_X1 U78 ( .A1(B[32]), .A2(A[32]), .ZN(n63) );
  OAI21_X1 U79 ( .B1(n67), .B2(n68), .A(n69), .ZN(n62) );
  XOR2_X1 U80 ( .A(n70), .B(n68), .Z(SUM[31]) );
  AOI21_X1 U81 ( .B1(n71), .B2(n72), .A(n73), .ZN(n68) );
  INV_X1 U82 ( .A(n74), .ZN(n71) );
  NAND2_X1 U83 ( .A1(n75), .A2(n69), .ZN(n70) );
  NAND2_X1 U84 ( .A1(B[31]), .A2(A[31]), .ZN(n69) );
  INV_X1 U85 ( .A(n67), .ZN(n75) );
  NOR2_X1 U86 ( .A1(B[31]), .A2(A[31]), .ZN(n67) );
  XOR2_X1 U87 ( .A(n72), .B(n76), .Z(SUM[30]) );
  NOR2_X1 U88 ( .A1(n73), .A2(n74), .ZN(n76) );
  NOR2_X1 U89 ( .A1(B[30]), .A2(A[30]), .ZN(n74) );
  AND2_X1 U90 ( .A1(B[30]), .A2(A[30]), .ZN(n73) );
  OAI21_X1 U91 ( .B1(n77), .B2(n78), .A(n79), .ZN(n72) );
  XOR2_X1 U92 ( .A(n80), .B(n78), .Z(SUM[29]) );
  AOI21_X1 U93 ( .B1(n81), .B2(n82), .A(n83), .ZN(n78) );
  INV_X1 U94 ( .A(n84), .ZN(n81) );
  NAND2_X1 U95 ( .A1(n85), .A2(n79), .ZN(n80) );
  NAND2_X1 U96 ( .A1(B[29]), .A2(A[29]), .ZN(n79) );
  INV_X1 U97 ( .A(n77), .ZN(n85) );
  NOR2_X1 U98 ( .A1(B[29]), .A2(A[29]), .ZN(n77) );
  XOR2_X1 U99 ( .A(n82), .B(n86), .Z(SUM[28]) );
  NOR2_X1 U100 ( .A1(n83), .A2(n84), .ZN(n86) );
  NOR2_X1 U101 ( .A1(B[28]), .A2(A[28]), .ZN(n84) );
  AND2_X1 U102 ( .A1(B[28]), .A2(A[28]), .ZN(n83) );
  OAI21_X1 U103 ( .B1(n87), .B2(n88), .A(n89), .ZN(n82) );
  XOR2_X1 U104 ( .A(n90), .B(n88), .Z(SUM[27]) );
  AOI21_X1 U105 ( .B1(n91), .B2(n92), .A(n93), .ZN(n88) );
  INV_X1 U106 ( .A(n94), .ZN(n92) );
  NAND2_X1 U107 ( .A1(n95), .A2(n89), .ZN(n90) );
  NAND2_X1 U108 ( .A1(B[27]), .A2(A[27]), .ZN(n89) );
  INV_X1 U109 ( .A(n87), .ZN(n95) );
  NOR2_X1 U110 ( .A1(B[27]), .A2(A[27]), .ZN(n87) );
  XOR2_X1 U111 ( .A(n91), .B(n96), .Z(SUM[26]) );
  NOR2_X1 U112 ( .A1(n93), .A2(n94), .ZN(n96) );
  NOR2_X1 U113 ( .A1(B[26]), .A2(A[26]), .ZN(n94) );
  AND2_X1 U114 ( .A1(B[26]), .A2(A[26]), .ZN(n93) );
  OAI21_X1 U115 ( .B1(n97), .B2(n98), .A(n99), .ZN(n91) );
  XOR2_X1 U116 ( .A(n100), .B(n98), .Z(SUM[25]) );
  AOI21_X1 U117 ( .B1(n101), .B2(n102), .A(n103), .ZN(n98) );
  INV_X1 U118 ( .A(n104), .ZN(n101) );
  NAND2_X1 U119 ( .A1(n105), .A2(n99), .ZN(n100) );
  NAND2_X1 U120 ( .A1(B[25]), .A2(A[25]), .ZN(n99) );
  INV_X1 U121 ( .A(n97), .ZN(n105) );
  NOR2_X1 U122 ( .A1(B[25]), .A2(A[25]), .ZN(n97) );
  XOR2_X1 U123 ( .A(n102), .B(n106), .Z(SUM[24]) );
  NOR2_X1 U124 ( .A1(n103), .A2(n104), .ZN(n106) );
  NOR2_X1 U125 ( .A1(B[24]), .A2(A[24]), .ZN(n104) );
  AND2_X1 U126 ( .A1(B[24]), .A2(A[24]), .ZN(n103) );
  OAI21_X1 U127 ( .B1(n107), .B2(n108), .A(n109), .ZN(n102) );
  XOR2_X1 U128 ( .A(n108), .B(n110), .Z(SUM[23]) );
  NAND2_X1 U129 ( .A1(n111), .A2(n109), .ZN(n110) );
  NAND2_X1 U130 ( .A1(B[23]), .A2(A[23]), .ZN(n109) );
  INV_X1 U131 ( .A(n107), .ZN(n111) );
  NOR2_X1 U132 ( .A1(B[23]), .A2(A[23]), .ZN(n107) );
  INV_X1 U133 ( .A(n112), .ZN(SUM[22]) );
  OAI21_X1 U134 ( .B1(B[22]), .B2(A[22]), .A(n108), .ZN(n112) );
  NAND2_X1 U135 ( .A1(B[22]), .A2(A[22]), .ZN(n108) );
endmodule


module iir_filter_DW02_mult_4 ( A, B, TC, PRODUCT );
  input [23:0] A;
  input [23:0] B;
  output [47:0] PRODUCT;
  input TC;
  wire   ab_23__23_, ab_23__22_, ab_23__21_, ab_23__20_, ab_23__19_,
         ab_23__18_, ab_23__17_, ab_23__16_, ab_23__15_, ab_23__14_,
         ab_23__13_, ab_23__12_, ab_23__11_, ab_23__10_, ab_23__9_, ab_23__8_,
         ab_23__7_, ab_23__6_, ab_23__5_, ab_23__4_, ab_23__3_, ab_23__2_,
         ab_23__1_, ab_23__0_, ab_22__23_, ab_22__22_, ab_22__21_, ab_22__20_,
         ab_22__19_, ab_22__18_, ab_22__17_, ab_22__16_, ab_22__15_,
         ab_22__14_, ab_22__13_, ab_22__12_, ab_22__11_, ab_22__10_, ab_22__9_,
         ab_22__8_, ab_22__7_, ab_22__6_, ab_22__5_, ab_22__4_, ab_22__3_,
         ab_22__2_, ab_22__1_, ab_22__0_, ab_21__23_, ab_21__22_, ab_21__21_,
         ab_21__20_, ab_21__19_, ab_21__18_, ab_21__17_, ab_21__16_,
         ab_21__15_, ab_21__14_, ab_21__13_, ab_21__12_, ab_21__11_,
         ab_21__10_, ab_21__9_, ab_21__8_, ab_21__7_, ab_21__6_, ab_21__5_,
         ab_21__4_, ab_21__3_, ab_21__2_, ab_21__1_, ab_21__0_, ab_20__23_,
         ab_20__22_, ab_20__21_, ab_20__20_, ab_20__19_, ab_20__18_,
         ab_20__17_, ab_20__16_, ab_20__15_, ab_20__14_, ab_20__13_,
         ab_20__12_, ab_20__11_, ab_20__10_, ab_20__9_, ab_20__8_, ab_20__7_,
         ab_20__6_, ab_20__5_, ab_20__4_, ab_20__3_, ab_20__2_, ab_20__1_,
         ab_20__0_, ab_19__23_, ab_19__22_, ab_19__21_, ab_19__20_, ab_19__19_,
         ab_19__18_, ab_19__17_, ab_19__16_, ab_19__15_, ab_19__14_,
         ab_19__13_, ab_19__12_, ab_19__11_, ab_19__10_, ab_19__9_, ab_19__8_,
         ab_19__7_, ab_19__6_, ab_19__5_, ab_19__4_, ab_19__3_, ab_19__2_,
         ab_19__1_, ab_19__0_, ab_18__23_, ab_18__22_, ab_18__21_, ab_18__20_,
         ab_18__19_, ab_18__18_, ab_18__17_, ab_18__16_, ab_18__15_,
         ab_18__14_, ab_18__13_, ab_18__12_, ab_18__11_, ab_18__10_, ab_18__9_,
         ab_18__8_, ab_18__7_, ab_18__6_, ab_18__5_, ab_18__4_, ab_18__3_,
         ab_18__2_, ab_18__1_, ab_18__0_, ab_17__23_, ab_17__22_, ab_17__21_,
         ab_17__20_, ab_17__19_, ab_17__18_, ab_17__17_, ab_17__16_,
         ab_17__15_, ab_17__14_, ab_17__13_, ab_17__12_, ab_17__11_,
         ab_17__10_, ab_17__9_, ab_17__8_, ab_17__7_, ab_17__6_, ab_17__5_,
         ab_17__4_, ab_17__3_, ab_17__2_, ab_17__1_, ab_17__0_, ab_16__23_,
         ab_16__22_, ab_16__21_, ab_16__20_, ab_16__19_, ab_16__18_,
         ab_16__17_, ab_16__16_, ab_16__15_, ab_16__14_, ab_16__13_,
         ab_16__12_, ab_16__11_, ab_16__10_, ab_16__9_, ab_16__8_, ab_16__7_,
         ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_, ab_16__1_,
         ab_16__0_, ab_15__23_, ab_15__22_, ab_15__21_, ab_15__20_, ab_15__19_,
         ab_15__18_, ab_15__17_, ab_15__16_, ab_15__15_, ab_15__14_,
         ab_15__13_, ab_15__12_, ab_15__11_, ab_15__10_, ab_15__9_, ab_15__8_,
         ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_, ab_15__3_, ab_15__2_,
         ab_15__1_, ab_15__0_, ab_14__23_, ab_14__22_, ab_14__21_, ab_14__20_,
         ab_14__19_, ab_14__18_, ab_14__17_, ab_14__16_, ab_14__15_,
         ab_14__14_, ab_14__13_, ab_14__12_, ab_14__11_, ab_14__10_, ab_14__9_,
         ab_14__8_, ab_14__7_, ab_14__6_, ab_14__5_, ab_14__4_, ab_14__3_,
         ab_14__2_, ab_14__1_, ab_14__0_, ab_13__23_, ab_13__22_, ab_13__21_,
         ab_13__20_, ab_13__19_, ab_13__18_, ab_13__17_, ab_13__16_,
         ab_13__15_, ab_13__14_, ab_13__13_, ab_13__12_, ab_13__11_,
         ab_13__10_, ab_13__9_, ab_13__8_, ab_13__7_, ab_13__6_, ab_13__5_,
         ab_13__4_, ab_13__3_, ab_13__2_, ab_13__1_, ab_13__0_, ab_12__23_,
         ab_12__22_, ab_12__21_, ab_12__20_, ab_12__19_, ab_12__18_,
         ab_12__17_, ab_12__16_, ab_12__15_, ab_12__14_, ab_12__13_,
         ab_12__12_, ab_12__11_, ab_12__10_, ab_12__9_, ab_12__8_, ab_12__7_,
         ab_12__6_, ab_12__5_, ab_12__4_, ab_12__3_, ab_12__2_, ab_12__1_,
         ab_12__0_, ab_11__23_, ab_11__22_, ab_11__21_, ab_11__20_, ab_11__19_,
         ab_11__18_, ab_11__17_, ab_11__16_, ab_11__15_, ab_11__14_,
         ab_11__13_, ab_11__12_, ab_11__11_, ab_11__10_, ab_11__9_, ab_11__8_,
         ab_11__7_, ab_11__6_, ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_,
         ab_11__1_, ab_11__0_, ab_10__23_, ab_10__22_, ab_10__21_, ab_10__20_,
         ab_10__19_, ab_10__18_, ab_10__17_, ab_10__16_, ab_10__15_,
         ab_10__14_, ab_10__13_, ab_10__12_, ab_10__11_, ab_10__10_, ab_10__9_,
         ab_10__8_, ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_,
         ab_10__2_, ab_10__1_, ab_10__0_, ab_9__23_, ab_9__22_, ab_9__21_,
         ab_9__20_, ab_9__19_, ab_9__18_, ab_9__17_, ab_9__16_, ab_9__15_,
         ab_9__14_, ab_9__13_, ab_9__12_, ab_9__11_, ab_9__10_, ab_9__9_,
         ab_9__8_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_,
         ab_9__1_, ab_9__0_, ab_8__23_, ab_8__22_, ab_8__21_, ab_8__20_,
         ab_8__19_, ab_8__18_, ab_8__17_, ab_8__16_, ab_8__15_, ab_8__14_,
         ab_8__13_, ab_8__12_, ab_8__11_, ab_8__10_, ab_8__9_, ab_8__8_,
         ab_8__7_, ab_8__6_, ab_8__5_, ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_,
         ab_8__0_, ab_7__23_, ab_7__22_, ab_7__21_, ab_7__20_, ab_7__19_,
         ab_7__18_, ab_7__17_, ab_7__16_, ab_7__15_, ab_7__14_, ab_7__13_,
         ab_7__12_, ab_7__11_, ab_7__10_, ab_7__9_, ab_7__8_, ab_7__7_,
         ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_,
         ab_6__23_, ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_, ab_6__18_,
         ab_6__17_, ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_, ab_6__12_,
         ab_6__11_, ab_6__10_, ab_6__9_, ab_6__8_, ab_6__7_, ab_6__6_,
         ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_, ab_5__23_,
         ab_5__22_, ab_5__21_, ab_5__20_, ab_5__19_, ab_5__18_, ab_5__17_,
         ab_5__16_, ab_5__15_, ab_5__14_, ab_5__13_, ab_5__12_, ab_5__11_,
         ab_5__10_, ab_5__9_, ab_5__8_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_,
         ab_5__3_, ab_5__2_, ab_5__1_, ab_5__0_, ab_4__23_, ab_4__22_,
         ab_4__21_, ab_4__20_, ab_4__19_, ab_4__18_, ab_4__17_, ab_4__16_,
         ab_4__15_, ab_4__14_, ab_4__13_, ab_4__12_, ab_4__11_, ab_4__10_,
         ab_4__9_, ab_4__8_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_,
         ab_4__2_, ab_4__1_, ab_4__0_, ab_3__23_, ab_3__22_, ab_3__21_,
         ab_3__20_, ab_3__19_, ab_3__18_, ab_3__17_, ab_3__16_, ab_3__15_,
         ab_3__14_, ab_3__13_, ab_3__12_, ab_3__11_, ab_3__10_, ab_3__9_,
         ab_3__8_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_, ab_3__2_,
         ab_3__1_, ab_3__0_, ab_2__23_, ab_2__22_, ab_2__21_, ab_2__20_,
         ab_2__19_, ab_2__18_, ab_2__17_, ab_2__16_, ab_2__15_, ab_2__14_,
         ab_2__13_, ab_2__12_, ab_2__11_, ab_2__10_, ab_2__9_, ab_2__8_,
         ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_,
         ab_2__0_, ab_1__23_, ab_1__22_, ab_1__21_, ab_1__20_, ab_1__19_,
         ab_1__18_, ab_1__17_, ab_1__16_, ab_1__15_, ab_1__14_, ab_1__13_,
         ab_1__12_, ab_1__11_, ab_1__10_, ab_1__9_, ab_1__8_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_0__23_,
         ab_0__22_, ab_0__21_, ab_0__20_, ab_0__19_, ab_0__18_, ab_0__17_,
         ab_0__16_, ab_0__15_, ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_,
         ab_0__10_, ab_0__9_, ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_23__23_, CARRYB_23__22_, CARRYB_23__21_,
         CARRYB_23__20_, CARRYB_23__19_, CARRYB_23__18_, CARRYB_23__17_,
         CARRYB_23__16_, CARRYB_23__15_, CARRYB_23__14_, CARRYB_23__13_,
         CARRYB_23__12_, CARRYB_23__11_, CARRYB_23__10_, CARRYB_23__9_,
         CARRYB_23__8_, CARRYB_23__7_, CARRYB_23__6_, CARRYB_23__5_,
         CARRYB_23__4_, CARRYB_23__3_, CARRYB_23__2_, CARRYB_23__1_,
         CARRYB_23__0_, CARRYB_22__22_, CARRYB_22__21_, CARRYB_22__20_,
         CARRYB_22__19_, CARRYB_22__18_, CARRYB_22__17_, CARRYB_22__16_,
         CARRYB_22__15_, CARRYB_22__14_, CARRYB_22__13_, CARRYB_22__12_,
         CARRYB_22__11_, CARRYB_22__10_, CARRYB_22__9_, CARRYB_22__8_,
         CARRYB_22__7_, CARRYB_22__6_, CARRYB_22__5_, CARRYB_22__4_,
         CARRYB_22__3_, CARRYB_22__2_, CARRYB_22__1_, CARRYB_22__0_,
         CARRYB_21__22_, CARRYB_21__21_, CARRYB_21__20_, CARRYB_21__19_,
         CARRYB_21__18_, CARRYB_21__17_, CARRYB_21__16_, CARRYB_21__15_,
         CARRYB_21__14_, CARRYB_21__13_, CARRYB_21__12_, CARRYB_21__11_,
         CARRYB_21__10_, CARRYB_21__9_, CARRYB_21__8_, CARRYB_21__7_,
         CARRYB_21__6_, CARRYB_21__5_, CARRYB_21__4_, CARRYB_21__3_,
         CARRYB_21__2_, CARRYB_21__1_, CARRYB_21__0_, CARRYB_20__22_,
         CARRYB_20__21_, CARRYB_20__20_, CARRYB_20__19_, CARRYB_20__18_,
         CARRYB_20__17_, CARRYB_20__16_, CARRYB_20__15_, CARRYB_20__14_,
         CARRYB_20__13_, CARRYB_20__12_, CARRYB_20__11_, CARRYB_20__10_,
         CARRYB_20__9_, CARRYB_20__8_, CARRYB_20__7_, CARRYB_20__6_,
         CARRYB_20__5_, CARRYB_20__4_, CARRYB_20__3_, CARRYB_20__2_,
         CARRYB_20__1_, CARRYB_20__0_, CARRYB_19__22_, CARRYB_19__21_,
         CARRYB_19__20_, CARRYB_19__19_, CARRYB_19__18_, CARRYB_19__17_,
         CARRYB_19__16_, CARRYB_19__15_, CARRYB_19__14_, CARRYB_19__13_,
         CARRYB_19__12_, CARRYB_19__11_, CARRYB_19__10_, CARRYB_19__9_,
         CARRYB_19__8_, CARRYB_19__7_, CARRYB_19__6_, CARRYB_19__5_,
         CARRYB_19__4_, CARRYB_19__3_, CARRYB_19__2_, CARRYB_19__1_,
         CARRYB_19__0_, CARRYB_18__22_, CARRYB_18__21_, CARRYB_18__20_,
         CARRYB_18__19_, CARRYB_18__18_, CARRYB_18__17_, CARRYB_18__16_,
         CARRYB_18__15_, CARRYB_18__14_, CARRYB_18__13_, CARRYB_18__12_,
         CARRYB_18__11_, CARRYB_18__10_, CARRYB_18__9_, CARRYB_18__8_,
         CARRYB_18__7_, CARRYB_18__6_, CARRYB_18__5_, CARRYB_18__4_,
         CARRYB_18__3_, CARRYB_18__2_, CARRYB_18__1_, CARRYB_18__0_,
         CARRYB_17__22_, CARRYB_17__21_, CARRYB_17__20_, CARRYB_17__19_,
         CARRYB_17__18_, CARRYB_17__17_, CARRYB_17__16_, CARRYB_17__15_,
         CARRYB_17__14_, CARRYB_17__13_, CARRYB_17__12_, CARRYB_17__11_,
         CARRYB_17__10_, CARRYB_17__9_, CARRYB_17__8_, CARRYB_17__7_,
         CARRYB_17__6_, CARRYB_17__5_, CARRYB_17__4_, CARRYB_17__3_,
         CARRYB_17__2_, CARRYB_17__1_, CARRYB_17__0_, CARRYB_16__22_,
         CARRYB_16__21_, CARRYB_16__20_, CARRYB_16__19_, CARRYB_16__18_,
         CARRYB_16__17_, CARRYB_16__16_, CARRYB_16__15_, CARRYB_16__14_,
         CARRYB_16__13_, CARRYB_16__12_, CARRYB_16__11_, CARRYB_16__10_,
         CARRYB_16__9_, CARRYB_16__8_, CARRYB_16__7_, CARRYB_16__6_,
         CARRYB_16__5_, CARRYB_16__4_, CARRYB_16__3_, CARRYB_16__2_,
         CARRYB_16__1_, CARRYB_16__0_, CARRYB_15__22_, CARRYB_15__21_,
         CARRYB_15__20_, CARRYB_15__19_, CARRYB_15__18_, CARRYB_15__17_,
         CARRYB_15__16_, CARRYB_15__15_, CARRYB_15__14_, CARRYB_15__13_,
         CARRYB_15__12_, CARRYB_15__11_, CARRYB_15__10_, CARRYB_15__9_,
         CARRYB_15__8_, CARRYB_15__7_, CARRYB_15__6_, CARRYB_15__5_,
         CARRYB_15__4_, CARRYB_15__3_, CARRYB_15__2_, CARRYB_15__1_,
         CARRYB_15__0_, CARRYB_14__22_, CARRYB_14__21_, CARRYB_14__20_,
         CARRYB_14__19_, CARRYB_14__18_, CARRYB_14__17_, CARRYB_14__16_,
         CARRYB_14__15_, CARRYB_14__14_, CARRYB_14__13_, CARRYB_14__12_,
         CARRYB_14__11_, CARRYB_14__10_, CARRYB_14__9_, CARRYB_14__8_,
         CARRYB_14__7_, CARRYB_14__6_, CARRYB_14__5_, CARRYB_14__4_,
         CARRYB_14__3_, CARRYB_14__2_, CARRYB_14__1_, CARRYB_14__0_,
         CARRYB_13__22_, CARRYB_13__21_, CARRYB_13__20_, CARRYB_13__19_,
         CARRYB_13__18_, CARRYB_13__17_, CARRYB_13__16_, CARRYB_13__15_,
         CARRYB_13__14_, CARRYB_13__13_, CARRYB_13__12_, CARRYB_13__11_,
         CARRYB_13__10_, CARRYB_13__9_, CARRYB_13__8_, CARRYB_13__7_,
         CARRYB_13__6_, CARRYB_13__5_, CARRYB_13__4_, CARRYB_13__3_,
         CARRYB_13__2_, CARRYB_13__1_, CARRYB_13__0_, CARRYB_12__22_,
         CARRYB_12__21_, CARRYB_12__20_, CARRYB_12__19_, CARRYB_12__18_,
         CARRYB_12__17_, CARRYB_12__16_, CARRYB_12__15_, CARRYB_12__14_,
         CARRYB_12__13_, CARRYB_12__12_, CARRYB_12__11_, CARRYB_12__10_,
         CARRYB_12__9_, CARRYB_12__8_, CARRYB_12__7_, CARRYB_12__6_,
         CARRYB_12__5_, CARRYB_12__4_, CARRYB_12__3_, CARRYB_12__2_,
         CARRYB_12__1_, CARRYB_12__0_, CARRYB_11__22_, CARRYB_11__21_,
         CARRYB_11__20_, CARRYB_11__19_, CARRYB_11__18_, CARRYB_11__17_,
         CARRYB_11__16_, CARRYB_11__15_, CARRYB_11__14_, CARRYB_11__13_,
         CARRYB_11__12_, CARRYB_11__11_, CARRYB_11__10_, CARRYB_11__9_,
         CARRYB_11__8_, CARRYB_11__7_, CARRYB_11__6_, CARRYB_11__5_,
         CARRYB_11__4_, CARRYB_11__3_, CARRYB_11__2_, CARRYB_11__1_,
         CARRYB_11__0_, CARRYB_10__22_, CARRYB_10__21_, CARRYB_10__20_,
         CARRYB_10__19_, CARRYB_10__18_, CARRYB_10__17_, CARRYB_10__16_,
         CARRYB_10__15_, CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_,
         CARRYB_10__11_, CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_,
         CARRYB_10__7_, CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_,
         CARRYB_10__3_, CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_,
         CARRYB_9__22_, CARRYB_9__21_, CARRYB_9__20_, CARRYB_9__19_,
         CARRYB_9__18_, CARRYB_9__17_, CARRYB_9__16_, CARRYB_9__15_,
         CARRYB_9__14_, CARRYB_9__13_, CARRYB_9__12_, CARRYB_9__11_,
         CARRYB_9__10_, CARRYB_9__9_, CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_,
         CARRYB_9__5_, CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_,
         CARRYB_9__0_, CARRYB_8__22_, CARRYB_8__21_, CARRYB_8__20_,
         CARRYB_8__19_, CARRYB_8__18_, CARRYB_8__17_, CARRYB_8__16_,
         CARRYB_8__15_, CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_,
         CARRYB_8__11_, CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_,
         CARRYB_8__7_, CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_,
         CARRYB_8__2_, CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__22_,
         CARRYB_7__21_, CARRYB_7__20_, CARRYB_7__19_, CARRYB_7__18_,
         CARRYB_7__17_, CARRYB_7__16_, CARRYB_7__15_, CARRYB_7__14_,
         CARRYB_7__13_, CARRYB_7__12_, CARRYB_7__11_, CARRYB_7__10_,
         CARRYB_7__9_, CARRYB_7__8_, CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_,
         CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_,
         CARRYB_6__22_, CARRYB_6__21_, CARRYB_6__20_, CARRYB_6__19_,
         CARRYB_6__18_, CARRYB_6__17_, CARRYB_6__16_, CARRYB_6__15_,
         CARRYB_6__14_, CARRYB_6__13_, CARRYB_6__12_, CARRYB_6__11_,
         CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_, CARRYB_6__7_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__22_, CARRYB_5__21_, CARRYB_5__20_,
         CARRYB_5__19_, CARRYB_5__18_, CARRYB_5__17_, CARRYB_5__16_,
         CARRYB_5__15_, CARRYB_5__14_, CARRYB_5__13_, CARRYB_5__12_,
         CARRYB_5__11_, CARRYB_5__10_, CARRYB_5__9_, CARRYB_5__8_,
         CARRYB_5__7_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__22_,
         CARRYB_4__21_, CARRYB_4__20_, CARRYB_4__19_, CARRYB_4__18_,
         CARRYB_4__17_, CARRYB_4__16_, CARRYB_4__15_, CARRYB_4__14_,
         CARRYB_4__13_, CARRYB_4__12_, CARRYB_4__11_, CARRYB_4__10_,
         CARRYB_4__9_, CARRYB_4__8_, CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__22_, CARRYB_3__21_, CARRYB_3__20_, CARRYB_3__19_,
         CARRYB_3__18_, CARRYB_3__17_, CARRYB_3__16_, CARRYB_3__15_,
         CARRYB_3__14_, CARRYB_3__13_, CARRYB_3__12_, CARRYB_3__11_,
         CARRYB_3__10_, CARRYB_3__9_, CARRYB_3__8_, CARRYB_3__7_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__22_, CARRYB_2__21_, CARRYB_2__20_,
         CARRYB_2__19_, CARRYB_2__18_, CARRYB_2__17_, CARRYB_2__16_,
         CARRYB_2__15_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__22_,
         CARRYB_1__21_, CARRYB_1__20_, CARRYB_1__19_, CARRYB_1__18_,
         CARRYB_1__17_, CARRYB_1__16_, CARRYB_1__15_, CARRYB_1__14_,
         CARRYB_1__13_, CARRYB_1__12_, CARRYB_1__11_, CARRYB_1__10_,
         CARRYB_1__9_, CARRYB_1__8_, CARRYB_1__7_, CARRYB_1__6_, CARRYB_1__5_,
         CARRYB_1__4_, CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_,
         SUMB_23__23_, SUMB_23__22_, SUMB_23__21_, SUMB_23__20_, SUMB_23__19_,
         SUMB_23__18_, SUMB_23__17_, SUMB_23__16_, SUMB_23__15_, SUMB_23__14_,
         SUMB_23__13_, SUMB_23__12_, SUMB_23__11_, SUMB_23__10_, SUMB_23__9_,
         SUMB_23__8_, SUMB_23__7_, SUMB_23__6_, SUMB_23__5_, SUMB_23__4_,
         SUMB_23__3_, SUMB_23__2_, SUMB_23__1_, SUMB_23__0_, SUMB_22__22_,
         SUMB_22__21_, SUMB_22__20_, SUMB_22__19_, SUMB_22__18_, SUMB_22__17_,
         SUMB_22__16_, SUMB_22__15_, SUMB_22__14_, SUMB_22__13_, SUMB_22__12_,
         SUMB_22__11_, SUMB_22__10_, SUMB_22__9_, SUMB_22__8_, SUMB_22__7_,
         SUMB_22__6_, SUMB_22__5_, SUMB_22__4_, SUMB_22__3_, SUMB_22__2_,
         SUMB_22__1_, SUMB_21__22_, SUMB_21__21_, SUMB_21__20_, SUMB_21__19_,
         SUMB_21__18_, SUMB_21__17_, SUMB_21__16_, SUMB_21__15_, SUMB_21__14_,
         SUMB_21__13_, SUMB_21__12_, SUMB_21__11_, SUMB_21__10_, SUMB_21__9_,
         SUMB_21__8_, SUMB_21__7_, SUMB_21__6_, SUMB_21__5_, SUMB_21__4_,
         SUMB_21__3_, SUMB_21__2_, SUMB_21__1_, SUMB_20__22_, SUMB_20__21_,
         SUMB_20__20_, SUMB_20__19_, SUMB_20__18_, SUMB_20__17_, SUMB_20__16_,
         SUMB_20__15_, SUMB_20__14_, SUMB_20__13_, SUMB_20__12_, SUMB_20__11_,
         SUMB_20__10_, SUMB_20__9_, SUMB_20__8_, SUMB_20__7_, SUMB_20__6_,
         SUMB_20__5_, SUMB_20__4_, SUMB_20__3_, SUMB_20__2_, SUMB_20__1_,
         SUMB_19__22_, SUMB_19__21_, SUMB_19__20_, SUMB_19__19_, SUMB_19__18_,
         SUMB_19__17_, SUMB_19__16_, SUMB_19__15_, SUMB_19__14_, SUMB_19__13_,
         SUMB_19__12_, SUMB_19__11_, SUMB_19__10_, SUMB_19__9_, SUMB_19__8_,
         SUMB_19__7_, SUMB_19__6_, SUMB_19__5_, SUMB_19__4_, SUMB_19__3_,
         SUMB_19__2_, SUMB_19__1_, SUMB_18__22_, SUMB_18__21_, SUMB_18__20_,
         SUMB_18__19_, SUMB_18__18_, SUMB_18__17_, SUMB_18__16_, SUMB_18__15_,
         SUMB_18__14_, SUMB_18__13_, SUMB_18__12_, SUMB_18__11_, SUMB_18__10_,
         SUMB_18__9_, SUMB_18__8_, SUMB_18__7_, SUMB_18__6_, SUMB_18__5_,
         SUMB_18__4_, SUMB_18__3_, SUMB_18__2_, SUMB_18__1_, SUMB_17__22_,
         SUMB_17__21_, SUMB_17__20_, SUMB_17__19_, SUMB_17__18_, SUMB_17__17_,
         SUMB_17__16_, SUMB_17__15_, SUMB_17__14_, SUMB_17__13_, SUMB_17__12_,
         SUMB_17__11_, SUMB_17__10_, SUMB_17__9_, SUMB_17__8_, SUMB_17__7_,
         SUMB_17__6_, SUMB_17__5_, SUMB_17__4_, SUMB_17__3_, SUMB_17__2_,
         SUMB_17__1_, SUMB_16__22_, SUMB_16__21_, SUMB_16__20_, SUMB_16__19_,
         SUMB_16__18_, SUMB_16__17_, SUMB_16__16_, SUMB_16__15_, SUMB_16__14_,
         SUMB_16__13_, SUMB_16__12_, SUMB_16__11_, SUMB_16__10_, SUMB_16__9_,
         SUMB_16__8_, SUMB_16__7_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_,
         SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, SUMB_15__22_, SUMB_15__21_,
         SUMB_15__20_, SUMB_15__19_, SUMB_15__18_, SUMB_15__17_, SUMB_15__16_,
         SUMB_15__15_, SUMB_15__14_, SUMB_15__13_, SUMB_15__12_, SUMB_15__11_,
         SUMB_15__10_, SUMB_15__9_, SUMB_15__8_, SUMB_15__7_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_14__22_, SUMB_14__21_, SUMB_14__20_, SUMB_14__19_, SUMB_14__18_,
         SUMB_14__17_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_, SUMB_14__13_,
         SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_, SUMB_14__8_,
         SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_,
         SUMB_14__2_, SUMB_14__1_, SUMB_13__22_, SUMB_13__21_, SUMB_13__20_,
         SUMB_13__19_, SUMB_13__18_, SUMB_13__17_, SUMB_13__16_, SUMB_13__15_,
         SUMB_13__14_, SUMB_13__13_, SUMB_13__12_, SUMB_13__11_, SUMB_13__10_,
         SUMB_13__9_, SUMB_13__8_, SUMB_13__7_, SUMB_13__6_, SUMB_13__5_,
         SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_, SUMB_12__22_,
         SUMB_12__21_, SUMB_12__20_, SUMB_12__19_, SUMB_12__18_, SUMB_12__17_,
         SUMB_12__16_, SUMB_12__15_, SUMB_12__14_, SUMB_12__13_, SUMB_12__12_,
         SUMB_12__11_, SUMB_12__10_, SUMB_12__9_, SUMB_12__8_, SUMB_12__7_,
         SUMB_12__6_, SUMB_12__5_, SUMB_12__4_, SUMB_12__3_, SUMB_12__2_,
         SUMB_12__1_, SUMB_11__22_, SUMB_11__21_, SUMB_11__20_, SUMB_11__19_,
         SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_, SUMB_11__14_,
         SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_, SUMB_11__9_,
         SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_, SUMB_11__4_,
         SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__22_, SUMB_10__21_,
         SUMB_10__20_, SUMB_10__19_, SUMB_10__18_, SUMB_10__17_, SUMB_10__16_,
         SUMB_10__15_, SUMB_10__14_, SUMB_10__13_, SUMB_10__12_, SUMB_10__11_,
         SUMB_10__10_, SUMB_10__9_, SUMB_10__8_, SUMB_10__7_, SUMB_10__6_,
         SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_,
         SUMB_9__22_, SUMB_9__21_, SUMB_9__20_, SUMB_9__19_, SUMB_9__18_,
         SUMB_9__17_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_, SUMB_9__13_,
         SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_, SUMB_9__8_,
         SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_,
         SUMB_9__2_, SUMB_9__1_, SUMB_8__22_, SUMB_8__21_, SUMB_8__20_,
         SUMB_8__19_, SUMB_8__18_, SUMB_8__17_, SUMB_8__16_, SUMB_8__15_,
         SUMB_8__14_, SUMB_8__13_, SUMB_8__12_, SUMB_8__11_, SUMB_8__10_,
         SUMB_8__9_, SUMB_8__8_, SUMB_8__7_, SUMB_8__6_, SUMB_8__5_,
         SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_, SUMB_7__22_,
         SUMB_7__21_, SUMB_7__20_, SUMB_7__19_, SUMB_7__18_, SUMB_7__17_,
         SUMB_7__16_, SUMB_7__15_, SUMB_7__14_, SUMB_7__13_, SUMB_7__12_,
         SUMB_7__11_, SUMB_7__10_, SUMB_7__9_, SUMB_7__8_, SUMB_7__7_,
         SUMB_7__6_, SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_,
         SUMB_7__1_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_, SUMB_6__19_,
         SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_, SUMB_6__14_,
         SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_, SUMB_6__9_,
         SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_,
         SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__22_, SUMB_5__21_,
         SUMB_5__20_, SUMB_5__19_, SUMB_5__18_, SUMB_5__17_, SUMB_5__16_,
         SUMB_5__15_, SUMB_5__14_, SUMB_5__13_, SUMB_5__12_, SUMB_5__11_,
         SUMB_5__10_, SUMB_5__9_, SUMB_5__8_, SUMB_5__7_, SUMB_5__6_,
         SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_,
         SUMB_4__22_, SUMB_4__21_, SUMB_4__20_, SUMB_4__19_, SUMB_4__18_,
         SUMB_4__17_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_, SUMB_4__13_,
         SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_, SUMB_4__8_,
         SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_,
         SUMB_4__2_, SUMB_4__1_, SUMB_3__22_, SUMB_3__21_, SUMB_3__20_,
         SUMB_3__19_, SUMB_3__18_, SUMB_3__17_, SUMB_3__16_, SUMB_3__15_,
         SUMB_3__14_, SUMB_3__13_, SUMB_3__12_, SUMB_3__11_, SUMB_3__10_,
         SUMB_3__9_, SUMB_3__8_, SUMB_3__7_, SUMB_3__6_, SUMB_3__5_,
         SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_, SUMB_2__22_,
         SUMB_2__21_, SUMB_2__20_, SUMB_2__19_, SUMB_2__18_, SUMB_2__17_,
         SUMB_2__16_, SUMB_2__15_, SUMB_2__14_, SUMB_2__13_, SUMB_2__12_,
         SUMB_2__11_, SUMB_2__10_, SUMB_2__9_, SUMB_2__8_, SUMB_2__7_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__22_, SUMB_1__21_, SUMB_1__20_, SUMB_1__19_,
         SUMB_1__18_, SUMB_1__17_, SUMB_1__16_, SUMB_1__15_, SUMB_1__14_,
         SUMB_1__13_, SUMB_1__12_, SUMB_1__11_, SUMB_1__10_, SUMB_1__9_,
         SUMB_1__8_, SUMB_1__7_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_,
         SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, QA, QB, A1_45_, A1_44_, A1_43_,
         A1_42_, A1_41_, A1_40_, A1_39_, A1_38_, A1_37_, A1_36_, A1_35_,
         A1_34_, A1_33_, A1_32_, A1_31_, A1_30_, A1_29_, A1_28_, A1_27_,
         A1_26_, A1_25_, A1_24_, A1_23_, A1_22_, A1_21_, A1_20_, A1_19_,
         A1_18_, A1_17_, A1_16_, A1_15_, A1_14_, A1_13_, A1_12_, A1_11_,
         A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_,
         A1_0_, A2_45_, A2_44_, A2_43_, A2_42_, A2_41_, A2_40_, A2_39_, A2_38_,
         A2_37_, A2_36_, A2_35_, A2_34_, A2_33_, A2_32_, A2_31_, A2_30_,
         A2_29_, A2_28_, A2_27_, A2_26_, A2_25_, A2_24_, A2_23_, A2_22_, n1,
         n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21;

  FA_X1 S14_23_0 ( .A(A[23]), .B(B[23]), .CI(SUMB_23__0_), .CO(A2_22_), .S(
        A1_21_) );
  FA_X1 S4_0 ( .A(ab_23__0_), .B(CARRYB_22__0_), .CI(SUMB_22__1_), .CO(
        CARRYB_23__0_), .S(SUMB_23__0_) );
  FA_X1 S4_1 ( .A(ab_23__1_), .B(CARRYB_22__1_), .CI(SUMB_22__2_), .CO(
        CARRYB_23__1_), .S(SUMB_23__1_) );
  FA_X1 S4_2 ( .A(ab_23__2_), .B(CARRYB_22__2_), .CI(SUMB_22__3_), .CO(
        CARRYB_23__2_), .S(SUMB_23__2_) );
  FA_X1 S4_3 ( .A(ab_23__3_), .B(CARRYB_22__3_), .CI(SUMB_22__4_), .CO(
        CARRYB_23__3_), .S(SUMB_23__3_) );
  FA_X1 S4_4 ( .A(ab_23__4_), .B(CARRYB_22__4_), .CI(SUMB_22__5_), .CO(
        CARRYB_23__4_), .S(SUMB_23__4_) );
  FA_X1 S4_5 ( .A(ab_23__5_), .B(CARRYB_22__5_), .CI(SUMB_22__6_), .CO(
        CARRYB_23__5_), .S(SUMB_23__5_) );
  FA_X1 S4_6 ( .A(ab_23__6_), .B(CARRYB_22__6_), .CI(SUMB_22__7_), .CO(
        CARRYB_23__6_), .S(SUMB_23__6_) );
  FA_X1 S4_7 ( .A(ab_23__7_), .B(CARRYB_22__7_), .CI(SUMB_22__8_), .CO(
        CARRYB_23__7_), .S(SUMB_23__7_) );
  FA_X1 S4_8 ( .A(ab_23__8_), .B(CARRYB_22__8_), .CI(SUMB_22__9_), .CO(
        CARRYB_23__8_), .S(SUMB_23__8_) );
  FA_X1 S4_9 ( .A(ab_23__9_), .B(CARRYB_22__9_), .CI(SUMB_22__10_), .CO(
        CARRYB_23__9_), .S(SUMB_23__9_) );
  FA_X1 S4_10 ( .A(ab_23__10_), .B(CARRYB_22__10_), .CI(SUMB_22__11_), .CO(
        CARRYB_23__10_), .S(SUMB_23__10_) );
  FA_X1 S4_11 ( .A(ab_23__11_), .B(CARRYB_22__11_), .CI(SUMB_22__12_), .CO(
        CARRYB_23__11_), .S(SUMB_23__11_) );
  FA_X1 S4_12 ( .A(ab_23__12_), .B(CARRYB_22__12_), .CI(SUMB_22__13_), .CO(
        CARRYB_23__12_), .S(SUMB_23__12_) );
  FA_X1 S4_13 ( .A(ab_23__13_), .B(CARRYB_22__13_), .CI(SUMB_22__14_), .CO(
        CARRYB_23__13_), .S(SUMB_23__13_) );
  FA_X1 S4_14 ( .A(ab_23__14_), .B(CARRYB_22__14_), .CI(SUMB_22__15_), .CO(
        CARRYB_23__14_), .S(SUMB_23__14_) );
  FA_X1 S4_15 ( .A(ab_23__15_), .B(CARRYB_22__15_), .CI(SUMB_22__16_), .CO(
        CARRYB_23__15_), .S(SUMB_23__15_) );
  FA_X1 S4_16 ( .A(ab_23__16_), .B(CARRYB_22__16_), .CI(SUMB_22__17_), .CO(
        CARRYB_23__16_), .S(SUMB_23__16_) );
  FA_X1 S4_17 ( .A(ab_23__17_), .B(CARRYB_22__17_), .CI(SUMB_22__18_), .CO(
        CARRYB_23__17_), .S(SUMB_23__17_) );
  FA_X1 S4_18 ( .A(ab_23__18_), .B(CARRYB_22__18_), .CI(SUMB_22__19_), .CO(
        CARRYB_23__18_), .S(SUMB_23__18_) );
  FA_X1 S4_19 ( .A(ab_23__19_), .B(CARRYB_22__19_), .CI(SUMB_22__20_), .CO(
        CARRYB_23__19_), .S(SUMB_23__19_) );
  FA_X1 S4_20 ( .A(ab_23__20_), .B(CARRYB_22__20_), .CI(SUMB_22__21_), .CO(
        CARRYB_23__20_), .S(SUMB_23__20_) );
  FA_X1 S4_21 ( .A(ab_23__21_), .B(CARRYB_22__21_), .CI(SUMB_22__22_), .CO(
        CARRYB_23__21_), .S(SUMB_23__21_) );
  FA_X1 S5_22 ( .A(ab_23__22_), .B(CARRYB_22__22_), .CI(ab_22__23_), .CO(
        CARRYB_23__22_), .S(SUMB_23__22_) );
  FA_X1 S14_23 ( .A(n3), .B(n1), .CI(ab_23__23_), .CO(CARRYB_23__23_), .S(
        SUMB_23__23_) );
  FA_X1 S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), .CO(
        CARRYB_22__0_), .S(A1_20_) );
  FA_X1 S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), .CO(
        CARRYB_22__1_), .S(SUMB_22__1_) );
  FA_X1 S2_22_2 ( .A(ab_22__2_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), .CO(
        CARRYB_22__2_), .S(SUMB_22__2_) );
  FA_X1 S2_22_3 ( .A(ab_22__3_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), .CO(
        CARRYB_22__3_), .S(SUMB_22__3_) );
  FA_X1 S2_22_4 ( .A(ab_22__4_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), .CO(
        CARRYB_22__4_), .S(SUMB_22__4_) );
  FA_X1 S2_22_5 ( .A(ab_22__5_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), .CO(
        CARRYB_22__5_), .S(SUMB_22__5_) );
  FA_X1 S2_22_6 ( .A(ab_22__6_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), .CO(
        CARRYB_22__6_), .S(SUMB_22__6_) );
  FA_X1 S2_22_7 ( .A(ab_22__7_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), .CO(
        CARRYB_22__7_), .S(SUMB_22__7_) );
  FA_X1 S2_22_8 ( .A(ab_22__8_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), .CO(
        CARRYB_22__8_), .S(SUMB_22__8_) );
  FA_X1 S2_22_9 ( .A(ab_22__9_), .B(CARRYB_21__9_), .CI(SUMB_21__10_), .CO(
        CARRYB_22__9_), .S(SUMB_22__9_) );
  FA_X1 S2_22_10 ( .A(ab_22__10_), .B(CARRYB_21__10_), .CI(SUMB_21__11_), .CO(
        CARRYB_22__10_), .S(SUMB_22__10_) );
  FA_X1 S2_22_11 ( .A(ab_22__11_), .B(CARRYB_21__11_), .CI(SUMB_21__12_), .CO(
        CARRYB_22__11_), .S(SUMB_22__11_) );
  FA_X1 S2_22_12 ( .A(ab_22__12_), .B(CARRYB_21__12_), .CI(SUMB_21__13_), .CO(
        CARRYB_22__12_), .S(SUMB_22__12_) );
  FA_X1 S2_22_13 ( .A(ab_22__13_), .B(CARRYB_21__13_), .CI(SUMB_21__14_), .CO(
        CARRYB_22__13_), .S(SUMB_22__13_) );
  FA_X1 S2_22_14 ( .A(ab_22__14_), .B(CARRYB_21__14_), .CI(SUMB_21__15_), .CO(
        CARRYB_22__14_), .S(SUMB_22__14_) );
  FA_X1 S2_22_15 ( .A(ab_22__15_), .B(CARRYB_21__15_), .CI(SUMB_21__16_), .CO(
        CARRYB_22__15_), .S(SUMB_22__15_) );
  FA_X1 S2_22_16 ( .A(ab_22__16_), .B(CARRYB_21__16_), .CI(SUMB_21__17_), .CO(
        CARRYB_22__16_), .S(SUMB_22__16_) );
  FA_X1 S2_22_17 ( .A(ab_22__17_), .B(CARRYB_21__17_), .CI(SUMB_21__18_), .CO(
        CARRYB_22__17_), .S(SUMB_22__17_) );
  FA_X1 S2_22_18 ( .A(ab_22__18_), .B(CARRYB_21__18_), .CI(SUMB_21__19_), .CO(
        CARRYB_22__18_), .S(SUMB_22__18_) );
  FA_X1 S2_22_19 ( .A(ab_22__19_), .B(CARRYB_21__19_), .CI(SUMB_21__20_), .CO(
        CARRYB_22__19_), .S(SUMB_22__19_) );
  FA_X1 S2_22_20 ( .A(ab_22__20_), .B(CARRYB_21__20_), .CI(SUMB_21__21_), .CO(
        CARRYB_22__20_), .S(SUMB_22__20_) );
  FA_X1 S2_22_21 ( .A(ab_22__21_), .B(CARRYB_21__21_), .CI(SUMB_21__22_), .CO(
        CARRYB_22__21_), .S(SUMB_22__21_) );
  FA_X1 S3_22_22 ( .A(ab_22__22_), .B(CARRYB_21__22_), .CI(ab_21__23_), .CO(
        CARRYB_22__22_), .S(SUMB_22__22_) );
  FA_X1 S1_21_0 ( .A(ab_21__0_), .B(CARRYB_20__0_), .CI(SUMB_20__1_), .CO(
        CARRYB_21__0_), .S(A1_19_) );
  FA_X1 S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), .CO(
        CARRYB_21__1_), .S(SUMB_21__1_) );
  FA_X1 S2_21_2 ( .A(ab_21__2_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), .CO(
        CARRYB_21__2_), .S(SUMB_21__2_) );
  FA_X1 S2_21_3 ( .A(ab_21__3_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), .CO(
        CARRYB_21__3_), .S(SUMB_21__3_) );
  FA_X1 S2_21_4 ( .A(ab_21__4_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), .CO(
        CARRYB_21__4_), .S(SUMB_21__4_) );
  FA_X1 S2_21_5 ( .A(ab_21__5_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), .CO(
        CARRYB_21__5_), .S(SUMB_21__5_) );
  FA_X1 S2_21_6 ( .A(ab_21__6_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), .CO(
        CARRYB_21__6_), .S(SUMB_21__6_) );
  FA_X1 S2_21_7 ( .A(ab_21__7_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), .CO(
        CARRYB_21__7_), .S(SUMB_21__7_) );
  FA_X1 S2_21_8 ( .A(ab_21__8_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), .CO(
        CARRYB_21__8_), .S(SUMB_21__8_) );
  FA_X1 S2_21_9 ( .A(ab_21__9_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), .CO(
        CARRYB_21__9_), .S(SUMB_21__9_) );
  FA_X1 S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .CI(SUMB_20__11_), .CO(
        CARRYB_21__10_), .S(SUMB_21__10_) );
  FA_X1 S2_21_11 ( .A(ab_21__11_), .B(CARRYB_20__11_), .CI(SUMB_20__12_), .CO(
        CARRYB_21__11_), .S(SUMB_21__11_) );
  FA_X1 S2_21_12 ( .A(ab_21__12_), .B(CARRYB_20__12_), .CI(SUMB_20__13_), .CO(
        CARRYB_21__12_), .S(SUMB_21__12_) );
  FA_X1 S2_21_13 ( .A(ab_21__13_), .B(CARRYB_20__13_), .CI(SUMB_20__14_), .CO(
        CARRYB_21__13_), .S(SUMB_21__13_) );
  FA_X1 S2_21_14 ( .A(ab_21__14_), .B(CARRYB_20__14_), .CI(SUMB_20__15_), .CO(
        CARRYB_21__14_), .S(SUMB_21__14_) );
  FA_X1 S2_21_15 ( .A(ab_21__15_), .B(CARRYB_20__15_), .CI(SUMB_20__16_), .CO(
        CARRYB_21__15_), .S(SUMB_21__15_) );
  FA_X1 S2_21_16 ( .A(ab_21__16_), .B(CARRYB_20__16_), .CI(SUMB_20__17_), .CO(
        CARRYB_21__16_), .S(SUMB_21__16_) );
  FA_X1 S2_21_17 ( .A(ab_21__17_), .B(CARRYB_20__17_), .CI(SUMB_20__18_), .CO(
        CARRYB_21__17_), .S(SUMB_21__17_) );
  FA_X1 S2_21_18 ( .A(ab_21__18_), .B(CARRYB_20__18_), .CI(SUMB_20__19_), .CO(
        CARRYB_21__18_), .S(SUMB_21__18_) );
  FA_X1 S2_21_19 ( .A(ab_21__19_), .B(CARRYB_20__19_), .CI(SUMB_20__20_), .CO(
        CARRYB_21__19_), .S(SUMB_21__19_) );
  FA_X1 S2_21_20 ( .A(ab_21__20_), .B(CARRYB_20__20_), .CI(SUMB_20__21_), .CO(
        CARRYB_21__20_), .S(SUMB_21__20_) );
  FA_X1 S2_21_21 ( .A(ab_21__21_), .B(CARRYB_20__21_), .CI(SUMB_20__22_), .CO(
        CARRYB_21__21_), .S(SUMB_21__21_) );
  FA_X1 S3_21_22 ( .A(ab_21__22_), .B(CARRYB_20__22_), .CI(ab_20__23_), .CO(
        CARRYB_21__22_), .S(SUMB_21__22_) );
  FA_X1 S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), .CO(
        CARRYB_20__0_), .S(A1_18_) );
  FA_X1 S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), .CO(
        CARRYB_20__1_), .S(SUMB_20__1_) );
  FA_X1 S2_20_2 ( .A(ab_20__2_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), .CO(
        CARRYB_20__2_), .S(SUMB_20__2_) );
  FA_X1 S2_20_3 ( .A(ab_20__3_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), .CO(
        CARRYB_20__3_), .S(SUMB_20__3_) );
  FA_X1 S2_20_4 ( .A(ab_20__4_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), .CO(
        CARRYB_20__4_), .S(SUMB_20__4_) );
  FA_X1 S2_20_5 ( .A(ab_20__5_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), .CO(
        CARRYB_20__5_), .S(SUMB_20__5_) );
  FA_X1 S2_20_6 ( .A(ab_20__6_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), .CO(
        CARRYB_20__6_), .S(SUMB_20__6_) );
  FA_X1 S2_20_7 ( .A(ab_20__7_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), .CO(
        CARRYB_20__7_), .S(SUMB_20__7_) );
  FA_X1 S2_20_8 ( .A(ab_20__8_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), .CO(
        CARRYB_20__8_), .S(SUMB_20__8_) );
  FA_X1 S2_20_9 ( .A(ab_20__9_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), .CO(
        CARRYB_20__9_), .S(SUMB_20__9_) );
  FA_X1 S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), .CO(
        CARRYB_20__10_), .S(SUMB_20__10_) );
  FA_X1 S2_20_11 ( .A(ab_20__11_), .B(CARRYB_19__11_), .CI(SUMB_19__12_), .CO(
        CARRYB_20__11_), .S(SUMB_20__11_) );
  FA_X1 S2_20_12 ( .A(ab_20__12_), .B(CARRYB_19__12_), .CI(SUMB_19__13_), .CO(
        CARRYB_20__12_), .S(SUMB_20__12_) );
  FA_X1 S2_20_13 ( .A(ab_20__13_), .B(CARRYB_19__13_), .CI(SUMB_19__14_), .CO(
        CARRYB_20__13_), .S(SUMB_20__13_) );
  FA_X1 S2_20_14 ( .A(ab_20__14_), .B(CARRYB_19__14_), .CI(SUMB_19__15_), .CO(
        CARRYB_20__14_), .S(SUMB_20__14_) );
  FA_X1 S2_20_15 ( .A(ab_20__15_), .B(CARRYB_19__15_), .CI(SUMB_19__16_), .CO(
        CARRYB_20__15_), .S(SUMB_20__15_) );
  FA_X1 S2_20_16 ( .A(ab_20__16_), .B(CARRYB_19__16_), .CI(SUMB_19__17_), .CO(
        CARRYB_20__16_), .S(SUMB_20__16_) );
  FA_X1 S2_20_17 ( .A(ab_20__17_), .B(CARRYB_19__17_), .CI(SUMB_19__18_), .CO(
        CARRYB_20__17_), .S(SUMB_20__17_) );
  FA_X1 S2_20_18 ( .A(ab_20__18_), .B(CARRYB_19__18_), .CI(SUMB_19__19_), .CO(
        CARRYB_20__18_), .S(SUMB_20__18_) );
  FA_X1 S2_20_19 ( .A(ab_20__19_), .B(CARRYB_19__19_), .CI(SUMB_19__20_), .CO(
        CARRYB_20__19_), .S(SUMB_20__19_) );
  FA_X1 S2_20_20 ( .A(ab_20__20_), .B(CARRYB_19__20_), .CI(SUMB_19__21_), .CO(
        CARRYB_20__20_), .S(SUMB_20__20_) );
  FA_X1 S2_20_21 ( .A(ab_20__21_), .B(CARRYB_19__21_), .CI(SUMB_19__22_), .CO(
        CARRYB_20__21_), .S(SUMB_20__21_) );
  FA_X1 S3_20_22 ( .A(ab_20__22_), .B(CARRYB_19__22_), .CI(ab_19__23_), .CO(
        CARRYB_20__22_), .S(SUMB_20__22_) );
  FA_X1 S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), .CO(
        CARRYB_19__0_), .S(A1_17_) );
  FA_X1 S2_19_1 ( .A(ab_19__1_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), .CO(
        CARRYB_19__1_), .S(SUMB_19__1_) );
  FA_X1 S2_19_2 ( .A(ab_19__2_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), .CO(
        CARRYB_19__2_), .S(SUMB_19__2_) );
  FA_X1 S2_19_3 ( .A(ab_19__3_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), .CO(
        CARRYB_19__3_), .S(SUMB_19__3_) );
  FA_X1 S2_19_4 ( .A(ab_19__4_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), .CO(
        CARRYB_19__4_), .S(SUMB_19__4_) );
  FA_X1 S2_19_5 ( .A(ab_19__5_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), .CO(
        CARRYB_19__5_), .S(SUMB_19__5_) );
  FA_X1 S2_19_6 ( .A(ab_19__6_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), .CO(
        CARRYB_19__6_), .S(SUMB_19__6_) );
  FA_X1 S2_19_7 ( .A(ab_19__7_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), .CO(
        CARRYB_19__7_), .S(SUMB_19__7_) );
  FA_X1 S2_19_8 ( .A(ab_19__8_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), .CO(
        CARRYB_19__8_), .S(SUMB_19__8_) );
  FA_X1 S2_19_9 ( .A(ab_19__9_), .B(CARRYB_18__9_), .CI(SUMB_18__10_), .CO(
        CARRYB_19__9_), .S(SUMB_19__9_) );
  FA_X1 S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), .CO(
        CARRYB_19__10_), .S(SUMB_19__10_) );
  FA_X1 S2_19_11 ( .A(ab_19__11_), .B(CARRYB_18__11_), .CI(SUMB_18__12_), .CO(
        CARRYB_19__11_), .S(SUMB_19__11_) );
  FA_X1 S2_19_12 ( .A(ab_19__12_), .B(CARRYB_18__12_), .CI(SUMB_18__13_), .CO(
        CARRYB_19__12_), .S(SUMB_19__12_) );
  FA_X1 S2_19_13 ( .A(ab_19__13_), .B(CARRYB_18__13_), .CI(SUMB_18__14_), .CO(
        CARRYB_19__13_), .S(SUMB_19__13_) );
  FA_X1 S2_19_14 ( .A(ab_19__14_), .B(CARRYB_18__14_), .CI(SUMB_18__15_), .CO(
        CARRYB_19__14_), .S(SUMB_19__14_) );
  FA_X1 S2_19_15 ( .A(ab_19__15_), .B(CARRYB_18__15_), .CI(SUMB_18__16_), .CO(
        CARRYB_19__15_), .S(SUMB_19__15_) );
  FA_X1 S2_19_16 ( .A(ab_19__16_), .B(CARRYB_18__16_), .CI(SUMB_18__17_), .CO(
        CARRYB_19__16_), .S(SUMB_19__16_) );
  FA_X1 S2_19_17 ( .A(ab_19__17_), .B(CARRYB_18__17_), .CI(SUMB_18__18_), .CO(
        CARRYB_19__17_), .S(SUMB_19__17_) );
  FA_X1 S2_19_18 ( .A(ab_19__18_), .B(CARRYB_18__18_), .CI(SUMB_18__19_), .CO(
        CARRYB_19__18_), .S(SUMB_19__18_) );
  FA_X1 S2_19_19 ( .A(ab_19__19_), .B(CARRYB_18__19_), .CI(SUMB_18__20_), .CO(
        CARRYB_19__19_), .S(SUMB_19__19_) );
  FA_X1 S2_19_20 ( .A(ab_19__20_), .B(CARRYB_18__20_), .CI(SUMB_18__21_), .CO(
        CARRYB_19__20_), .S(SUMB_19__20_) );
  FA_X1 S2_19_21 ( .A(ab_19__21_), .B(CARRYB_18__21_), .CI(SUMB_18__22_), .CO(
        CARRYB_19__21_), .S(SUMB_19__21_) );
  FA_X1 S3_19_22 ( .A(ab_19__22_), .B(CARRYB_18__22_), .CI(ab_18__23_), .CO(
        CARRYB_19__22_), .S(SUMB_19__22_) );
  FA_X1 S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), .CO(
        CARRYB_18__0_), .S(A1_16_) );
  FA_X1 S2_18_1 ( .A(ab_18__1_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), .CO(
        CARRYB_18__1_), .S(SUMB_18__1_) );
  FA_X1 S2_18_2 ( .A(ab_18__2_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), .CO(
        CARRYB_18__2_), .S(SUMB_18__2_) );
  FA_X1 S2_18_3 ( .A(ab_18__3_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), .CO(
        CARRYB_18__3_), .S(SUMB_18__3_) );
  FA_X1 S2_18_4 ( .A(ab_18__4_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), .CO(
        CARRYB_18__4_), .S(SUMB_18__4_) );
  FA_X1 S2_18_5 ( .A(ab_18__5_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), .CO(
        CARRYB_18__5_), .S(SUMB_18__5_) );
  FA_X1 S2_18_6 ( .A(ab_18__6_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), .CO(
        CARRYB_18__6_), .S(SUMB_18__6_) );
  FA_X1 S2_18_7 ( .A(ab_18__7_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), .CO(
        CARRYB_18__7_), .S(SUMB_18__7_) );
  FA_X1 S2_18_8 ( .A(ab_18__8_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), .CO(
        CARRYB_18__8_), .S(SUMB_18__8_) );
  FA_X1 S2_18_9 ( .A(ab_18__9_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), .CO(
        CARRYB_18__9_), .S(SUMB_18__9_) );
  FA_X1 S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), .CO(
        CARRYB_18__10_), .S(SUMB_18__10_) );
  FA_X1 S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), .CO(
        CARRYB_18__11_), .S(SUMB_18__11_) );
  FA_X1 S2_18_12 ( .A(ab_18__12_), .B(CARRYB_17__12_), .CI(SUMB_17__13_), .CO(
        CARRYB_18__12_), .S(SUMB_18__12_) );
  FA_X1 S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .CI(SUMB_17__14_), .CO(
        CARRYB_18__13_), .S(SUMB_18__13_) );
  FA_X1 S2_18_14 ( .A(ab_18__14_), .B(CARRYB_17__14_), .CI(SUMB_17__15_), .CO(
        CARRYB_18__14_), .S(SUMB_18__14_) );
  FA_X1 S2_18_15 ( .A(ab_18__15_), .B(CARRYB_17__15_), .CI(SUMB_17__16_), .CO(
        CARRYB_18__15_), .S(SUMB_18__15_) );
  FA_X1 S2_18_16 ( .A(ab_18__16_), .B(CARRYB_17__16_), .CI(SUMB_17__17_), .CO(
        CARRYB_18__16_), .S(SUMB_18__16_) );
  FA_X1 S2_18_17 ( .A(ab_18__17_), .B(CARRYB_17__17_), .CI(SUMB_17__18_), .CO(
        CARRYB_18__17_), .S(SUMB_18__17_) );
  FA_X1 S2_18_18 ( .A(ab_18__18_), .B(CARRYB_17__18_), .CI(SUMB_17__19_), .CO(
        CARRYB_18__18_), .S(SUMB_18__18_) );
  FA_X1 S2_18_19 ( .A(ab_18__19_), .B(CARRYB_17__19_), .CI(SUMB_17__20_), .CO(
        CARRYB_18__19_), .S(SUMB_18__19_) );
  FA_X1 S2_18_20 ( .A(ab_18__20_), .B(CARRYB_17__20_), .CI(SUMB_17__21_), .CO(
        CARRYB_18__20_), .S(SUMB_18__20_) );
  FA_X1 S2_18_21 ( .A(ab_18__21_), .B(CARRYB_17__21_), .CI(SUMB_17__22_), .CO(
        CARRYB_18__21_), .S(SUMB_18__21_) );
  FA_X1 S3_18_22 ( .A(ab_18__22_), .B(CARRYB_17__22_), .CI(ab_17__23_), .CO(
        CARRYB_18__22_), .S(SUMB_18__22_) );
  FA_X1 S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), .CO(
        CARRYB_17__0_), .S(A1_15_) );
  FA_X1 S2_17_1 ( .A(ab_17__1_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), .CO(
        CARRYB_17__1_), .S(SUMB_17__1_) );
  FA_X1 S2_17_2 ( .A(ab_17__2_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), .CO(
        CARRYB_17__2_), .S(SUMB_17__2_) );
  FA_X1 S2_17_3 ( .A(ab_17__3_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), .CO(
        CARRYB_17__3_), .S(SUMB_17__3_) );
  FA_X1 S2_17_4 ( .A(ab_17__4_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), .CO(
        CARRYB_17__4_), .S(SUMB_17__4_) );
  FA_X1 S2_17_5 ( .A(ab_17__5_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), .CO(
        CARRYB_17__5_), .S(SUMB_17__5_) );
  FA_X1 S2_17_6 ( .A(ab_17__6_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), .CO(
        CARRYB_17__6_), .S(SUMB_17__6_) );
  FA_X1 S2_17_7 ( .A(ab_17__7_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), .CO(
        CARRYB_17__7_), .S(SUMB_17__7_) );
  FA_X1 S2_17_8 ( .A(ab_17__8_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), .CO(
        CARRYB_17__8_), .S(SUMB_17__8_) );
  FA_X1 S2_17_9 ( .A(ab_17__9_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), .CO(
        CARRYB_17__9_), .S(SUMB_17__9_) );
  FA_X1 S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), .CO(
        CARRYB_17__10_), .S(SUMB_17__10_) );
  FA_X1 S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), .CO(
        CARRYB_17__11_), .S(SUMB_17__11_) );
  FA_X1 S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), .CO(
        CARRYB_17__12_), .S(SUMB_17__12_) );
  FA_X1 S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), .CO(
        CARRYB_17__13_), .S(SUMB_17__13_) );
  FA_X1 S2_17_14 ( .A(ab_17__14_), .B(CARRYB_16__14_), .CI(SUMB_16__15_), .CO(
        CARRYB_17__14_), .S(SUMB_17__14_) );
  FA_X1 S2_17_15 ( .A(ab_17__15_), .B(CARRYB_16__15_), .CI(SUMB_16__16_), .CO(
        CARRYB_17__15_), .S(SUMB_17__15_) );
  FA_X1 S2_17_16 ( .A(ab_17__16_), .B(CARRYB_16__16_), .CI(SUMB_16__17_), .CO(
        CARRYB_17__16_), .S(SUMB_17__16_) );
  FA_X1 S2_17_17 ( .A(ab_17__17_), .B(CARRYB_16__17_), .CI(SUMB_16__18_), .CO(
        CARRYB_17__17_), .S(SUMB_17__17_) );
  FA_X1 S2_17_18 ( .A(ab_17__18_), .B(CARRYB_16__18_), .CI(SUMB_16__19_), .CO(
        CARRYB_17__18_), .S(SUMB_17__18_) );
  FA_X1 S2_17_19 ( .A(ab_17__19_), .B(CARRYB_16__19_), .CI(SUMB_16__20_), .CO(
        CARRYB_17__19_), .S(SUMB_17__19_) );
  FA_X1 S2_17_20 ( .A(ab_17__20_), .B(CARRYB_16__20_), .CI(SUMB_16__21_), .CO(
        CARRYB_17__20_), .S(SUMB_17__20_) );
  FA_X1 S2_17_21 ( .A(ab_17__21_), .B(CARRYB_16__21_), .CI(SUMB_16__22_), .CO(
        CARRYB_17__21_), .S(SUMB_17__21_) );
  FA_X1 S3_17_22 ( .A(ab_17__22_), .B(CARRYB_16__22_), .CI(ab_16__23_), .CO(
        CARRYB_17__22_), .S(SUMB_17__22_) );
  FA_X1 S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(A1_14_) );
  FA_X1 S2_16_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  FA_X1 S2_16_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  FA_X1 S2_16_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  FA_X1 S2_16_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  FA_X1 S2_16_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  FA_X1 S2_16_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  FA_X1 S2_16_7 ( .A(ab_16__7_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), .CO(
        CARRYB_16__7_), .S(SUMB_16__7_) );
  FA_X1 S2_16_8 ( .A(ab_16__8_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), .CO(
        CARRYB_16__8_), .S(SUMB_16__8_) );
  FA_X1 S2_16_9 ( .A(ab_16__9_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), .CO(
        CARRYB_16__9_), .S(SUMB_16__9_) );
  FA_X1 S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), .CO(
        CARRYB_16__10_), .S(SUMB_16__10_) );
  FA_X1 S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), .CO(
        CARRYB_16__11_), .S(SUMB_16__11_) );
  FA_X1 S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), .CO(
        CARRYB_16__12_), .S(SUMB_16__12_) );
  FA_X1 S2_16_13 ( .A(ab_16__13_), .B(CARRYB_15__13_), .CI(SUMB_15__14_), .CO(
        CARRYB_16__13_), .S(SUMB_16__13_) );
  FA_X1 S2_16_14 ( .A(ab_16__14_), .B(CARRYB_15__14_), .CI(SUMB_15__15_), .CO(
        CARRYB_16__14_), .S(SUMB_16__14_) );
  FA_X1 S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .CI(SUMB_15__16_), .CO(
        CARRYB_16__15_), .S(SUMB_16__15_) );
  FA_X1 S2_16_16 ( .A(ab_16__16_), .B(CARRYB_15__16_), .CI(SUMB_15__17_), .CO(
        CARRYB_16__16_), .S(SUMB_16__16_) );
  FA_X1 S2_16_17 ( .A(ab_16__17_), .B(CARRYB_15__17_), .CI(SUMB_15__18_), .CO(
        CARRYB_16__17_), .S(SUMB_16__17_) );
  FA_X1 S2_16_18 ( .A(ab_16__18_), .B(CARRYB_15__18_), .CI(SUMB_15__19_), .CO(
        CARRYB_16__18_), .S(SUMB_16__18_) );
  FA_X1 S2_16_19 ( .A(ab_16__19_), .B(CARRYB_15__19_), .CI(SUMB_15__20_), .CO(
        CARRYB_16__19_), .S(SUMB_16__19_) );
  FA_X1 S2_16_20 ( .A(ab_16__20_), .B(CARRYB_15__20_), .CI(SUMB_15__21_), .CO(
        CARRYB_16__20_), .S(SUMB_16__20_) );
  FA_X1 S2_16_21 ( .A(ab_16__21_), .B(CARRYB_15__21_), .CI(SUMB_15__22_), .CO(
        CARRYB_16__21_), .S(SUMB_16__21_) );
  FA_X1 S3_16_22 ( .A(ab_16__22_), .B(CARRYB_15__22_), .CI(ab_15__23_), .CO(
        CARRYB_16__22_), .S(SUMB_16__22_) );
  FA_X1 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  FA_X1 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  FA_X1 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  FA_X1 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  FA_X1 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  FA_X1 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  FA_X1 S2_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  FA_X1 S2_15_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), .CO(
        CARRYB_15__7_), .S(SUMB_15__7_) );
  FA_X1 S2_15_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), .CO(
        CARRYB_15__8_), .S(SUMB_15__8_) );
  FA_X1 S2_15_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), .CO(
        CARRYB_15__9_), .S(SUMB_15__9_) );
  FA_X1 S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), .CO(
        CARRYB_15__10_), .S(SUMB_15__10_) );
  FA_X1 S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), .CO(
        CARRYB_15__11_), .S(SUMB_15__11_) );
  FA_X1 S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), .CO(
        CARRYB_15__12_), .S(SUMB_15__12_) );
  FA_X1 S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), .CO(
        CARRYB_15__13_), .S(SUMB_15__13_) );
  FA_X1 S2_15_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), .CO(
        CARRYB_15__14_), .S(SUMB_15__14_) );
  FA_X1 S2_15_15 ( .A(ab_15__15_), .B(CARRYB_14__15_), .CI(SUMB_14__16_), .CO(
        CARRYB_15__15_), .S(SUMB_15__15_) );
  FA_X1 S2_15_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .CI(SUMB_14__17_), .CO(
        CARRYB_15__16_), .S(SUMB_15__16_) );
  FA_X1 S2_15_17 ( .A(ab_15__17_), .B(CARRYB_14__17_), .CI(SUMB_14__18_), .CO(
        CARRYB_15__17_), .S(SUMB_15__17_) );
  FA_X1 S2_15_18 ( .A(ab_15__18_), .B(CARRYB_14__18_), .CI(SUMB_14__19_), .CO(
        CARRYB_15__18_), .S(SUMB_15__18_) );
  FA_X1 S2_15_19 ( .A(ab_15__19_), .B(CARRYB_14__19_), .CI(SUMB_14__20_), .CO(
        CARRYB_15__19_), .S(SUMB_15__19_) );
  FA_X1 S2_15_20 ( .A(ab_15__20_), .B(CARRYB_14__20_), .CI(SUMB_14__21_), .CO(
        CARRYB_15__20_), .S(SUMB_15__20_) );
  FA_X1 S2_15_21 ( .A(ab_15__21_), .B(CARRYB_14__21_), .CI(SUMB_14__22_), .CO(
        CARRYB_15__21_), .S(SUMB_15__21_) );
  FA_X1 S3_15_22 ( .A(ab_15__22_), .B(CARRYB_14__22_), .CI(ab_14__23_), .CO(
        CARRYB_15__22_), .S(SUMB_15__22_) );
  FA_X1 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  FA_X1 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  FA_X1 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  FA_X1 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  FA_X1 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  FA_X1 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  FA_X1 S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  FA_X1 S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), .CO(
        CARRYB_14__7_), .S(SUMB_14__7_) );
  FA_X1 S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), .CO(
        CARRYB_14__8_), .S(SUMB_14__8_) );
  FA_X1 S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), .CO(
        CARRYB_14__9_), .S(SUMB_14__9_) );
  FA_X1 S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), .CO(
        CARRYB_14__10_), .S(SUMB_14__10_) );
  FA_X1 S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), .CO(
        CARRYB_14__11_), .S(SUMB_14__11_) );
  FA_X1 S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), .CO(
        CARRYB_14__12_), .S(SUMB_14__12_) );
  FA_X1 S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), .CO(
        CARRYB_14__13_), .S(SUMB_14__13_) );
  FA_X1 S2_14_14 ( .A(ab_14__14_), .B(CARRYB_13__14_), .CI(SUMB_13__15_), .CO(
        CARRYB_14__14_), .S(SUMB_14__14_) );
  FA_X1 S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), .CO(
        CARRYB_14__15_), .S(SUMB_14__15_) );
  FA_X1 S2_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), .CO(
        CARRYB_14__16_), .S(SUMB_14__16_) );
  FA_X1 S2_14_17 ( .A(ab_14__17_), .B(CARRYB_13__17_), .CI(SUMB_13__18_), .CO(
        CARRYB_14__17_), .S(SUMB_14__17_) );
  FA_X1 S2_14_18 ( .A(ab_14__18_), .B(CARRYB_13__18_), .CI(SUMB_13__19_), .CO(
        CARRYB_14__18_), .S(SUMB_14__18_) );
  FA_X1 S2_14_19 ( .A(ab_14__19_), .B(CARRYB_13__19_), .CI(SUMB_13__20_), .CO(
        CARRYB_14__19_), .S(SUMB_14__19_) );
  FA_X1 S2_14_20 ( .A(ab_14__20_), .B(CARRYB_13__20_), .CI(SUMB_13__21_), .CO(
        CARRYB_14__20_), .S(SUMB_14__20_) );
  FA_X1 S2_14_21 ( .A(ab_14__21_), .B(CARRYB_13__21_), .CI(SUMB_13__22_), .CO(
        CARRYB_14__21_), .S(SUMB_14__21_) );
  FA_X1 S3_14_22 ( .A(ab_14__22_), .B(CARRYB_13__22_), .CI(ab_13__23_), .CO(
        CARRYB_14__22_), .S(SUMB_14__22_) );
  FA_X1 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  FA_X1 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  FA_X1 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  FA_X1 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  FA_X1 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  FA_X1 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  FA_X1 S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  FA_X1 S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), .CO(
        CARRYB_13__7_), .S(SUMB_13__7_) );
  FA_X1 S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), .CO(
        CARRYB_13__8_), .S(SUMB_13__8_) );
  FA_X1 S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), .CO(
        CARRYB_13__9_), .S(SUMB_13__9_) );
  FA_X1 S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), .CO(
        CARRYB_13__10_), .S(SUMB_13__10_) );
  FA_X1 S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), .CO(
        CARRYB_13__11_), .S(SUMB_13__11_) );
  FA_X1 S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), .CO(
        CARRYB_13__12_), .S(SUMB_13__12_) );
  FA_X1 S2_13_13 ( .A(ab_13__13_), .B(CARRYB_12__13_), .CI(SUMB_12__14_), .CO(
        CARRYB_13__13_), .S(SUMB_13__13_) );
  FA_X1 S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), .CO(
        CARRYB_13__14_), .S(SUMB_13__14_) );
  FA_X1 S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), .CO(
        CARRYB_13__15_), .S(SUMB_13__15_) );
  FA_X1 S2_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), .CO(
        CARRYB_13__16_), .S(SUMB_13__16_) );
  FA_X1 S2_13_17 ( .A(ab_13__17_), .B(CARRYB_12__17_), .CI(SUMB_12__18_), .CO(
        CARRYB_13__17_), .S(SUMB_13__17_) );
  FA_X1 S2_13_18 ( .A(ab_13__18_), .B(CARRYB_12__18_), .CI(SUMB_12__19_), .CO(
        CARRYB_13__18_), .S(SUMB_13__18_) );
  FA_X1 S2_13_19 ( .A(ab_13__19_), .B(CARRYB_12__19_), .CI(SUMB_12__20_), .CO(
        CARRYB_13__19_), .S(SUMB_13__19_) );
  FA_X1 S2_13_20 ( .A(ab_13__20_), .B(CARRYB_12__20_), .CI(SUMB_12__21_), .CO(
        CARRYB_13__20_), .S(SUMB_13__20_) );
  FA_X1 S2_13_21 ( .A(ab_13__21_), .B(CARRYB_12__21_), .CI(SUMB_12__22_), .CO(
        CARRYB_13__21_), .S(SUMB_13__21_) );
  FA_X1 S3_13_22 ( .A(ab_13__22_), .B(CARRYB_12__22_), .CI(ab_12__23_), .CO(
        CARRYB_13__22_), .S(SUMB_13__22_) );
  FA_X1 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  FA_X1 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  FA_X1 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  FA_X1 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  FA_X1 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  FA_X1 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  FA_X1 S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  FA_X1 S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), .CO(
        CARRYB_12__7_), .S(SUMB_12__7_) );
  FA_X1 S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), .CO(
        CARRYB_12__8_), .S(SUMB_12__8_) );
  FA_X1 S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), .CO(
        CARRYB_12__9_), .S(SUMB_12__9_) );
  FA_X1 S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), .CO(
        CARRYB_12__10_), .S(SUMB_12__10_) );
  FA_X1 S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), .CO(
        CARRYB_12__11_), .S(SUMB_12__11_) );
  FA_X1 S2_12_12 ( .A(ab_12__12_), .B(CARRYB_11__12_), .CI(SUMB_11__13_), .CO(
        CARRYB_12__12_), .S(SUMB_12__12_) );
  FA_X1 S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), .CO(
        CARRYB_12__13_), .S(SUMB_12__13_) );
  FA_X1 S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), .CO(
        CARRYB_12__14_), .S(SUMB_12__14_) );
  FA_X1 S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), .CO(
        CARRYB_12__15_), .S(SUMB_12__15_) );
  FA_X1 S2_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), .CO(
        CARRYB_12__16_), .S(SUMB_12__16_) );
  FA_X1 S2_12_17 ( .A(ab_12__17_), .B(CARRYB_11__17_), .CI(SUMB_11__18_), .CO(
        CARRYB_12__17_), .S(SUMB_12__17_) );
  FA_X1 S2_12_18 ( .A(ab_12__18_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), .CO(
        CARRYB_12__18_), .S(SUMB_12__18_) );
  FA_X1 S2_12_19 ( .A(ab_12__19_), .B(CARRYB_11__19_), .CI(SUMB_11__20_), .CO(
        CARRYB_12__19_), .S(SUMB_12__19_) );
  FA_X1 S2_12_20 ( .A(ab_12__20_), .B(CARRYB_11__20_), .CI(SUMB_11__21_), .CO(
        CARRYB_12__20_), .S(SUMB_12__20_) );
  FA_X1 S2_12_21 ( .A(ab_12__21_), .B(CARRYB_11__21_), .CI(SUMB_11__22_), .CO(
        CARRYB_12__21_), .S(SUMB_12__21_) );
  FA_X1 S3_12_22 ( .A(ab_12__22_), .B(CARRYB_11__22_), .CI(ab_11__23_), .CO(
        CARRYB_12__22_), .S(SUMB_12__22_) );
  FA_X1 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  FA_X1 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  FA_X1 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  FA_X1 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  FA_X1 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  FA_X1 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  FA_X1 S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  FA_X1 S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), .CO(
        CARRYB_11__7_), .S(SUMB_11__7_) );
  FA_X1 S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), .CO(
        CARRYB_11__8_), .S(SUMB_11__8_) );
  FA_X1 S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), .CO(
        CARRYB_11__9_), .S(SUMB_11__9_) );
  FA_X1 S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), .CO(
        CARRYB_11__10_), .S(SUMB_11__10_) );
  FA_X1 S2_11_11 ( .A(ab_11__11_), .B(CARRYB_10__11_), .CI(SUMB_10__12_), .CO(
        CARRYB_11__11_), .S(SUMB_11__11_) );
  FA_X1 S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), .CO(
        CARRYB_11__12_), .S(SUMB_11__12_) );
  FA_X1 S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), .CO(
        CARRYB_11__13_), .S(SUMB_11__13_) );
  FA_X1 S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), .CO(
        CARRYB_11__14_), .S(SUMB_11__14_) );
  FA_X1 S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), .CO(
        CARRYB_11__15_), .S(SUMB_11__15_) );
  FA_X1 S2_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(SUMB_10__17_), .CO(
        CARRYB_11__16_), .S(SUMB_11__16_) );
  FA_X1 S2_11_17 ( .A(ab_11__17_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), .CO(
        CARRYB_11__17_), .S(SUMB_11__17_) );
  FA_X1 S2_11_18 ( .A(ab_11__18_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), .CO(
        CARRYB_11__18_), .S(SUMB_11__18_) );
  FA_X1 S2_11_19 ( .A(ab_11__19_), .B(CARRYB_10__19_), .CI(SUMB_10__20_), .CO(
        CARRYB_11__19_), .S(SUMB_11__19_) );
  FA_X1 S2_11_20 ( .A(ab_11__20_), .B(CARRYB_10__20_), .CI(SUMB_10__21_), .CO(
        CARRYB_11__20_), .S(SUMB_11__20_) );
  FA_X1 S2_11_21 ( .A(ab_11__21_), .B(CARRYB_10__21_), .CI(SUMB_10__22_), .CO(
        CARRYB_11__21_), .S(SUMB_11__21_) );
  FA_X1 S3_11_22 ( .A(ab_11__22_), .B(CARRYB_10__22_), .CI(ab_10__23_), .CO(
        CARRYB_11__22_), .S(SUMB_11__22_) );
  FA_X1 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  FA_X1 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  FA_X1 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  FA_X1 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  FA_X1 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  FA_X1 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  FA_X1 S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  FA_X1 S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  FA_X1 S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  FA_X1 S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  FA_X1 S2_10_10 ( .A(ab_10__10_), .B(CARRYB_9__10_), .CI(SUMB_9__11_), .CO(
        CARRYB_10__10_), .S(SUMB_10__10_) );
  FA_X1 S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), .CO(
        CARRYB_10__11_), .S(SUMB_10__11_) );
  FA_X1 S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), .CO(
        CARRYB_10__12_), .S(SUMB_10__12_) );
  FA_X1 S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), .CO(
        CARRYB_10__13_), .S(SUMB_10__13_) );
  FA_X1 S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), .CO(
        CARRYB_10__14_), .S(SUMB_10__14_) );
  FA_X1 S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), .CO(
        CARRYB_10__15_), .S(SUMB_10__15_) );
  FA_X1 S2_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), .CO(
        CARRYB_10__16_), .S(SUMB_10__16_) );
  FA_X1 S2_10_17 ( .A(ab_10__17_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), .CO(
        CARRYB_10__17_), .S(SUMB_10__17_) );
  FA_X1 S2_10_18 ( .A(ab_10__18_), .B(CARRYB_9__18_), .CI(SUMB_9__19_), .CO(
        CARRYB_10__18_), .S(SUMB_10__18_) );
  FA_X1 S2_10_19 ( .A(ab_10__19_), .B(CARRYB_9__19_), .CI(SUMB_9__20_), .CO(
        CARRYB_10__19_), .S(SUMB_10__19_) );
  FA_X1 S2_10_20 ( .A(ab_10__20_), .B(CARRYB_9__20_), .CI(SUMB_9__21_), .CO(
        CARRYB_10__20_), .S(SUMB_10__20_) );
  FA_X1 S2_10_21 ( .A(ab_10__21_), .B(CARRYB_9__21_), .CI(SUMB_9__22_), .CO(
        CARRYB_10__21_), .S(SUMB_10__21_) );
  FA_X1 S3_10_22 ( .A(ab_10__22_), .B(CARRYB_9__22_), .CI(ab_9__23_), .CO(
        CARRYB_10__22_), .S(SUMB_10__22_) );
  FA_X1 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  FA_X1 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  FA_X1 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  FA_X1 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  FA_X1 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  FA_X1 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  FA_X1 S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  FA_X1 S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  FA_X1 S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  FA_X1 S2_9_9 ( .A(ab_9__9_), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  FA_X1 S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), .CO(
        CARRYB_9__10_), .S(SUMB_9__10_) );
  FA_X1 S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), .CO(
        CARRYB_9__11_), .S(SUMB_9__11_) );
  FA_X1 S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), .CO(
        CARRYB_9__12_), .S(SUMB_9__12_) );
  FA_X1 S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), .CO(
        CARRYB_9__13_), .S(SUMB_9__13_) );
  FA_X1 S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), .CO(
        CARRYB_9__14_), .S(SUMB_9__14_) );
  FA_X1 S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), .CO(
        CARRYB_9__15_), .S(SUMB_9__15_) );
  FA_X1 S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), .CO(
        CARRYB_9__16_), .S(SUMB_9__16_) );
  FA_X1 S2_9_17 ( .A(ab_9__17_), .B(CARRYB_8__17_), .CI(SUMB_8__18_), .CO(
        CARRYB_9__17_), .S(SUMB_9__17_) );
  FA_X1 S2_9_18 ( .A(ab_9__18_), .B(CARRYB_8__18_), .CI(SUMB_8__19_), .CO(
        CARRYB_9__18_), .S(SUMB_9__18_) );
  FA_X1 S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), .CO(
        CARRYB_9__19_), .S(SUMB_9__19_) );
  FA_X1 S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(SUMB_8__21_), .CO(
        CARRYB_9__20_), .S(SUMB_9__20_) );
  FA_X1 S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), .CO(
        CARRYB_9__21_), .S(SUMB_9__21_) );
  FA_X1 S3_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .CI(ab_8__23_), .CO(
        CARRYB_9__22_), .S(SUMB_9__22_) );
  FA_X1 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  FA_X1 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  FA_X1 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  FA_X1 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  FA_X1 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  FA_X1 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  FA_X1 S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  FA_X1 S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  FA_X1 S2_8_8 ( .A(ab_8__8_), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  FA_X1 S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  FA_X1 S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), .CO(
        CARRYB_8__10_), .S(SUMB_8__10_) );
  FA_X1 S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), .CO(
        CARRYB_8__11_), .S(SUMB_8__11_) );
  FA_X1 S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), .CO(
        CARRYB_8__12_), .S(SUMB_8__12_) );
  FA_X1 S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), .CO(
        CARRYB_8__13_), .S(SUMB_8__13_) );
  FA_X1 S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), .CO(
        CARRYB_8__14_), .S(SUMB_8__14_) );
  FA_X1 S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), .CO(
        CARRYB_8__15_), .S(SUMB_8__15_) );
  FA_X1 S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), .CO(
        CARRYB_8__16_), .S(SUMB_8__16_) );
  FA_X1 S2_8_17 ( .A(ab_8__17_), .B(CARRYB_7__17_), .CI(SUMB_7__18_), .CO(
        CARRYB_8__17_), .S(SUMB_8__17_) );
  FA_X1 S2_8_18 ( .A(ab_8__18_), .B(CARRYB_7__18_), .CI(SUMB_7__19_), .CO(
        CARRYB_8__18_), .S(SUMB_8__18_) );
  FA_X1 S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), .CO(
        CARRYB_8__19_), .S(SUMB_8__19_) );
  FA_X1 S2_8_20 ( .A(ab_8__20_), .B(CARRYB_7__20_), .CI(SUMB_7__21_), .CO(
        CARRYB_8__20_), .S(SUMB_8__20_) );
  FA_X1 S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), .CO(
        CARRYB_8__21_), .S(SUMB_8__21_) );
  FA_X1 S3_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(ab_7__23_), .CO(
        CARRYB_8__22_), .S(SUMB_8__22_) );
  FA_X1 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(A1_5_) );
  FA_X1 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S2_7_7 ( .A(ab_7__7_), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  FA_X1 S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  FA_X1 S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  FA_X1 S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), .CO(
        CARRYB_7__10_), .S(SUMB_7__10_) );
  FA_X1 S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), .CO(
        CARRYB_7__11_), .S(SUMB_7__11_) );
  FA_X1 S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), .CO(
        CARRYB_7__12_), .S(SUMB_7__12_) );
  FA_X1 S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), .CO(
        CARRYB_7__13_), .S(SUMB_7__13_) );
  FA_X1 S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), .CO(
        CARRYB_7__14_), .S(SUMB_7__14_) );
  FA_X1 S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), .CO(
        CARRYB_7__15_), .S(SUMB_7__15_) );
  FA_X1 S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), .CO(
        CARRYB_7__16_), .S(SUMB_7__16_) );
  FA_X1 S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), .CO(
        CARRYB_7__17_), .S(SUMB_7__17_) );
  FA_X1 S2_7_18 ( .A(ab_7__18_), .B(CARRYB_6__18_), .CI(SUMB_6__19_), .CO(
        CARRYB_7__18_), .S(SUMB_7__18_) );
  FA_X1 S2_7_19 ( .A(ab_7__19_), .B(CARRYB_6__19_), .CI(SUMB_6__20_), .CO(
        CARRYB_7__19_), .S(SUMB_7__19_) );
  FA_X1 S2_7_20 ( .A(ab_7__20_), .B(CARRYB_6__20_), .CI(SUMB_6__21_), .CO(
        CARRYB_7__20_), .S(SUMB_7__20_) );
  FA_X1 S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), .CO(
        CARRYB_7__21_), .S(SUMB_7__21_) );
  FA_X1 S3_7_22 ( .A(ab_7__22_), .B(CARRYB_6__22_), .CI(ab_6__23_), .CO(
        CARRYB_7__22_), .S(SUMB_7__22_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S2_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  FA_X1 S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  FA_X1 S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  FA_X1 S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), .CO(
        CARRYB_6__10_), .S(SUMB_6__10_) );
  FA_X1 S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), .CO(
        CARRYB_6__11_), .S(SUMB_6__11_) );
  FA_X1 S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), .CO(
        CARRYB_6__12_), .S(SUMB_6__12_) );
  FA_X1 S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), .CO(
        CARRYB_6__13_), .S(SUMB_6__13_) );
  FA_X1 S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), .CO(
        CARRYB_6__14_), .S(SUMB_6__14_) );
  FA_X1 S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), .CO(
        CARRYB_6__15_), .S(SUMB_6__15_) );
  FA_X1 S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), .CO(
        CARRYB_6__16_), .S(SUMB_6__16_) );
  FA_X1 S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), .CO(
        CARRYB_6__17_), .S(SUMB_6__17_) );
  FA_X1 S2_6_18 ( .A(ab_6__18_), .B(CARRYB_5__18_), .CI(SUMB_5__19_), .CO(
        CARRYB_6__18_), .S(SUMB_6__18_) );
  FA_X1 S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), .CO(
        CARRYB_6__19_), .S(SUMB_6__19_) );
  FA_X1 S2_6_20 ( .A(ab_6__20_), .B(CARRYB_5__20_), .CI(SUMB_5__21_), .CO(
        CARRYB_6__20_), .S(SUMB_6__20_) );
  FA_X1 S2_6_21 ( .A(ab_6__21_), .B(CARRYB_5__21_), .CI(SUMB_5__22_), .CO(
        CARRYB_6__21_), .S(SUMB_6__21_) );
  FA_X1 S3_6_22 ( .A(ab_6__22_), .B(CARRYB_5__22_), .CI(ab_5__23_), .CO(
        CARRYB_6__22_), .S(SUMB_6__22_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  FA_X1 S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  FA_X1 S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  FA_X1 S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), .CO(
        CARRYB_5__10_), .S(SUMB_5__10_) );
  FA_X1 S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), .CO(
        CARRYB_5__11_), .S(SUMB_5__11_) );
  FA_X1 S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), .CO(
        CARRYB_5__12_), .S(SUMB_5__12_) );
  FA_X1 S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), .CO(
        CARRYB_5__13_), .S(SUMB_5__13_) );
  FA_X1 S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), .CO(
        CARRYB_5__14_), .S(SUMB_5__14_) );
  FA_X1 S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), .CO(
        CARRYB_5__15_), .S(SUMB_5__15_) );
  FA_X1 S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), .CO(
        CARRYB_5__16_), .S(SUMB_5__16_) );
  FA_X1 S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), .CO(
        CARRYB_5__17_), .S(SUMB_5__17_) );
  FA_X1 S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), .CO(
        CARRYB_5__18_), .S(SUMB_5__18_) );
  FA_X1 S2_5_19 ( .A(ab_5__19_), .B(CARRYB_4__19_), .CI(SUMB_4__20_), .CO(
        CARRYB_5__19_), .S(SUMB_5__19_) );
  FA_X1 S2_5_20 ( .A(ab_5__20_), .B(CARRYB_4__20_), .CI(SUMB_4__21_), .CO(
        CARRYB_5__20_), .S(SUMB_5__20_) );
  FA_X1 S2_5_21 ( .A(ab_5__21_), .B(CARRYB_4__21_), .CI(SUMB_4__22_), .CO(
        CARRYB_5__21_), .S(SUMB_5__21_) );
  FA_X1 S3_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(ab_4__23_), .CO(
        CARRYB_5__22_), .S(SUMB_5__22_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  FA_X1 S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  FA_X1 S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  FA_X1 S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), .CO(
        CARRYB_4__10_), .S(SUMB_4__10_) );
  FA_X1 S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), .CO(
        CARRYB_4__11_), .S(SUMB_4__11_) );
  FA_X1 S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), .CO(
        CARRYB_4__12_), .S(SUMB_4__12_) );
  FA_X1 S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), .CO(
        CARRYB_4__13_), .S(SUMB_4__13_) );
  FA_X1 S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), .CO(
        CARRYB_4__14_), .S(SUMB_4__14_) );
  FA_X1 S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), .CO(
        CARRYB_4__15_), .S(SUMB_4__15_) );
  FA_X1 S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), .CO(
        CARRYB_4__16_), .S(SUMB_4__16_) );
  FA_X1 S2_4_17 ( .A(ab_4__17_), .B(CARRYB_3__17_), .CI(SUMB_3__18_), .CO(
        CARRYB_4__17_), .S(SUMB_4__17_) );
  FA_X1 S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), .CO(
        CARRYB_4__18_), .S(SUMB_4__18_) );
  FA_X1 S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), .CO(
        CARRYB_4__19_), .S(SUMB_4__19_) );
  FA_X1 S2_4_20 ( .A(ab_4__20_), .B(CARRYB_3__20_), .CI(SUMB_3__21_), .CO(
        CARRYB_4__20_), .S(SUMB_4__20_) );
  FA_X1 S2_4_21 ( .A(ab_4__21_), .B(CARRYB_3__21_), .CI(SUMB_3__22_), .CO(
        CARRYB_4__21_), .S(SUMB_4__21_) );
  FA_X1 S3_4_22 ( .A(ab_4__22_), .B(CARRYB_3__22_), .CI(ab_3__23_), .CO(
        CARRYB_4__22_), .S(SUMB_4__22_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  FA_X1 S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  FA_X1 S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  FA_X1 S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), .CO(
        CARRYB_3__10_), .S(SUMB_3__10_) );
  FA_X1 S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), .CO(
        CARRYB_3__11_), .S(SUMB_3__11_) );
  FA_X1 S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), .CO(
        CARRYB_3__12_), .S(SUMB_3__12_) );
  FA_X1 S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), .CO(
        CARRYB_3__13_), .S(SUMB_3__13_) );
  FA_X1 S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), .CO(
        CARRYB_3__14_), .S(SUMB_3__14_) );
  FA_X1 S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), .CO(
        CARRYB_3__15_), .S(SUMB_3__15_) );
  FA_X1 S2_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(SUMB_2__17_), .CO(
        CARRYB_3__16_), .S(SUMB_3__16_) );
  FA_X1 S2_3_17 ( .A(ab_3__17_), .B(CARRYB_2__17_), .CI(SUMB_2__18_), .CO(
        CARRYB_3__17_), .S(SUMB_3__17_) );
  FA_X1 S2_3_18 ( .A(ab_3__18_), .B(CARRYB_2__18_), .CI(SUMB_2__19_), .CO(
        CARRYB_3__18_), .S(SUMB_3__18_) );
  FA_X1 S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), .CO(
        CARRYB_3__19_), .S(SUMB_3__19_) );
  FA_X1 S2_3_20 ( .A(ab_3__20_), .B(CARRYB_2__20_), .CI(SUMB_2__21_), .CO(
        CARRYB_3__20_), .S(SUMB_3__20_) );
  FA_X1 S2_3_21 ( .A(ab_3__21_), .B(CARRYB_2__21_), .CI(SUMB_2__22_), .CO(
        CARRYB_3__21_), .S(SUMB_3__21_) );
  FA_X1 S3_3_22 ( .A(ab_3__22_), .B(CARRYB_2__22_), .CI(ab_2__23_), .CO(
        CARRYB_3__22_), .S(SUMB_3__22_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S2_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(SUMB_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  FA_X1 S2_2_7 ( .A(ab_2__7_), .B(CARRYB_1__7_), .CI(SUMB_1__8_), .CO(
        CARRYB_2__7_), .S(SUMB_2__7_) );
  FA_X1 S2_2_8 ( .A(ab_2__8_), .B(CARRYB_1__8_), .CI(SUMB_1__9_), .CO(
        CARRYB_2__8_), .S(SUMB_2__8_) );
  FA_X1 S2_2_9 ( .A(ab_2__9_), .B(CARRYB_1__9_), .CI(SUMB_1__10_), .CO(
        CARRYB_2__9_), .S(SUMB_2__9_) );
  FA_X1 S2_2_10 ( .A(ab_2__10_), .B(CARRYB_1__10_), .CI(SUMB_1__11_), .CO(
        CARRYB_2__10_), .S(SUMB_2__10_) );
  FA_X1 S2_2_11 ( .A(ab_2__11_), .B(CARRYB_1__11_), .CI(SUMB_1__12_), .CO(
        CARRYB_2__11_), .S(SUMB_2__11_) );
  FA_X1 S2_2_12 ( .A(ab_2__12_), .B(CARRYB_1__12_), .CI(SUMB_1__13_), .CO(
        CARRYB_2__12_), .S(SUMB_2__12_) );
  FA_X1 S2_2_13 ( .A(ab_2__13_), .B(CARRYB_1__13_), .CI(SUMB_1__14_), .CO(
        CARRYB_2__13_), .S(SUMB_2__13_) );
  FA_X1 S2_2_14 ( .A(ab_2__14_), .B(CARRYB_1__14_), .CI(SUMB_1__15_), .CO(
        CARRYB_2__14_), .S(SUMB_2__14_) );
  FA_X1 S2_2_15 ( .A(ab_2__15_), .B(CARRYB_1__15_), .CI(SUMB_1__16_), .CO(
        CARRYB_2__15_), .S(SUMB_2__15_) );
  FA_X1 S2_2_16 ( .A(ab_2__16_), .B(CARRYB_1__16_), .CI(SUMB_1__17_), .CO(
        CARRYB_2__16_), .S(SUMB_2__16_) );
  FA_X1 S2_2_17 ( .A(ab_2__17_), .B(CARRYB_1__17_), .CI(SUMB_1__18_), .CO(
        CARRYB_2__17_), .S(SUMB_2__17_) );
  FA_X1 S2_2_18 ( .A(ab_2__18_), .B(CARRYB_1__18_), .CI(SUMB_1__19_), .CO(
        CARRYB_2__18_), .S(SUMB_2__18_) );
  FA_X1 S2_2_19 ( .A(ab_2__19_), .B(CARRYB_1__19_), .CI(SUMB_1__20_), .CO(
        CARRYB_2__19_), .S(SUMB_2__19_) );
  FA_X1 S2_2_20 ( .A(ab_2__20_), .B(CARRYB_1__20_), .CI(SUMB_1__21_), .CO(
        CARRYB_2__20_), .S(SUMB_2__20_) );
  FA_X1 S2_2_21 ( .A(ab_2__21_), .B(CARRYB_1__21_), .CI(SUMB_1__22_), .CO(
        CARRYB_2__21_), .S(SUMB_2__21_) );
  FA_X1 S3_2_22 ( .A(ab_2__22_), .B(CARRYB_1__22_), .CI(ab_1__23_), .CO(
        CARRYB_2__22_), .S(SUMB_2__22_) );
  iir_filter_DW01_add_8 FS_1 ( .A({A1_45_, A1_44_, A1_43_, A1_42_, A1_41_, 
        A1_40_, A1_39_, A1_38_, A1_37_, A1_36_, A1_35_, A1_34_, A1_33_, A1_32_, 
        A1_31_, A1_30_, A1_29_, A1_28_, A1_27_, A1_26_, A1_25_, A1_24_, A1_23_, 
        A1_22_, A1_21_, A1_20_, A1_19_, A1_18_, A1_17_, A1_16_, A1_15_, A1_14_, 
        A1_13_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, A1_5_, 
        A1_4_, A1_3_, A1_2_, A1_1_, A1_0_}), .B({A2_45_, A2_44_, A2_43_, 
        A2_42_, A2_41_, A2_40_, A2_39_, A2_38_, A2_37_, A2_36_, A2_35_, A2_34_, 
        A2_33_, A2_32_, A2_31_, A2_30_, A2_29_, A2_28_, A2_27_, A2_26_, A2_25_, 
        A2_24_, A2_23_, A2_22_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({PRODUCT[47], SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, PRODUCT[44:22], SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21}) );
  BUF_X1 U2 ( .A(QB), .Z(n1) );
  BUF_X1 U3 ( .A(QB), .Z(n2) );
  BUF_X1 U4 ( .A(QA), .Z(n3) );
  BUF_X1 U5 ( .A(QA), .Z(n4) );
  INV_X1 U6 ( .A(B[22]), .ZN(n15) );
  INV_X1 U7 ( .A(B[21]), .ZN(n16) );
  INV_X1 U8 ( .A(B[20]), .ZN(n17) );
  INV_X1 U9 ( .A(B[19]), .ZN(n19) );
  INV_X1 U10 ( .A(B[18]), .ZN(n20) );
  INV_X1 U11 ( .A(B[17]), .ZN(n21) );
  INV_X1 U12 ( .A(B[16]), .ZN(n22) );
  INV_X1 U13 ( .A(B[15]), .ZN(n23) );
  INV_X1 U14 ( .A(B[14]), .ZN(n24) );
  INV_X1 U15 ( .A(B[13]), .ZN(n25) );
  INV_X1 U16 ( .A(B[12]), .ZN(n26) );
  INV_X1 U17 ( .A(B[11]), .ZN(n27) );
  INV_X1 U18 ( .A(B[10]), .ZN(n28) );
  INV_X1 U19 ( .A(B[9]), .ZN(n7) );
  INV_X1 U20 ( .A(B[8]), .ZN(n8) );
  INV_X1 U21 ( .A(B[7]), .ZN(n9) );
  INV_X1 U22 ( .A(B[6]), .ZN(n10) );
  INV_X1 U23 ( .A(B[5]), .ZN(n11) );
  INV_X1 U24 ( .A(B[4]), .ZN(n12) );
  INV_X1 U25 ( .A(B[3]), .ZN(n13) );
  INV_X1 U26 ( .A(B[2]), .ZN(n14) );
  INV_X1 U27 ( .A(A[2]), .ZN(n36) );
  INV_X1 U28 ( .A(A[3]), .ZN(n35) );
  INV_X1 U29 ( .A(A[4]), .ZN(n34) );
  INV_X1 U30 ( .A(A[5]), .ZN(n33) );
  INV_X1 U31 ( .A(A[6]), .ZN(n32) );
  INV_X1 U32 ( .A(B[1]), .ZN(n18) );
  INV_X1 U33 ( .A(A[1]), .ZN(n40) );
  INV_X1 U34 ( .A(B[0]), .ZN(n29) );
  INV_X1 U35 ( .A(A[0]), .ZN(n51) );
  INV_X1 U36 ( .A(A[7]), .ZN(n31) );
  INV_X1 U37 ( .A(A[8]), .ZN(n30) );
  INV_X1 U38 ( .A(A[10]), .ZN(n50) );
  INV_X1 U39 ( .A(A[11]), .ZN(n49) );
  INV_X1 U40 ( .A(A[12]), .ZN(n48) );
  INV_X1 U41 ( .A(A[13]), .ZN(n47) );
  INV_X1 U42 ( .A(A[14]), .ZN(n46) );
  INV_X1 U43 ( .A(A[9]), .ZN(n6) );
  INV_X1 U44 ( .A(A[22]), .ZN(n37) );
  INV_X1 U45 ( .A(A[15]), .ZN(n45) );
  INV_X1 U46 ( .A(A[16]), .ZN(n44) );
  INV_X1 U47 ( .A(A[17]), .ZN(n43) );
  INV_X1 U48 ( .A(A[18]), .ZN(n42) );
  INV_X1 U49 ( .A(A[19]), .ZN(n41) );
  INV_X1 U50 ( .A(A[20]), .ZN(n39) );
  INV_X1 U51 ( .A(A[21]), .ZN(n38) );
  AND2_X1 U52 ( .A1(SUMB_23__23_), .A2(CARRYB_23__22_), .ZN(A2_45_) );
  XOR2_X1 U53 ( .A(CARRYB_23__22_), .B(SUMB_23__23_), .Z(A1_44_) );
  AND2_X1 U54 ( .A1(SUMB_23__22_), .A2(CARRYB_23__21_), .ZN(A2_44_) );
  XOR2_X1 U55 ( .A(CARRYB_23__21_), .B(SUMB_23__22_), .Z(A1_43_) );
  AND2_X1 U56 ( .A1(SUMB_23__21_), .A2(CARRYB_23__20_), .ZN(A2_43_) );
  XOR2_X1 U57 ( .A(CARRYB_23__20_), .B(SUMB_23__21_), .Z(A1_42_) );
  AND2_X1 U58 ( .A1(SUMB_23__20_), .A2(CARRYB_23__19_), .ZN(A2_42_) );
  XOR2_X1 U59 ( .A(CARRYB_23__19_), .B(SUMB_23__20_), .Z(A1_41_) );
  AND2_X1 U60 ( .A1(SUMB_23__19_), .A2(CARRYB_23__18_), .ZN(A2_41_) );
  XOR2_X1 U61 ( .A(CARRYB_23__18_), .B(SUMB_23__19_), .Z(A1_40_) );
  AND2_X1 U62 ( .A1(SUMB_23__18_), .A2(CARRYB_23__17_), .ZN(A2_40_) );
  XOR2_X1 U63 ( .A(CARRYB_23__17_), .B(SUMB_23__18_), .Z(A1_39_) );
  AND2_X1 U64 ( .A1(SUMB_23__17_), .A2(CARRYB_23__16_), .ZN(A2_39_) );
  XOR2_X1 U65 ( .A(CARRYB_23__16_), .B(SUMB_23__17_), .Z(A1_38_) );
  AND2_X1 U66 ( .A1(SUMB_23__16_), .A2(CARRYB_23__15_), .ZN(A2_38_) );
  XOR2_X1 U67 ( .A(CARRYB_23__15_), .B(SUMB_23__16_), .Z(A1_37_) );
  AND2_X1 U68 ( .A1(SUMB_23__15_), .A2(CARRYB_23__14_), .ZN(A2_37_) );
  XOR2_X1 U69 ( .A(CARRYB_23__14_), .B(SUMB_23__15_), .Z(A1_36_) );
  AND2_X1 U70 ( .A1(SUMB_23__14_), .A2(CARRYB_23__13_), .ZN(A2_36_) );
  XOR2_X1 U71 ( .A(CARRYB_23__13_), .B(SUMB_23__14_), .Z(A1_35_) );
  AND2_X1 U72 ( .A1(SUMB_23__13_), .A2(CARRYB_23__12_), .ZN(A2_35_) );
  XOR2_X1 U73 ( .A(CARRYB_23__12_), .B(SUMB_23__13_), .Z(A1_34_) );
  AND2_X1 U74 ( .A1(SUMB_23__12_), .A2(CARRYB_23__11_), .ZN(A2_34_) );
  XOR2_X1 U75 ( .A(CARRYB_23__11_), .B(SUMB_23__12_), .Z(A1_33_) );
  AND2_X1 U76 ( .A1(SUMB_23__11_), .A2(CARRYB_23__10_), .ZN(A2_33_) );
  XOR2_X1 U77 ( .A(CARRYB_23__10_), .B(SUMB_23__11_), .Z(A1_32_) );
  AND2_X1 U78 ( .A1(SUMB_23__10_), .A2(CARRYB_23__9_), .ZN(A2_32_) );
  XOR2_X1 U79 ( .A(CARRYB_23__9_), .B(SUMB_23__10_), .Z(A1_31_) );
  AND2_X1 U80 ( .A1(SUMB_23__9_), .A2(CARRYB_23__8_), .ZN(A2_31_) );
  XOR2_X1 U81 ( .A(CARRYB_23__8_), .B(SUMB_23__9_), .Z(A1_30_) );
  AND2_X1 U82 ( .A1(SUMB_23__8_), .A2(CARRYB_23__7_), .ZN(A2_30_) );
  XOR2_X1 U83 ( .A(CARRYB_23__7_), .B(SUMB_23__8_), .Z(A1_29_) );
  AND2_X1 U84 ( .A1(SUMB_23__7_), .A2(CARRYB_23__6_), .ZN(A2_29_) );
  XOR2_X1 U85 ( .A(CARRYB_23__6_), .B(SUMB_23__7_), .Z(A1_28_) );
  AND2_X1 U86 ( .A1(SUMB_23__6_), .A2(CARRYB_23__5_), .ZN(A2_28_) );
  XOR2_X1 U87 ( .A(CARRYB_23__5_), .B(SUMB_23__6_), .Z(A1_27_) );
  AND2_X1 U88 ( .A1(SUMB_23__5_), .A2(CARRYB_23__4_), .ZN(A2_27_) );
  XOR2_X1 U89 ( .A(CARRYB_23__4_), .B(SUMB_23__5_), .Z(A1_26_) );
  AND2_X1 U90 ( .A1(SUMB_23__4_), .A2(CARRYB_23__3_), .ZN(A2_26_) );
  XOR2_X1 U91 ( .A(CARRYB_23__3_), .B(SUMB_23__4_), .Z(A1_25_) );
  AND2_X1 U92 ( .A1(SUMB_23__3_), .A2(CARRYB_23__2_), .ZN(A2_25_) );
  XOR2_X1 U93 ( .A(CARRYB_23__2_), .B(SUMB_23__3_), .Z(A1_24_) );
  AND2_X1 U94 ( .A1(SUMB_23__2_), .A2(CARRYB_23__1_), .ZN(A2_24_) );
  XOR2_X1 U95 ( .A(CARRYB_23__1_), .B(SUMB_23__2_), .Z(A1_23_) );
  AND2_X1 U96 ( .A1(SUMB_23__1_), .A2(CARRYB_23__0_), .ZN(A2_23_) );
  XOR2_X1 U97 ( .A(CARRYB_23__0_), .B(SUMB_23__1_), .Z(A1_22_) );
  AND2_X1 U98 ( .A1(ab_1__22_), .A2(ab_0__23_), .ZN(CARRYB_1__22_) );
  XOR2_X1 U99 ( .A(ab_1__22_), .B(ab_0__23_), .Z(SUMB_1__22_) );
  AND2_X1 U100 ( .A1(ab_1__21_), .A2(ab_0__22_), .ZN(CARRYB_1__21_) );
  XOR2_X1 U101 ( .A(ab_1__21_), .B(ab_0__22_), .Z(SUMB_1__21_) );
  AND2_X1 U102 ( .A1(ab_1__20_), .A2(ab_0__21_), .ZN(CARRYB_1__20_) );
  XOR2_X1 U103 ( .A(ab_1__20_), .B(ab_0__21_), .Z(SUMB_1__20_) );
  AND2_X1 U104 ( .A1(ab_1__19_), .A2(ab_0__20_), .ZN(CARRYB_1__19_) );
  XOR2_X1 U105 ( .A(ab_1__19_), .B(ab_0__20_), .Z(SUMB_1__19_) );
  AND2_X1 U106 ( .A1(ab_1__18_), .A2(ab_0__19_), .ZN(CARRYB_1__18_) );
  XOR2_X1 U107 ( .A(ab_1__18_), .B(ab_0__19_), .Z(SUMB_1__18_) );
  AND2_X1 U108 ( .A1(ab_1__17_), .A2(ab_0__18_), .ZN(CARRYB_1__17_) );
  XOR2_X1 U109 ( .A(ab_1__17_), .B(ab_0__18_), .Z(SUMB_1__17_) );
  AND2_X1 U110 ( .A1(ab_1__16_), .A2(ab_0__17_), .ZN(CARRYB_1__16_) );
  XOR2_X1 U111 ( .A(ab_1__16_), .B(ab_0__17_), .Z(SUMB_1__16_) );
  AND2_X1 U112 ( .A1(ab_1__15_), .A2(ab_0__16_), .ZN(CARRYB_1__15_) );
  XOR2_X1 U113 ( .A(ab_1__15_), .B(ab_0__16_), .Z(SUMB_1__15_) );
  AND2_X1 U114 ( .A1(ab_1__14_), .A2(ab_0__15_), .ZN(CARRYB_1__14_) );
  XOR2_X1 U115 ( .A(ab_1__14_), .B(ab_0__15_), .Z(SUMB_1__14_) );
  AND2_X1 U116 ( .A1(ab_1__13_), .A2(ab_0__14_), .ZN(CARRYB_1__13_) );
  XOR2_X1 U117 ( .A(ab_1__13_), .B(ab_0__14_), .Z(SUMB_1__13_) );
  AND2_X1 U118 ( .A1(ab_1__12_), .A2(ab_0__13_), .ZN(CARRYB_1__12_) );
  XOR2_X1 U119 ( .A(ab_1__12_), .B(ab_0__13_), .Z(SUMB_1__12_) );
  AND2_X1 U120 ( .A1(ab_1__11_), .A2(ab_0__12_), .ZN(CARRYB_1__11_) );
  XOR2_X1 U121 ( .A(ab_1__11_), .B(ab_0__12_), .Z(SUMB_1__11_) );
  AND2_X1 U122 ( .A1(ab_1__10_), .A2(ab_0__11_), .ZN(CARRYB_1__10_) );
  XOR2_X1 U123 ( .A(ab_1__10_), .B(ab_0__11_), .Z(SUMB_1__10_) );
  AND2_X1 U124 ( .A1(ab_1__9_), .A2(ab_0__10_), .ZN(CARRYB_1__9_) );
  XOR2_X1 U125 ( .A(ab_1__9_), .B(ab_0__10_), .Z(SUMB_1__9_) );
  AND2_X1 U126 ( .A1(ab_1__8_), .A2(ab_0__9_), .ZN(CARRYB_1__8_) );
  XOR2_X1 U127 ( .A(ab_1__8_), .B(ab_0__9_), .Z(SUMB_1__8_) );
  AND2_X1 U128 ( .A1(ab_1__7_), .A2(ab_0__8_), .ZN(CARRYB_1__7_) );
  XOR2_X1 U129 ( .A(ab_1__7_), .B(ab_0__8_), .Z(SUMB_1__7_) );
  AND2_X1 U130 ( .A1(ab_1__6_), .A2(ab_0__7_), .ZN(CARRYB_1__6_) );
  XOR2_X1 U131 ( .A(ab_1__6_), .B(ab_0__7_), .Z(SUMB_1__6_) );
  AND2_X1 U132 ( .A1(ab_1__5_), .A2(ab_0__6_), .ZN(CARRYB_1__5_) );
  XOR2_X1 U133 ( .A(ab_1__5_), .B(ab_0__6_), .Z(SUMB_1__5_) );
  AND2_X1 U134 ( .A1(ab_1__4_), .A2(ab_0__5_), .ZN(CARRYB_1__4_) );
  XOR2_X1 U135 ( .A(ab_1__4_), .B(ab_0__5_), .Z(SUMB_1__4_) );
  AND2_X1 U136 ( .A1(ab_1__3_), .A2(ab_0__4_), .ZN(CARRYB_1__3_) );
  XOR2_X1 U137 ( .A(ab_1__3_), .B(ab_0__4_), .Z(SUMB_1__3_) );
  AND2_X1 U138 ( .A1(ab_1__2_), .A2(ab_0__3_), .ZN(CARRYB_1__2_) );
  XOR2_X1 U139 ( .A(ab_1__2_), .B(ab_0__3_), .Z(SUMB_1__2_) );
  AND2_X1 U140 ( .A1(ab_1__1_), .A2(ab_0__2_), .ZN(CARRYB_1__1_) );
  XOR2_X1 U141 ( .A(ab_1__1_), .B(ab_0__2_), .Z(SUMB_1__1_) );
  NOR2_X1 U142 ( .A1(n6), .A2(n7), .ZN(ab_9__9_) );
  NOR2_X1 U143 ( .A1(n6), .A2(n8), .ZN(ab_9__8_) );
  NOR2_X1 U144 ( .A1(n6), .A2(n9), .ZN(ab_9__7_) );
  NOR2_X1 U145 ( .A1(n6), .A2(n10), .ZN(ab_9__6_) );
  NOR2_X1 U146 ( .A1(n6), .A2(n11), .ZN(ab_9__5_) );
  NOR2_X1 U147 ( .A1(n6), .A2(n12), .ZN(ab_9__4_) );
  NOR2_X1 U148 ( .A1(n6), .A2(n13), .ZN(ab_9__3_) );
  NOR2_X1 U149 ( .A1(n6), .A2(n14), .ZN(ab_9__2_) );
  NOR2_X1 U150 ( .A1(A[9]), .A2(n1), .ZN(ab_9__23_) );
  NOR2_X1 U151 ( .A1(n6), .A2(n15), .ZN(ab_9__22_) );
  NOR2_X1 U152 ( .A1(n6), .A2(n16), .ZN(ab_9__21_) );
  NOR2_X1 U153 ( .A1(n6), .A2(n17), .ZN(ab_9__20_) );
  NOR2_X1 U154 ( .A1(n6), .A2(n18), .ZN(ab_9__1_) );
  NOR2_X1 U155 ( .A1(n6), .A2(n19), .ZN(ab_9__19_) );
  NOR2_X1 U156 ( .A1(n6), .A2(n20), .ZN(ab_9__18_) );
  NOR2_X1 U157 ( .A1(n6), .A2(n21), .ZN(ab_9__17_) );
  NOR2_X1 U158 ( .A1(n6), .A2(n22), .ZN(ab_9__16_) );
  NOR2_X1 U159 ( .A1(n6), .A2(n23), .ZN(ab_9__15_) );
  NOR2_X1 U160 ( .A1(n6), .A2(n24), .ZN(ab_9__14_) );
  NOR2_X1 U161 ( .A1(n6), .A2(n25), .ZN(ab_9__13_) );
  NOR2_X1 U162 ( .A1(n6), .A2(n26), .ZN(ab_9__12_) );
  NOR2_X1 U163 ( .A1(n6), .A2(n27), .ZN(ab_9__11_) );
  NOR2_X1 U164 ( .A1(n6), .A2(n28), .ZN(ab_9__10_) );
  NOR2_X1 U165 ( .A1(n6), .A2(n29), .ZN(ab_9__0_) );
  NOR2_X1 U166 ( .A1(n7), .A2(n30), .ZN(ab_8__9_) );
  NOR2_X1 U167 ( .A1(n8), .A2(n30), .ZN(ab_8__8_) );
  NOR2_X1 U168 ( .A1(n9), .A2(n30), .ZN(ab_8__7_) );
  NOR2_X1 U169 ( .A1(n10), .A2(n30), .ZN(ab_8__6_) );
  NOR2_X1 U170 ( .A1(n11), .A2(n30), .ZN(ab_8__5_) );
  NOR2_X1 U171 ( .A1(n12), .A2(n30), .ZN(ab_8__4_) );
  NOR2_X1 U172 ( .A1(n13), .A2(n30), .ZN(ab_8__3_) );
  NOR2_X1 U173 ( .A1(n14), .A2(n30), .ZN(ab_8__2_) );
  NOR2_X1 U174 ( .A1(A[8]), .A2(n1), .ZN(ab_8__23_) );
  NOR2_X1 U175 ( .A1(n15), .A2(n30), .ZN(ab_8__22_) );
  NOR2_X1 U176 ( .A1(n16), .A2(n30), .ZN(ab_8__21_) );
  NOR2_X1 U177 ( .A1(n17), .A2(n30), .ZN(ab_8__20_) );
  NOR2_X1 U178 ( .A1(n18), .A2(n30), .ZN(ab_8__1_) );
  NOR2_X1 U179 ( .A1(n19), .A2(n30), .ZN(ab_8__19_) );
  NOR2_X1 U180 ( .A1(n20), .A2(n30), .ZN(ab_8__18_) );
  NOR2_X1 U181 ( .A1(n21), .A2(n30), .ZN(ab_8__17_) );
  NOR2_X1 U182 ( .A1(n22), .A2(n30), .ZN(ab_8__16_) );
  NOR2_X1 U183 ( .A1(n23), .A2(n30), .ZN(ab_8__15_) );
  NOR2_X1 U184 ( .A1(n24), .A2(n30), .ZN(ab_8__14_) );
  NOR2_X1 U185 ( .A1(n25), .A2(n30), .ZN(ab_8__13_) );
  NOR2_X1 U186 ( .A1(n26), .A2(n30), .ZN(ab_8__12_) );
  NOR2_X1 U187 ( .A1(n27), .A2(n30), .ZN(ab_8__11_) );
  NOR2_X1 U188 ( .A1(n28), .A2(n30), .ZN(ab_8__10_) );
  NOR2_X1 U189 ( .A1(n29), .A2(n30), .ZN(ab_8__0_) );
  NOR2_X1 U190 ( .A1(n7), .A2(n31), .ZN(ab_7__9_) );
  NOR2_X1 U191 ( .A1(n8), .A2(n31), .ZN(ab_7__8_) );
  NOR2_X1 U192 ( .A1(n9), .A2(n31), .ZN(ab_7__7_) );
  NOR2_X1 U193 ( .A1(n10), .A2(n31), .ZN(ab_7__6_) );
  NOR2_X1 U194 ( .A1(n11), .A2(n31), .ZN(ab_7__5_) );
  NOR2_X1 U195 ( .A1(n12), .A2(n31), .ZN(ab_7__4_) );
  NOR2_X1 U196 ( .A1(n13), .A2(n31), .ZN(ab_7__3_) );
  NOR2_X1 U197 ( .A1(n14), .A2(n31), .ZN(ab_7__2_) );
  NOR2_X1 U198 ( .A1(A[7]), .A2(n1), .ZN(ab_7__23_) );
  NOR2_X1 U199 ( .A1(n15), .A2(n31), .ZN(ab_7__22_) );
  NOR2_X1 U200 ( .A1(n16), .A2(n31), .ZN(ab_7__21_) );
  NOR2_X1 U201 ( .A1(n17), .A2(n31), .ZN(ab_7__20_) );
  NOR2_X1 U202 ( .A1(n18), .A2(n31), .ZN(ab_7__1_) );
  NOR2_X1 U203 ( .A1(n19), .A2(n31), .ZN(ab_7__19_) );
  NOR2_X1 U204 ( .A1(n20), .A2(n31), .ZN(ab_7__18_) );
  NOR2_X1 U205 ( .A1(n21), .A2(n31), .ZN(ab_7__17_) );
  NOR2_X1 U206 ( .A1(n22), .A2(n31), .ZN(ab_7__16_) );
  NOR2_X1 U207 ( .A1(n23), .A2(n31), .ZN(ab_7__15_) );
  NOR2_X1 U208 ( .A1(n24), .A2(n31), .ZN(ab_7__14_) );
  NOR2_X1 U209 ( .A1(n25), .A2(n31), .ZN(ab_7__13_) );
  NOR2_X1 U210 ( .A1(n26), .A2(n31), .ZN(ab_7__12_) );
  NOR2_X1 U211 ( .A1(n27), .A2(n31), .ZN(ab_7__11_) );
  NOR2_X1 U212 ( .A1(n28), .A2(n31), .ZN(ab_7__10_) );
  NOR2_X1 U213 ( .A1(n29), .A2(n31), .ZN(ab_7__0_) );
  NOR2_X1 U214 ( .A1(n7), .A2(n32), .ZN(ab_6__9_) );
  NOR2_X1 U215 ( .A1(n8), .A2(n32), .ZN(ab_6__8_) );
  NOR2_X1 U216 ( .A1(n9), .A2(n32), .ZN(ab_6__7_) );
  NOR2_X1 U217 ( .A1(n10), .A2(n32), .ZN(ab_6__6_) );
  NOR2_X1 U218 ( .A1(n11), .A2(n32), .ZN(ab_6__5_) );
  NOR2_X1 U219 ( .A1(n12), .A2(n32), .ZN(ab_6__4_) );
  NOR2_X1 U220 ( .A1(n13), .A2(n32), .ZN(ab_6__3_) );
  NOR2_X1 U221 ( .A1(n14), .A2(n32), .ZN(ab_6__2_) );
  NOR2_X1 U222 ( .A1(A[6]), .A2(n1), .ZN(ab_6__23_) );
  NOR2_X1 U223 ( .A1(n15), .A2(n32), .ZN(ab_6__22_) );
  NOR2_X1 U224 ( .A1(n16), .A2(n32), .ZN(ab_6__21_) );
  NOR2_X1 U225 ( .A1(n17), .A2(n32), .ZN(ab_6__20_) );
  NOR2_X1 U226 ( .A1(n18), .A2(n32), .ZN(ab_6__1_) );
  NOR2_X1 U227 ( .A1(n19), .A2(n32), .ZN(ab_6__19_) );
  NOR2_X1 U228 ( .A1(n20), .A2(n32), .ZN(ab_6__18_) );
  NOR2_X1 U229 ( .A1(n21), .A2(n32), .ZN(ab_6__17_) );
  NOR2_X1 U230 ( .A1(n22), .A2(n32), .ZN(ab_6__16_) );
  NOR2_X1 U231 ( .A1(n23), .A2(n32), .ZN(ab_6__15_) );
  NOR2_X1 U232 ( .A1(n24), .A2(n32), .ZN(ab_6__14_) );
  NOR2_X1 U233 ( .A1(n25), .A2(n32), .ZN(ab_6__13_) );
  NOR2_X1 U234 ( .A1(n26), .A2(n32), .ZN(ab_6__12_) );
  NOR2_X1 U235 ( .A1(n27), .A2(n32), .ZN(ab_6__11_) );
  NOR2_X1 U236 ( .A1(n28), .A2(n32), .ZN(ab_6__10_) );
  NOR2_X1 U237 ( .A1(n29), .A2(n32), .ZN(ab_6__0_) );
  NOR2_X1 U238 ( .A1(n7), .A2(n33), .ZN(ab_5__9_) );
  NOR2_X1 U239 ( .A1(n8), .A2(n33), .ZN(ab_5__8_) );
  NOR2_X1 U240 ( .A1(n9), .A2(n33), .ZN(ab_5__7_) );
  NOR2_X1 U241 ( .A1(n10), .A2(n33), .ZN(ab_5__6_) );
  NOR2_X1 U242 ( .A1(n11), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U243 ( .A1(n12), .A2(n33), .ZN(ab_5__4_) );
  NOR2_X1 U244 ( .A1(n13), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U245 ( .A1(n14), .A2(n33), .ZN(ab_5__2_) );
  NOR2_X1 U246 ( .A1(A[5]), .A2(n1), .ZN(ab_5__23_) );
  NOR2_X1 U247 ( .A1(n15), .A2(n33), .ZN(ab_5__22_) );
  NOR2_X1 U248 ( .A1(n16), .A2(n33), .ZN(ab_5__21_) );
  NOR2_X1 U249 ( .A1(n17), .A2(n33), .ZN(ab_5__20_) );
  NOR2_X1 U250 ( .A1(n18), .A2(n33), .ZN(ab_5__1_) );
  NOR2_X1 U251 ( .A1(n19), .A2(n33), .ZN(ab_5__19_) );
  NOR2_X1 U252 ( .A1(n20), .A2(n33), .ZN(ab_5__18_) );
  NOR2_X1 U253 ( .A1(n21), .A2(n33), .ZN(ab_5__17_) );
  NOR2_X1 U254 ( .A1(n22), .A2(n33), .ZN(ab_5__16_) );
  NOR2_X1 U255 ( .A1(n23), .A2(n33), .ZN(ab_5__15_) );
  NOR2_X1 U256 ( .A1(n24), .A2(n33), .ZN(ab_5__14_) );
  NOR2_X1 U257 ( .A1(n25), .A2(n33), .ZN(ab_5__13_) );
  NOR2_X1 U258 ( .A1(n26), .A2(n33), .ZN(ab_5__12_) );
  NOR2_X1 U259 ( .A1(n27), .A2(n33), .ZN(ab_5__11_) );
  NOR2_X1 U260 ( .A1(n28), .A2(n33), .ZN(ab_5__10_) );
  NOR2_X1 U261 ( .A1(n29), .A2(n33), .ZN(ab_5__0_) );
  NOR2_X1 U262 ( .A1(n7), .A2(n34), .ZN(ab_4__9_) );
  NOR2_X1 U263 ( .A1(n8), .A2(n34), .ZN(ab_4__8_) );
  NOR2_X1 U264 ( .A1(n9), .A2(n34), .ZN(ab_4__7_) );
  NOR2_X1 U265 ( .A1(n10), .A2(n34), .ZN(ab_4__6_) );
  NOR2_X1 U266 ( .A1(n11), .A2(n34), .ZN(ab_4__5_) );
  NOR2_X1 U267 ( .A1(n12), .A2(n34), .ZN(ab_4__4_) );
  NOR2_X1 U268 ( .A1(n13), .A2(n34), .ZN(ab_4__3_) );
  NOR2_X1 U269 ( .A1(n14), .A2(n34), .ZN(ab_4__2_) );
  NOR2_X1 U270 ( .A1(A[4]), .A2(n1), .ZN(ab_4__23_) );
  NOR2_X1 U271 ( .A1(n15), .A2(n34), .ZN(ab_4__22_) );
  NOR2_X1 U272 ( .A1(n16), .A2(n34), .ZN(ab_4__21_) );
  NOR2_X1 U273 ( .A1(n17), .A2(n34), .ZN(ab_4__20_) );
  NOR2_X1 U274 ( .A1(n18), .A2(n34), .ZN(ab_4__1_) );
  NOR2_X1 U275 ( .A1(n19), .A2(n34), .ZN(ab_4__19_) );
  NOR2_X1 U276 ( .A1(n20), .A2(n34), .ZN(ab_4__18_) );
  NOR2_X1 U277 ( .A1(n21), .A2(n34), .ZN(ab_4__17_) );
  NOR2_X1 U278 ( .A1(n22), .A2(n34), .ZN(ab_4__16_) );
  NOR2_X1 U279 ( .A1(n23), .A2(n34), .ZN(ab_4__15_) );
  NOR2_X1 U280 ( .A1(n24), .A2(n34), .ZN(ab_4__14_) );
  NOR2_X1 U281 ( .A1(n25), .A2(n34), .ZN(ab_4__13_) );
  NOR2_X1 U282 ( .A1(n26), .A2(n34), .ZN(ab_4__12_) );
  NOR2_X1 U283 ( .A1(n27), .A2(n34), .ZN(ab_4__11_) );
  NOR2_X1 U284 ( .A1(n28), .A2(n34), .ZN(ab_4__10_) );
  NOR2_X1 U285 ( .A1(n29), .A2(n34), .ZN(ab_4__0_) );
  NOR2_X1 U286 ( .A1(n7), .A2(n35), .ZN(ab_3__9_) );
  NOR2_X1 U287 ( .A1(n8), .A2(n35), .ZN(ab_3__8_) );
  NOR2_X1 U288 ( .A1(n9), .A2(n35), .ZN(ab_3__7_) );
  NOR2_X1 U289 ( .A1(n10), .A2(n35), .ZN(ab_3__6_) );
  NOR2_X1 U290 ( .A1(n11), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U291 ( .A1(n12), .A2(n35), .ZN(ab_3__4_) );
  NOR2_X1 U292 ( .A1(n13), .A2(n35), .ZN(ab_3__3_) );
  NOR2_X1 U293 ( .A1(n14), .A2(n35), .ZN(ab_3__2_) );
  NOR2_X1 U294 ( .A1(A[3]), .A2(n1), .ZN(ab_3__23_) );
  NOR2_X1 U295 ( .A1(n15), .A2(n35), .ZN(ab_3__22_) );
  NOR2_X1 U296 ( .A1(n16), .A2(n35), .ZN(ab_3__21_) );
  NOR2_X1 U297 ( .A1(n17), .A2(n35), .ZN(ab_3__20_) );
  NOR2_X1 U298 ( .A1(n18), .A2(n35), .ZN(ab_3__1_) );
  NOR2_X1 U299 ( .A1(n19), .A2(n35), .ZN(ab_3__19_) );
  NOR2_X1 U300 ( .A1(n20), .A2(n35), .ZN(ab_3__18_) );
  NOR2_X1 U301 ( .A1(n21), .A2(n35), .ZN(ab_3__17_) );
  NOR2_X1 U302 ( .A1(n22), .A2(n35), .ZN(ab_3__16_) );
  NOR2_X1 U303 ( .A1(n23), .A2(n35), .ZN(ab_3__15_) );
  NOR2_X1 U304 ( .A1(n24), .A2(n35), .ZN(ab_3__14_) );
  NOR2_X1 U305 ( .A1(n25), .A2(n35), .ZN(ab_3__13_) );
  NOR2_X1 U306 ( .A1(n26), .A2(n35), .ZN(ab_3__12_) );
  NOR2_X1 U307 ( .A1(n27), .A2(n35), .ZN(ab_3__11_) );
  NOR2_X1 U308 ( .A1(n28), .A2(n35), .ZN(ab_3__10_) );
  NOR2_X1 U309 ( .A1(n29), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U310 ( .A1(n7), .A2(n36), .ZN(ab_2__9_) );
  NOR2_X1 U311 ( .A1(n8), .A2(n36), .ZN(ab_2__8_) );
  NOR2_X1 U312 ( .A1(n9), .A2(n36), .ZN(ab_2__7_) );
  NOR2_X1 U313 ( .A1(n10), .A2(n36), .ZN(ab_2__6_) );
  NOR2_X1 U314 ( .A1(n11), .A2(n36), .ZN(ab_2__5_) );
  NOR2_X1 U315 ( .A1(n12), .A2(n36), .ZN(ab_2__4_) );
  NOR2_X1 U316 ( .A1(n13), .A2(n36), .ZN(ab_2__3_) );
  NOR2_X1 U317 ( .A1(n14), .A2(n36), .ZN(ab_2__2_) );
  NOR2_X1 U318 ( .A1(A[2]), .A2(n1), .ZN(ab_2__23_) );
  NOR2_X1 U319 ( .A1(n15), .A2(n36), .ZN(ab_2__22_) );
  NOR2_X1 U320 ( .A1(n16), .A2(n36), .ZN(ab_2__21_) );
  NOR2_X1 U321 ( .A1(n17), .A2(n36), .ZN(ab_2__20_) );
  NOR2_X1 U322 ( .A1(n18), .A2(n36), .ZN(ab_2__1_) );
  NOR2_X1 U323 ( .A1(n19), .A2(n36), .ZN(ab_2__19_) );
  NOR2_X1 U324 ( .A1(n20), .A2(n36), .ZN(ab_2__18_) );
  NOR2_X1 U325 ( .A1(n21), .A2(n36), .ZN(ab_2__17_) );
  NOR2_X1 U326 ( .A1(n22), .A2(n36), .ZN(ab_2__16_) );
  NOR2_X1 U327 ( .A1(n23), .A2(n36), .ZN(ab_2__15_) );
  NOR2_X1 U328 ( .A1(n24), .A2(n36), .ZN(ab_2__14_) );
  NOR2_X1 U329 ( .A1(n25), .A2(n36), .ZN(ab_2__13_) );
  NOR2_X1 U330 ( .A1(n26), .A2(n36), .ZN(ab_2__12_) );
  NOR2_X1 U331 ( .A1(n27), .A2(n36), .ZN(ab_2__11_) );
  NOR2_X1 U332 ( .A1(n28), .A2(n36), .ZN(ab_2__10_) );
  NOR2_X1 U333 ( .A1(n29), .A2(n36), .ZN(ab_2__0_) );
  NOR2_X1 U334 ( .A1(B[9]), .A2(n4), .ZN(ab_23__9_) );
  NOR2_X1 U335 ( .A1(B[8]), .A2(n4), .ZN(ab_23__8_) );
  NOR2_X1 U336 ( .A1(B[7]), .A2(n4), .ZN(ab_23__7_) );
  NOR2_X1 U337 ( .A1(B[6]), .A2(n4), .ZN(ab_23__6_) );
  NOR2_X1 U338 ( .A1(B[5]), .A2(n3), .ZN(ab_23__5_) );
  NOR2_X1 U339 ( .A1(B[4]), .A2(n3), .ZN(ab_23__4_) );
  NOR2_X1 U340 ( .A1(B[3]), .A2(n3), .ZN(ab_23__3_) );
  NOR2_X1 U341 ( .A1(B[2]), .A2(n3), .ZN(ab_23__2_) );
  NOR2_X1 U342 ( .A1(n1), .A2(n3), .ZN(ab_23__23_) );
  NOR2_X1 U343 ( .A1(B[22]), .A2(n3), .ZN(ab_23__22_) );
  NOR2_X1 U344 ( .A1(B[21]), .A2(n3), .ZN(ab_23__21_) );
  NOR2_X1 U345 ( .A1(B[20]), .A2(n3), .ZN(ab_23__20_) );
  NOR2_X1 U346 ( .A1(B[1]), .A2(n3), .ZN(ab_23__1_) );
  NOR2_X1 U347 ( .A1(B[19]), .A2(n3), .ZN(ab_23__19_) );
  NOR2_X1 U348 ( .A1(B[18]), .A2(n3), .ZN(ab_23__18_) );
  NOR2_X1 U349 ( .A1(B[17]), .A2(n3), .ZN(ab_23__17_) );
  NOR2_X1 U350 ( .A1(B[16]), .A2(n3), .ZN(ab_23__16_) );
  NOR2_X1 U351 ( .A1(B[15]), .A2(n3), .ZN(ab_23__15_) );
  NOR2_X1 U352 ( .A1(B[14]), .A2(n3), .ZN(ab_23__14_) );
  NOR2_X1 U353 ( .A1(B[13]), .A2(n3), .ZN(ab_23__13_) );
  NOR2_X1 U354 ( .A1(B[12]), .A2(n3), .ZN(ab_23__12_) );
  NOR2_X1 U355 ( .A1(B[11]), .A2(n3), .ZN(ab_23__11_) );
  NOR2_X1 U356 ( .A1(B[10]), .A2(n3), .ZN(ab_23__10_) );
  NOR2_X1 U357 ( .A1(B[0]), .A2(n3), .ZN(ab_23__0_) );
  NOR2_X1 U358 ( .A1(n7), .A2(n37), .ZN(ab_22__9_) );
  NOR2_X1 U359 ( .A1(n8), .A2(n37), .ZN(ab_22__8_) );
  NOR2_X1 U360 ( .A1(n9), .A2(n37), .ZN(ab_22__7_) );
  NOR2_X1 U361 ( .A1(n10), .A2(n37), .ZN(ab_22__6_) );
  NOR2_X1 U362 ( .A1(n11), .A2(n37), .ZN(ab_22__5_) );
  NOR2_X1 U363 ( .A1(n12), .A2(n37), .ZN(ab_22__4_) );
  NOR2_X1 U364 ( .A1(n13), .A2(n37), .ZN(ab_22__3_) );
  NOR2_X1 U365 ( .A1(n14), .A2(n37), .ZN(ab_22__2_) );
  NOR2_X1 U366 ( .A1(A[22]), .A2(n1), .ZN(ab_22__23_) );
  NOR2_X1 U367 ( .A1(n15), .A2(n37), .ZN(ab_22__22_) );
  NOR2_X1 U368 ( .A1(n16), .A2(n37), .ZN(ab_22__21_) );
  NOR2_X1 U369 ( .A1(n17), .A2(n37), .ZN(ab_22__20_) );
  NOR2_X1 U370 ( .A1(n18), .A2(n37), .ZN(ab_22__1_) );
  NOR2_X1 U371 ( .A1(n19), .A2(n37), .ZN(ab_22__19_) );
  NOR2_X1 U372 ( .A1(n20), .A2(n37), .ZN(ab_22__18_) );
  NOR2_X1 U373 ( .A1(n21), .A2(n37), .ZN(ab_22__17_) );
  NOR2_X1 U374 ( .A1(n22), .A2(n37), .ZN(ab_22__16_) );
  NOR2_X1 U375 ( .A1(n23), .A2(n37), .ZN(ab_22__15_) );
  NOR2_X1 U376 ( .A1(n24), .A2(n37), .ZN(ab_22__14_) );
  NOR2_X1 U377 ( .A1(n25), .A2(n37), .ZN(ab_22__13_) );
  NOR2_X1 U378 ( .A1(n26), .A2(n37), .ZN(ab_22__12_) );
  NOR2_X1 U379 ( .A1(n27), .A2(n37), .ZN(ab_22__11_) );
  NOR2_X1 U380 ( .A1(n28), .A2(n37), .ZN(ab_22__10_) );
  NOR2_X1 U381 ( .A1(n29), .A2(n37), .ZN(ab_22__0_) );
  NOR2_X1 U382 ( .A1(n7), .A2(n38), .ZN(ab_21__9_) );
  NOR2_X1 U383 ( .A1(n8), .A2(n38), .ZN(ab_21__8_) );
  NOR2_X1 U384 ( .A1(n9), .A2(n38), .ZN(ab_21__7_) );
  NOR2_X1 U385 ( .A1(n10), .A2(n38), .ZN(ab_21__6_) );
  NOR2_X1 U386 ( .A1(n11), .A2(n38), .ZN(ab_21__5_) );
  NOR2_X1 U387 ( .A1(n12), .A2(n38), .ZN(ab_21__4_) );
  NOR2_X1 U388 ( .A1(n13), .A2(n38), .ZN(ab_21__3_) );
  NOR2_X1 U389 ( .A1(n14), .A2(n38), .ZN(ab_21__2_) );
  NOR2_X1 U390 ( .A1(A[21]), .A2(n1), .ZN(ab_21__23_) );
  NOR2_X1 U391 ( .A1(n15), .A2(n38), .ZN(ab_21__22_) );
  NOR2_X1 U392 ( .A1(n16), .A2(n38), .ZN(ab_21__21_) );
  NOR2_X1 U393 ( .A1(n17), .A2(n38), .ZN(ab_21__20_) );
  NOR2_X1 U394 ( .A1(n18), .A2(n38), .ZN(ab_21__1_) );
  NOR2_X1 U395 ( .A1(n19), .A2(n38), .ZN(ab_21__19_) );
  NOR2_X1 U396 ( .A1(n20), .A2(n38), .ZN(ab_21__18_) );
  NOR2_X1 U397 ( .A1(n21), .A2(n38), .ZN(ab_21__17_) );
  NOR2_X1 U398 ( .A1(n22), .A2(n38), .ZN(ab_21__16_) );
  NOR2_X1 U399 ( .A1(n23), .A2(n38), .ZN(ab_21__15_) );
  NOR2_X1 U400 ( .A1(n24), .A2(n38), .ZN(ab_21__14_) );
  NOR2_X1 U401 ( .A1(n25), .A2(n38), .ZN(ab_21__13_) );
  NOR2_X1 U402 ( .A1(n26), .A2(n38), .ZN(ab_21__12_) );
  NOR2_X1 U403 ( .A1(n27), .A2(n38), .ZN(ab_21__11_) );
  NOR2_X1 U404 ( .A1(n28), .A2(n38), .ZN(ab_21__10_) );
  NOR2_X1 U405 ( .A1(n29), .A2(n38), .ZN(ab_21__0_) );
  NOR2_X1 U406 ( .A1(n7), .A2(n39), .ZN(ab_20__9_) );
  NOR2_X1 U407 ( .A1(n8), .A2(n39), .ZN(ab_20__8_) );
  NOR2_X1 U408 ( .A1(n9), .A2(n39), .ZN(ab_20__7_) );
  NOR2_X1 U409 ( .A1(n10), .A2(n39), .ZN(ab_20__6_) );
  NOR2_X1 U410 ( .A1(n11), .A2(n39), .ZN(ab_20__5_) );
  NOR2_X1 U411 ( .A1(n12), .A2(n39), .ZN(ab_20__4_) );
  NOR2_X1 U412 ( .A1(n13), .A2(n39), .ZN(ab_20__3_) );
  NOR2_X1 U413 ( .A1(n14), .A2(n39), .ZN(ab_20__2_) );
  NOR2_X1 U414 ( .A1(A[20]), .A2(n1), .ZN(ab_20__23_) );
  NOR2_X1 U415 ( .A1(n15), .A2(n39), .ZN(ab_20__22_) );
  NOR2_X1 U416 ( .A1(n16), .A2(n39), .ZN(ab_20__21_) );
  NOR2_X1 U417 ( .A1(n17), .A2(n39), .ZN(ab_20__20_) );
  NOR2_X1 U418 ( .A1(n18), .A2(n39), .ZN(ab_20__1_) );
  NOR2_X1 U419 ( .A1(n19), .A2(n39), .ZN(ab_20__19_) );
  NOR2_X1 U420 ( .A1(n20), .A2(n39), .ZN(ab_20__18_) );
  NOR2_X1 U421 ( .A1(n21), .A2(n39), .ZN(ab_20__17_) );
  NOR2_X1 U422 ( .A1(n22), .A2(n39), .ZN(ab_20__16_) );
  NOR2_X1 U423 ( .A1(n23), .A2(n39), .ZN(ab_20__15_) );
  NOR2_X1 U424 ( .A1(n24), .A2(n39), .ZN(ab_20__14_) );
  NOR2_X1 U425 ( .A1(n25), .A2(n39), .ZN(ab_20__13_) );
  NOR2_X1 U426 ( .A1(n26), .A2(n39), .ZN(ab_20__12_) );
  NOR2_X1 U427 ( .A1(n27), .A2(n39), .ZN(ab_20__11_) );
  NOR2_X1 U428 ( .A1(n28), .A2(n39), .ZN(ab_20__10_) );
  NOR2_X1 U429 ( .A1(n29), .A2(n39), .ZN(ab_20__0_) );
  NOR2_X1 U430 ( .A1(n7), .A2(n40), .ZN(ab_1__9_) );
  NOR2_X1 U431 ( .A1(n8), .A2(n40), .ZN(ab_1__8_) );
  NOR2_X1 U432 ( .A1(n9), .A2(n40), .ZN(ab_1__7_) );
  NOR2_X1 U433 ( .A1(n10), .A2(n40), .ZN(ab_1__6_) );
  NOR2_X1 U434 ( .A1(n11), .A2(n40), .ZN(ab_1__5_) );
  NOR2_X1 U435 ( .A1(n12), .A2(n40), .ZN(ab_1__4_) );
  NOR2_X1 U436 ( .A1(n13), .A2(n40), .ZN(ab_1__3_) );
  NOR2_X1 U437 ( .A1(n14), .A2(n40), .ZN(ab_1__2_) );
  NOR2_X1 U438 ( .A1(A[1]), .A2(n1), .ZN(ab_1__23_) );
  NOR2_X1 U439 ( .A1(n15), .A2(n40), .ZN(ab_1__22_) );
  NOR2_X1 U440 ( .A1(n16), .A2(n40), .ZN(ab_1__21_) );
  NOR2_X1 U441 ( .A1(n17), .A2(n40), .ZN(ab_1__20_) );
  NOR2_X1 U442 ( .A1(n19), .A2(n40), .ZN(ab_1__19_) );
  NOR2_X1 U443 ( .A1(n20), .A2(n40), .ZN(ab_1__18_) );
  NOR2_X1 U444 ( .A1(n21), .A2(n40), .ZN(ab_1__17_) );
  NOR2_X1 U445 ( .A1(n22), .A2(n40), .ZN(ab_1__16_) );
  NOR2_X1 U446 ( .A1(n23), .A2(n40), .ZN(ab_1__15_) );
  NOR2_X1 U447 ( .A1(n24), .A2(n40), .ZN(ab_1__14_) );
  NOR2_X1 U448 ( .A1(n25), .A2(n40), .ZN(ab_1__13_) );
  NOR2_X1 U449 ( .A1(n26), .A2(n40), .ZN(ab_1__12_) );
  NOR2_X1 U450 ( .A1(n27), .A2(n40), .ZN(ab_1__11_) );
  NOR2_X1 U451 ( .A1(n28), .A2(n40), .ZN(ab_1__10_) );
  NOR2_X1 U452 ( .A1(n7), .A2(n41), .ZN(ab_19__9_) );
  NOR2_X1 U453 ( .A1(n8), .A2(n41), .ZN(ab_19__8_) );
  NOR2_X1 U454 ( .A1(n9), .A2(n41), .ZN(ab_19__7_) );
  NOR2_X1 U455 ( .A1(n10), .A2(n41), .ZN(ab_19__6_) );
  NOR2_X1 U456 ( .A1(n11), .A2(n41), .ZN(ab_19__5_) );
  NOR2_X1 U457 ( .A1(n12), .A2(n41), .ZN(ab_19__4_) );
  NOR2_X1 U458 ( .A1(n13), .A2(n41), .ZN(ab_19__3_) );
  NOR2_X1 U459 ( .A1(n14), .A2(n41), .ZN(ab_19__2_) );
  NOR2_X1 U460 ( .A1(A[19]), .A2(n1), .ZN(ab_19__23_) );
  NOR2_X1 U461 ( .A1(n15), .A2(n41), .ZN(ab_19__22_) );
  NOR2_X1 U462 ( .A1(n16), .A2(n41), .ZN(ab_19__21_) );
  NOR2_X1 U463 ( .A1(n17), .A2(n41), .ZN(ab_19__20_) );
  NOR2_X1 U464 ( .A1(n18), .A2(n41), .ZN(ab_19__1_) );
  NOR2_X1 U465 ( .A1(n19), .A2(n41), .ZN(ab_19__19_) );
  NOR2_X1 U466 ( .A1(n20), .A2(n41), .ZN(ab_19__18_) );
  NOR2_X1 U467 ( .A1(n21), .A2(n41), .ZN(ab_19__17_) );
  NOR2_X1 U468 ( .A1(n22), .A2(n41), .ZN(ab_19__16_) );
  NOR2_X1 U469 ( .A1(n23), .A2(n41), .ZN(ab_19__15_) );
  NOR2_X1 U470 ( .A1(n24), .A2(n41), .ZN(ab_19__14_) );
  NOR2_X1 U471 ( .A1(n25), .A2(n41), .ZN(ab_19__13_) );
  NOR2_X1 U472 ( .A1(n26), .A2(n41), .ZN(ab_19__12_) );
  NOR2_X1 U473 ( .A1(n27), .A2(n41), .ZN(ab_19__11_) );
  NOR2_X1 U474 ( .A1(n28), .A2(n41), .ZN(ab_19__10_) );
  NOR2_X1 U475 ( .A1(n29), .A2(n41), .ZN(ab_19__0_) );
  NOR2_X1 U476 ( .A1(n7), .A2(n42), .ZN(ab_18__9_) );
  NOR2_X1 U477 ( .A1(n8), .A2(n42), .ZN(ab_18__8_) );
  NOR2_X1 U478 ( .A1(n9), .A2(n42), .ZN(ab_18__7_) );
  NOR2_X1 U479 ( .A1(n10), .A2(n42), .ZN(ab_18__6_) );
  NOR2_X1 U480 ( .A1(n11), .A2(n42), .ZN(ab_18__5_) );
  NOR2_X1 U481 ( .A1(n12), .A2(n42), .ZN(ab_18__4_) );
  NOR2_X1 U482 ( .A1(n13), .A2(n42), .ZN(ab_18__3_) );
  NOR2_X1 U483 ( .A1(n14), .A2(n42), .ZN(ab_18__2_) );
  NOR2_X1 U484 ( .A1(A[18]), .A2(n1), .ZN(ab_18__23_) );
  NOR2_X1 U485 ( .A1(n15), .A2(n42), .ZN(ab_18__22_) );
  NOR2_X1 U486 ( .A1(n16), .A2(n42), .ZN(ab_18__21_) );
  NOR2_X1 U487 ( .A1(n17), .A2(n42), .ZN(ab_18__20_) );
  NOR2_X1 U488 ( .A1(n18), .A2(n42), .ZN(ab_18__1_) );
  NOR2_X1 U489 ( .A1(n19), .A2(n42), .ZN(ab_18__19_) );
  NOR2_X1 U490 ( .A1(n20), .A2(n42), .ZN(ab_18__18_) );
  NOR2_X1 U491 ( .A1(n21), .A2(n42), .ZN(ab_18__17_) );
  NOR2_X1 U492 ( .A1(n22), .A2(n42), .ZN(ab_18__16_) );
  NOR2_X1 U493 ( .A1(n23), .A2(n42), .ZN(ab_18__15_) );
  NOR2_X1 U494 ( .A1(n24), .A2(n42), .ZN(ab_18__14_) );
  NOR2_X1 U495 ( .A1(n25), .A2(n42), .ZN(ab_18__13_) );
  NOR2_X1 U496 ( .A1(n26), .A2(n42), .ZN(ab_18__12_) );
  NOR2_X1 U497 ( .A1(n27), .A2(n42), .ZN(ab_18__11_) );
  NOR2_X1 U498 ( .A1(n28), .A2(n42), .ZN(ab_18__10_) );
  NOR2_X1 U499 ( .A1(n29), .A2(n42), .ZN(ab_18__0_) );
  NOR2_X1 U500 ( .A1(n7), .A2(n43), .ZN(ab_17__9_) );
  NOR2_X1 U501 ( .A1(n8), .A2(n43), .ZN(ab_17__8_) );
  NOR2_X1 U502 ( .A1(n9), .A2(n43), .ZN(ab_17__7_) );
  NOR2_X1 U503 ( .A1(n10), .A2(n43), .ZN(ab_17__6_) );
  NOR2_X1 U504 ( .A1(n11), .A2(n43), .ZN(ab_17__5_) );
  NOR2_X1 U505 ( .A1(n12), .A2(n43), .ZN(ab_17__4_) );
  NOR2_X1 U506 ( .A1(n13), .A2(n43), .ZN(ab_17__3_) );
  NOR2_X1 U507 ( .A1(n14), .A2(n43), .ZN(ab_17__2_) );
  NOR2_X1 U508 ( .A1(A[17]), .A2(n1), .ZN(ab_17__23_) );
  NOR2_X1 U509 ( .A1(n15), .A2(n43), .ZN(ab_17__22_) );
  NOR2_X1 U510 ( .A1(n16), .A2(n43), .ZN(ab_17__21_) );
  NOR2_X1 U511 ( .A1(n17), .A2(n43), .ZN(ab_17__20_) );
  NOR2_X1 U512 ( .A1(n18), .A2(n43), .ZN(ab_17__1_) );
  NOR2_X1 U513 ( .A1(n19), .A2(n43), .ZN(ab_17__19_) );
  NOR2_X1 U514 ( .A1(n20), .A2(n43), .ZN(ab_17__18_) );
  NOR2_X1 U515 ( .A1(n21), .A2(n43), .ZN(ab_17__17_) );
  NOR2_X1 U516 ( .A1(n22), .A2(n43), .ZN(ab_17__16_) );
  NOR2_X1 U517 ( .A1(n23), .A2(n43), .ZN(ab_17__15_) );
  NOR2_X1 U518 ( .A1(n24), .A2(n43), .ZN(ab_17__14_) );
  NOR2_X1 U519 ( .A1(n25), .A2(n43), .ZN(ab_17__13_) );
  NOR2_X1 U520 ( .A1(n26), .A2(n43), .ZN(ab_17__12_) );
  NOR2_X1 U521 ( .A1(n27), .A2(n43), .ZN(ab_17__11_) );
  NOR2_X1 U522 ( .A1(n28), .A2(n43), .ZN(ab_17__10_) );
  NOR2_X1 U523 ( .A1(n29), .A2(n43), .ZN(ab_17__0_) );
  NOR2_X1 U524 ( .A1(n7), .A2(n44), .ZN(ab_16__9_) );
  NOR2_X1 U525 ( .A1(n8), .A2(n44), .ZN(ab_16__8_) );
  NOR2_X1 U526 ( .A1(n9), .A2(n44), .ZN(ab_16__7_) );
  NOR2_X1 U527 ( .A1(n10), .A2(n44), .ZN(ab_16__6_) );
  NOR2_X1 U528 ( .A1(n11), .A2(n44), .ZN(ab_16__5_) );
  NOR2_X1 U529 ( .A1(n12), .A2(n44), .ZN(ab_16__4_) );
  NOR2_X1 U530 ( .A1(n13), .A2(n44), .ZN(ab_16__3_) );
  NOR2_X1 U531 ( .A1(n14), .A2(n44), .ZN(ab_16__2_) );
  NOR2_X1 U532 ( .A1(A[16]), .A2(n1), .ZN(ab_16__23_) );
  NOR2_X1 U533 ( .A1(n15), .A2(n44), .ZN(ab_16__22_) );
  NOR2_X1 U534 ( .A1(n16), .A2(n44), .ZN(ab_16__21_) );
  NOR2_X1 U535 ( .A1(n17), .A2(n44), .ZN(ab_16__20_) );
  NOR2_X1 U536 ( .A1(n18), .A2(n44), .ZN(ab_16__1_) );
  NOR2_X1 U537 ( .A1(n19), .A2(n44), .ZN(ab_16__19_) );
  NOR2_X1 U538 ( .A1(n20), .A2(n44), .ZN(ab_16__18_) );
  NOR2_X1 U539 ( .A1(n21), .A2(n44), .ZN(ab_16__17_) );
  NOR2_X1 U540 ( .A1(n22), .A2(n44), .ZN(ab_16__16_) );
  NOR2_X1 U541 ( .A1(n23), .A2(n44), .ZN(ab_16__15_) );
  NOR2_X1 U542 ( .A1(n24), .A2(n44), .ZN(ab_16__14_) );
  NOR2_X1 U543 ( .A1(n25), .A2(n44), .ZN(ab_16__13_) );
  NOR2_X1 U544 ( .A1(n26), .A2(n44), .ZN(ab_16__12_) );
  NOR2_X1 U545 ( .A1(n27), .A2(n44), .ZN(ab_16__11_) );
  NOR2_X1 U546 ( .A1(n28), .A2(n44), .ZN(ab_16__10_) );
  NOR2_X1 U547 ( .A1(n29), .A2(n44), .ZN(ab_16__0_) );
  NOR2_X1 U548 ( .A1(n7), .A2(n45), .ZN(ab_15__9_) );
  NOR2_X1 U549 ( .A1(n8), .A2(n45), .ZN(ab_15__8_) );
  NOR2_X1 U550 ( .A1(n9), .A2(n45), .ZN(ab_15__7_) );
  NOR2_X1 U551 ( .A1(n10), .A2(n45), .ZN(ab_15__6_) );
  NOR2_X1 U552 ( .A1(n11), .A2(n45), .ZN(ab_15__5_) );
  NOR2_X1 U553 ( .A1(n12), .A2(n45), .ZN(ab_15__4_) );
  NOR2_X1 U554 ( .A1(n13), .A2(n45), .ZN(ab_15__3_) );
  NOR2_X1 U555 ( .A1(n14), .A2(n45), .ZN(ab_15__2_) );
  NOR2_X1 U556 ( .A1(A[15]), .A2(n1), .ZN(ab_15__23_) );
  NOR2_X1 U557 ( .A1(n15), .A2(n45), .ZN(ab_15__22_) );
  NOR2_X1 U558 ( .A1(n16), .A2(n45), .ZN(ab_15__21_) );
  NOR2_X1 U559 ( .A1(n17), .A2(n45), .ZN(ab_15__20_) );
  NOR2_X1 U560 ( .A1(n18), .A2(n45), .ZN(ab_15__1_) );
  NOR2_X1 U561 ( .A1(n19), .A2(n45), .ZN(ab_15__19_) );
  NOR2_X1 U562 ( .A1(n20), .A2(n45), .ZN(ab_15__18_) );
  NOR2_X1 U563 ( .A1(n21), .A2(n45), .ZN(ab_15__17_) );
  NOR2_X1 U564 ( .A1(n22), .A2(n45), .ZN(ab_15__16_) );
  NOR2_X1 U565 ( .A1(n23), .A2(n45), .ZN(ab_15__15_) );
  NOR2_X1 U566 ( .A1(n24), .A2(n45), .ZN(ab_15__14_) );
  NOR2_X1 U567 ( .A1(n25), .A2(n45), .ZN(ab_15__13_) );
  NOR2_X1 U568 ( .A1(n26), .A2(n45), .ZN(ab_15__12_) );
  NOR2_X1 U569 ( .A1(n27), .A2(n45), .ZN(ab_15__11_) );
  NOR2_X1 U570 ( .A1(n28), .A2(n45), .ZN(ab_15__10_) );
  NOR2_X1 U571 ( .A1(n29), .A2(n45), .ZN(ab_15__0_) );
  NOR2_X1 U572 ( .A1(n7), .A2(n46), .ZN(ab_14__9_) );
  NOR2_X1 U573 ( .A1(n8), .A2(n46), .ZN(ab_14__8_) );
  NOR2_X1 U574 ( .A1(n9), .A2(n46), .ZN(ab_14__7_) );
  NOR2_X1 U575 ( .A1(n10), .A2(n46), .ZN(ab_14__6_) );
  NOR2_X1 U576 ( .A1(n11), .A2(n46), .ZN(ab_14__5_) );
  NOR2_X1 U577 ( .A1(n12), .A2(n46), .ZN(ab_14__4_) );
  NOR2_X1 U578 ( .A1(n13), .A2(n46), .ZN(ab_14__3_) );
  NOR2_X1 U579 ( .A1(n14), .A2(n46), .ZN(ab_14__2_) );
  NOR2_X1 U580 ( .A1(A[14]), .A2(n2), .ZN(ab_14__23_) );
  NOR2_X1 U581 ( .A1(n15), .A2(n46), .ZN(ab_14__22_) );
  NOR2_X1 U582 ( .A1(n16), .A2(n46), .ZN(ab_14__21_) );
  NOR2_X1 U583 ( .A1(n17), .A2(n46), .ZN(ab_14__20_) );
  NOR2_X1 U584 ( .A1(n18), .A2(n46), .ZN(ab_14__1_) );
  NOR2_X1 U585 ( .A1(n19), .A2(n46), .ZN(ab_14__19_) );
  NOR2_X1 U586 ( .A1(n20), .A2(n46), .ZN(ab_14__18_) );
  NOR2_X1 U587 ( .A1(n21), .A2(n46), .ZN(ab_14__17_) );
  NOR2_X1 U588 ( .A1(n22), .A2(n46), .ZN(ab_14__16_) );
  NOR2_X1 U589 ( .A1(n23), .A2(n46), .ZN(ab_14__15_) );
  NOR2_X1 U590 ( .A1(n24), .A2(n46), .ZN(ab_14__14_) );
  NOR2_X1 U591 ( .A1(n25), .A2(n46), .ZN(ab_14__13_) );
  NOR2_X1 U592 ( .A1(n26), .A2(n46), .ZN(ab_14__12_) );
  NOR2_X1 U593 ( .A1(n27), .A2(n46), .ZN(ab_14__11_) );
  NOR2_X1 U594 ( .A1(n28), .A2(n46), .ZN(ab_14__10_) );
  NOR2_X1 U595 ( .A1(n29), .A2(n46), .ZN(ab_14__0_) );
  NOR2_X1 U596 ( .A1(n7), .A2(n47), .ZN(ab_13__9_) );
  NOR2_X1 U597 ( .A1(n8), .A2(n47), .ZN(ab_13__8_) );
  NOR2_X1 U598 ( .A1(n9), .A2(n47), .ZN(ab_13__7_) );
  NOR2_X1 U599 ( .A1(n10), .A2(n47), .ZN(ab_13__6_) );
  NOR2_X1 U600 ( .A1(n11), .A2(n47), .ZN(ab_13__5_) );
  NOR2_X1 U601 ( .A1(n12), .A2(n47), .ZN(ab_13__4_) );
  NOR2_X1 U602 ( .A1(n13), .A2(n47), .ZN(ab_13__3_) );
  NOR2_X1 U603 ( .A1(n14), .A2(n47), .ZN(ab_13__2_) );
  NOR2_X1 U604 ( .A1(A[13]), .A2(n2), .ZN(ab_13__23_) );
  NOR2_X1 U605 ( .A1(n15), .A2(n47), .ZN(ab_13__22_) );
  NOR2_X1 U606 ( .A1(n16), .A2(n47), .ZN(ab_13__21_) );
  NOR2_X1 U607 ( .A1(n17), .A2(n47), .ZN(ab_13__20_) );
  NOR2_X1 U608 ( .A1(n18), .A2(n47), .ZN(ab_13__1_) );
  NOR2_X1 U609 ( .A1(n19), .A2(n47), .ZN(ab_13__19_) );
  NOR2_X1 U610 ( .A1(n20), .A2(n47), .ZN(ab_13__18_) );
  NOR2_X1 U611 ( .A1(n21), .A2(n47), .ZN(ab_13__17_) );
  NOR2_X1 U612 ( .A1(n22), .A2(n47), .ZN(ab_13__16_) );
  NOR2_X1 U613 ( .A1(n23), .A2(n47), .ZN(ab_13__15_) );
  NOR2_X1 U614 ( .A1(n24), .A2(n47), .ZN(ab_13__14_) );
  NOR2_X1 U615 ( .A1(n25), .A2(n47), .ZN(ab_13__13_) );
  NOR2_X1 U616 ( .A1(n26), .A2(n47), .ZN(ab_13__12_) );
  NOR2_X1 U617 ( .A1(n27), .A2(n47), .ZN(ab_13__11_) );
  NOR2_X1 U618 ( .A1(n28), .A2(n47), .ZN(ab_13__10_) );
  NOR2_X1 U619 ( .A1(n29), .A2(n47), .ZN(ab_13__0_) );
  NOR2_X1 U620 ( .A1(n7), .A2(n48), .ZN(ab_12__9_) );
  NOR2_X1 U621 ( .A1(n8), .A2(n48), .ZN(ab_12__8_) );
  NOR2_X1 U622 ( .A1(n9), .A2(n48), .ZN(ab_12__7_) );
  NOR2_X1 U623 ( .A1(n10), .A2(n48), .ZN(ab_12__6_) );
  NOR2_X1 U624 ( .A1(n11), .A2(n48), .ZN(ab_12__5_) );
  NOR2_X1 U625 ( .A1(n12), .A2(n48), .ZN(ab_12__4_) );
  NOR2_X1 U626 ( .A1(n13), .A2(n48), .ZN(ab_12__3_) );
  NOR2_X1 U627 ( .A1(n14), .A2(n48), .ZN(ab_12__2_) );
  NOR2_X1 U628 ( .A1(A[12]), .A2(n2), .ZN(ab_12__23_) );
  NOR2_X1 U629 ( .A1(n15), .A2(n48), .ZN(ab_12__22_) );
  NOR2_X1 U630 ( .A1(n16), .A2(n48), .ZN(ab_12__21_) );
  NOR2_X1 U631 ( .A1(n17), .A2(n48), .ZN(ab_12__20_) );
  NOR2_X1 U632 ( .A1(n18), .A2(n48), .ZN(ab_12__1_) );
  NOR2_X1 U633 ( .A1(n19), .A2(n48), .ZN(ab_12__19_) );
  NOR2_X1 U634 ( .A1(n20), .A2(n48), .ZN(ab_12__18_) );
  NOR2_X1 U635 ( .A1(n21), .A2(n48), .ZN(ab_12__17_) );
  NOR2_X1 U636 ( .A1(n22), .A2(n48), .ZN(ab_12__16_) );
  NOR2_X1 U637 ( .A1(n23), .A2(n48), .ZN(ab_12__15_) );
  NOR2_X1 U638 ( .A1(n24), .A2(n48), .ZN(ab_12__14_) );
  NOR2_X1 U639 ( .A1(n25), .A2(n48), .ZN(ab_12__13_) );
  NOR2_X1 U640 ( .A1(n26), .A2(n48), .ZN(ab_12__12_) );
  NOR2_X1 U641 ( .A1(n27), .A2(n48), .ZN(ab_12__11_) );
  NOR2_X1 U642 ( .A1(n28), .A2(n48), .ZN(ab_12__10_) );
  NOR2_X1 U643 ( .A1(n29), .A2(n48), .ZN(ab_12__0_) );
  NOR2_X1 U644 ( .A1(n7), .A2(n49), .ZN(ab_11__9_) );
  NOR2_X1 U645 ( .A1(n8), .A2(n49), .ZN(ab_11__8_) );
  NOR2_X1 U646 ( .A1(n9), .A2(n49), .ZN(ab_11__7_) );
  NOR2_X1 U647 ( .A1(n10), .A2(n49), .ZN(ab_11__6_) );
  NOR2_X1 U648 ( .A1(n11), .A2(n49), .ZN(ab_11__5_) );
  NOR2_X1 U649 ( .A1(n12), .A2(n49), .ZN(ab_11__4_) );
  NOR2_X1 U650 ( .A1(n13), .A2(n49), .ZN(ab_11__3_) );
  NOR2_X1 U651 ( .A1(n14), .A2(n49), .ZN(ab_11__2_) );
  NOR2_X1 U652 ( .A1(A[11]), .A2(n2), .ZN(ab_11__23_) );
  NOR2_X1 U653 ( .A1(n15), .A2(n49), .ZN(ab_11__22_) );
  NOR2_X1 U654 ( .A1(n16), .A2(n49), .ZN(ab_11__21_) );
  NOR2_X1 U655 ( .A1(n17), .A2(n49), .ZN(ab_11__20_) );
  NOR2_X1 U656 ( .A1(n18), .A2(n49), .ZN(ab_11__1_) );
  NOR2_X1 U657 ( .A1(n19), .A2(n49), .ZN(ab_11__19_) );
  NOR2_X1 U658 ( .A1(n20), .A2(n49), .ZN(ab_11__18_) );
  NOR2_X1 U659 ( .A1(n21), .A2(n49), .ZN(ab_11__17_) );
  NOR2_X1 U660 ( .A1(n22), .A2(n49), .ZN(ab_11__16_) );
  NOR2_X1 U661 ( .A1(n23), .A2(n49), .ZN(ab_11__15_) );
  NOR2_X1 U662 ( .A1(n24), .A2(n49), .ZN(ab_11__14_) );
  NOR2_X1 U663 ( .A1(n25), .A2(n49), .ZN(ab_11__13_) );
  NOR2_X1 U664 ( .A1(n26), .A2(n49), .ZN(ab_11__12_) );
  NOR2_X1 U665 ( .A1(n27), .A2(n49), .ZN(ab_11__11_) );
  NOR2_X1 U666 ( .A1(n28), .A2(n49), .ZN(ab_11__10_) );
  NOR2_X1 U667 ( .A1(n29), .A2(n49), .ZN(ab_11__0_) );
  NOR2_X1 U668 ( .A1(n7), .A2(n50), .ZN(ab_10__9_) );
  NOR2_X1 U669 ( .A1(n8), .A2(n50), .ZN(ab_10__8_) );
  NOR2_X1 U670 ( .A1(n9), .A2(n50), .ZN(ab_10__7_) );
  NOR2_X1 U671 ( .A1(n10), .A2(n50), .ZN(ab_10__6_) );
  NOR2_X1 U672 ( .A1(n11), .A2(n50), .ZN(ab_10__5_) );
  NOR2_X1 U673 ( .A1(n12), .A2(n50), .ZN(ab_10__4_) );
  NOR2_X1 U674 ( .A1(n13), .A2(n50), .ZN(ab_10__3_) );
  NOR2_X1 U675 ( .A1(n14), .A2(n50), .ZN(ab_10__2_) );
  NOR2_X1 U676 ( .A1(A[10]), .A2(n2), .ZN(ab_10__23_) );
  NOR2_X1 U677 ( .A1(n15), .A2(n50), .ZN(ab_10__22_) );
  NOR2_X1 U678 ( .A1(n16), .A2(n50), .ZN(ab_10__21_) );
  NOR2_X1 U679 ( .A1(n17), .A2(n50), .ZN(ab_10__20_) );
  NOR2_X1 U680 ( .A1(n18), .A2(n50), .ZN(ab_10__1_) );
  NOR2_X1 U681 ( .A1(n19), .A2(n50), .ZN(ab_10__19_) );
  NOR2_X1 U682 ( .A1(n20), .A2(n50), .ZN(ab_10__18_) );
  NOR2_X1 U683 ( .A1(n21), .A2(n50), .ZN(ab_10__17_) );
  NOR2_X1 U684 ( .A1(n22), .A2(n50), .ZN(ab_10__16_) );
  NOR2_X1 U685 ( .A1(n23), .A2(n50), .ZN(ab_10__15_) );
  NOR2_X1 U686 ( .A1(n24), .A2(n50), .ZN(ab_10__14_) );
  NOR2_X1 U687 ( .A1(n25), .A2(n50), .ZN(ab_10__13_) );
  NOR2_X1 U688 ( .A1(n26), .A2(n50), .ZN(ab_10__12_) );
  NOR2_X1 U689 ( .A1(n27), .A2(n50), .ZN(ab_10__11_) );
  NOR2_X1 U690 ( .A1(n28), .A2(n50), .ZN(ab_10__10_) );
  NOR2_X1 U691 ( .A1(n29), .A2(n50), .ZN(ab_10__0_) );
  NOR2_X1 U692 ( .A1(n7), .A2(n51), .ZN(ab_0__9_) );
  NOR2_X1 U693 ( .A1(n8), .A2(n51), .ZN(ab_0__8_) );
  NOR2_X1 U694 ( .A1(n9), .A2(n51), .ZN(ab_0__7_) );
  NOR2_X1 U695 ( .A1(n10), .A2(n51), .ZN(ab_0__6_) );
  NOR2_X1 U696 ( .A1(n11), .A2(n51), .ZN(ab_0__5_) );
  NOR2_X1 U697 ( .A1(n12), .A2(n51), .ZN(ab_0__4_) );
  NOR2_X1 U698 ( .A1(n13), .A2(n51), .ZN(ab_0__3_) );
  NOR2_X1 U699 ( .A1(n14), .A2(n51), .ZN(ab_0__2_) );
  NOR2_X1 U700 ( .A1(A[0]), .A2(n1), .ZN(ab_0__23_) );
  NOR2_X1 U701 ( .A1(n15), .A2(n51), .ZN(ab_0__22_) );
  NOR2_X1 U702 ( .A1(n16), .A2(n51), .ZN(ab_0__21_) );
  NOR2_X1 U703 ( .A1(n17), .A2(n51), .ZN(ab_0__20_) );
  NOR2_X1 U704 ( .A1(n19), .A2(n51), .ZN(ab_0__19_) );
  NOR2_X1 U705 ( .A1(n20), .A2(n51), .ZN(ab_0__18_) );
  NOR2_X1 U706 ( .A1(n21), .A2(n51), .ZN(ab_0__17_) );
  NOR2_X1 U707 ( .A1(n22), .A2(n51), .ZN(ab_0__16_) );
  NOR2_X1 U708 ( .A1(n23), .A2(n51), .ZN(ab_0__15_) );
  NOR2_X1 U709 ( .A1(n24), .A2(n51), .ZN(ab_0__14_) );
  NOR2_X1 U710 ( .A1(n25), .A2(n51), .ZN(ab_0__13_) );
  NOR2_X1 U711 ( .A1(n26), .A2(n51), .ZN(ab_0__12_) );
  NOR2_X1 U712 ( .A1(n27), .A2(n51), .ZN(ab_0__11_) );
  NOR2_X1 U713 ( .A1(n28), .A2(n51), .ZN(ab_0__10_) );
  INV_X1 U714 ( .A(B[23]), .ZN(QB) );
  INV_X1 U715 ( .A(A[23]), .ZN(QA) );
  AND3_X1 U716 ( .A1(ab_1__1_), .A2(B[0]), .A3(A[0]), .ZN(CARRYB_1__0_) );
  NOR2_X1 U717 ( .A1(n40), .A2(n18), .ZN(ab_1__1_) );
  INV_X1 U719 ( .A(CARRYB_23__23_), .ZN(A1_45_) );
endmodule


module iir_filter_DW01_add_7 ( A, B, CI, SUM, CO );
  input [45:0] A;
  input [45:0] B;
  output [45:0] SUM;
  input CI;
  output CO;
  wire   A_21_, A_20_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112;
  assign SUM[21] = A_21_;
  assign A_21_ = A[21];
  assign SUM[20] = A_20_;
  assign A_20_ = A[20];

  XOR2_X1 U2 ( .A(n1), .B(n2), .Z(SUM[45]) );
  XOR2_X1 U3 ( .A(B[45]), .B(A[45]), .Z(n2) );
  OAI21_X1 U4 ( .B1(n3), .B2(n4), .A(n5), .ZN(n1) );
  OAI21_X1 U5 ( .B1(A[44]), .B2(n6), .A(B[44]), .ZN(n5) );
  INV_X1 U6 ( .A(n3), .ZN(n6) );
  INV_X1 U7 ( .A(A[44]), .ZN(n4) );
  AOI21_X1 U8 ( .B1(A[43]), .B2(B[43]), .A(n7), .ZN(n3) );
  INV_X1 U9 ( .A(n8), .ZN(n7) );
  OAI22_X1 U10 ( .A1(n9), .A2(n10), .B1(A[43]), .B2(B[43]), .ZN(n8) );
  AOI21_X1 U11 ( .B1(n11), .B2(n12), .A(n13), .ZN(n9) );
  NAND3_X1 U12 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n12) );
  AOI21_X1 U13 ( .B1(n17), .B2(n16), .A(n18), .ZN(n11) );
  INV_X1 U14 ( .A(n19), .ZN(n18) );
  XOR2_X1 U15 ( .A(n20), .B(n21), .Z(SUM[42]) );
  NOR2_X1 U16 ( .A1(n10), .A2(n13), .ZN(n21) );
  NOR2_X1 U17 ( .A1(B[42]), .A2(A[42]), .ZN(n13) );
  AND2_X1 U18 ( .A1(B[42]), .A2(A[42]), .ZN(n10) );
  OAI21_X1 U19 ( .B1(n22), .B2(n23), .A(n19), .ZN(n20) );
  XOR2_X1 U20 ( .A(n24), .B(n23), .Z(SUM[41]) );
  AOI21_X1 U21 ( .B1(n15), .B2(n14), .A(n17), .ZN(n23) );
  INV_X1 U22 ( .A(n25), .ZN(n15) );
  NAND2_X1 U23 ( .A1(n16), .A2(n19), .ZN(n24) );
  NAND2_X1 U24 ( .A1(B[41]), .A2(A[41]), .ZN(n19) );
  INV_X1 U25 ( .A(n22), .ZN(n16) );
  NOR2_X1 U26 ( .A1(B[41]), .A2(A[41]), .ZN(n22) );
  XOR2_X1 U27 ( .A(n14), .B(n26), .Z(SUM[40]) );
  NOR2_X1 U28 ( .A1(n17), .A2(n25), .ZN(n26) );
  NOR2_X1 U29 ( .A1(B[40]), .A2(A[40]), .ZN(n25) );
  AND2_X1 U30 ( .A1(B[40]), .A2(A[40]), .ZN(n17) );
  OAI21_X1 U31 ( .B1(n27), .B2(n28), .A(n29), .ZN(n14) );
  XOR2_X1 U32 ( .A(n30), .B(n28), .Z(SUM[39]) );
  AOI21_X1 U33 ( .B1(n31), .B2(n32), .A(n33), .ZN(n28) );
  INV_X1 U34 ( .A(n34), .ZN(n31) );
  NAND2_X1 U35 ( .A1(n35), .A2(n29), .ZN(n30) );
  NAND2_X1 U36 ( .A1(B[39]), .A2(A[39]), .ZN(n29) );
  INV_X1 U37 ( .A(n27), .ZN(n35) );
  NOR2_X1 U38 ( .A1(B[39]), .A2(A[39]), .ZN(n27) );
  XOR2_X1 U39 ( .A(n32), .B(n36), .Z(SUM[38]) );
  NOR2_X1 U40 ( .A1(n33), .A2(n34), .ZN(n36) );
  NOR2_X1 U41 ( .A1(B[38]), .A2(A[38]), .ZN(n34) );
  AND2_X1 U42 ( .A1(B[38]), .A2(A[38]), .ZN(n33) );
  OAI21_X1 U43 ( .B1(n37), .B2(n38), .A(n39), .ZN(n32) );
  XOR2_X1 U44 ( .A(n40), .B(n38), .Z(SUM[37]) );
  AOI21_X1 U45 ( .B1(n41), .B2(n42), .A(n43), .ZN(n38) );
  INV_X1 U46 ( .A(n44), .ZN(n41) );
  NAND2_X1 U47 ( .A1(n45), .A2(n39), .ZN(n40) );
  NAND2_X1 U48 ( .A1(B[37]), .A2(A[37]), .ZN(n39) );
  INV_X1 U49 ( .A(n37), .ZN(n45) );
  NOR2_X1 U50 ( .A1(B[37]), .A2(A[37]), .ZN(n37) );
  XOR2_X1 U51 ( .A(n42), .B(n46), .Z(SUM[36]) );
  NOR2_X1 U52 ( .A1(n43), .A2(n44), .ZN(n46) );
  NOR2_X1 U53 ( .A1(B[36]), .A2(A[36]), .ZN(n44) );
  AND2_X1 U54 ( .A1(B[36]), .A2(A[36]), .ZN(n43) );
  OAI21_X1 U55 ( .B1(n47), .B2(n48), .A(n49), .ZN(n42) );
  XOR2_X1 U56 ( .A(n50), .B(n48), .Z(SUM[35]) );
  AOI21_X1 U57 ( .B1(n51), .B2(n52), .A(n53), .ZN(n48) );
  INV_X1 U58 ( .A(n54), .ZN(n51) );
  NAND2_X1 U59 ( .A1(n55), .A2(n49), .ZN(n50) );
  NAND2_X1 U60 ( .A1(B[35]), .A2(A[35]), .ZN(n49) );
  INV_X1 U61 ( .A(n47), .ZN(n55) );
  NOR2_X1 U62 ( .A1(B[35]), .A2(A[35]), .ZN(n47) );
  XOR2_X1 U63 ( .A(n52), .B(n56), .Z(SUM[34]) );
  NOR2_X1 U64 ( .A1(n53), .A2(n54), .ZN(n56) );
  NOR2_X1 U65 ( .A1(B[34]), .A2(A[34]), .ZN(n54) );
  AND2_X1 U66 ( .A1(B[34]), .A2(A[34]), .ZN(n53) );
  OAI21_X1 U67 ( .B1(n57), .B2(n58), .A(n59), .ZN(n52) );
  XOR2_X1 U68 ( .A(n60), .B(n58), .Z(SUM[33]) );
  AOI21_X1 U69 ( .B1(n61), .B2(n62), .A(n63), .ZN(n58) );
  INV_X1 U70 ( .A(n64), .ZN(n61) );
  NAND2_X1 U71 ( .A1(n65), .A2(n59), .ZN(n60) );
  NAND2_X1 U72 ( .A1(B[33]), .A2(A[33]), .ZN(n59) );
  INV_X1 U73 ( .A(n57), .ZN(n65) );
  NOR2_X1 U74 ( .A1(B[33]), .A2(A[33]), .ZN(n57) );
  XOR2_X1 U75 ( .A(n62), .B(n66), .Z(SUM[32]) );
  NOR2_X1 U76 ( .A1(n63), .A2(n64), .ZN(n66) );
  NOR2_X1 U77 ( .A1(B[32]), .A2(A[32]), .ZN(n64) );
  AND2_X1 U78 ( .A1(B[32]), .A2(A[32]), .ZN(n63) );
  OAI21_X1 U79 ( .B1(n67), .B2(n68), .A(n69), .ZN(n62) );
  XOR2_X1 U80 ( .A(n70), .B(n68), .Z(SUM[31]) );
  AOI21_X1 U81 ( .B1(n71), .B2(n72), .A(n73), .ZN(n68) );
  INV_X1 U82 ( .A(n74), .ZN(n71) );
  NAND2_X1 U83 ( .A1(n75), .A2(n69), .ZN(n70) );
  NAND2_X1 U84 ( .A1(B[31]), .A2(A[31]), .ZN(n69) );
  INV_X1 U85 ( .A(n67), .ZN(n75) );
  NOR2_X1 U86 ( .A1(B[31]), .A2(A[31]), .ZN(n67) );
  XOR2_X1 U87 ( .A(n72), .B(n76), .Z(SUM[30]) );
  NOR2_X1 U88 ( .A1(n73), .A2(n74), .ZN(n76) );
  NOR2_X1 U89 ( .A1(B[30]), .A2(A[30]), .ZN(n74) );
  AND2_X1 U90 ( .A1(B[30]), .A2(A[30]), .ZN(n73) );
  OAI21_X1 U91 ( .B1(n77), .B2(n78), .A(n79), .ZN(n72) );
  XOR2_X1 U92 ( .A(n80), .B(n78), .Z(SUM[29]) );
  AOI21_X1 U93 ( .B1(n81), .B2(n82), .A(n83), .ZN(n78) );
  INV_X1 U94 ( .A(n84), .ZN(n81) );
  NAND2_X1 U95 ( .A1(n85), .A2(n79), .ZN(n80) );
  NAND2_X1 U96 ( .A1(B[29]), .A2(A[29]), .ZN(n79) );
  INV_X1 U97 ( .A(n77), .ZN(n85) );
  NOR2_X1 U98 ( .A1(B[29]), .A2(A[29]), .ZN(n77) );
  XOR2_X1 U99 ( .A(n82), .B(n86), .Z(SUM[28]) );
  NOR2_X1 U100 ( .A1(n83), .A2(n84), .ZN(n86) );
  NOR2_X1 U101 ( .A1(B[28]), .A2(A[28]), .ZN(n84) );
  AND2_X1 U102 ( .A1(B[28]), .A2(A[28]), .ZN(n83) );
  OAI21_X1 U103 ( .B1(n87), .B2(n88), .A(n89), .ZN(n82) );
  XOR2_X1 U104 ( .A(n90), .B(n88), .Z(SUM[27]) );
  AOI21_X1 U105 ( .B1(n91), .B2(n92), .A(n93), .ZN(n88) );
  INV_X1 U106 ( .A(n94), .ZN(n92) );
  NAND2_X1 U107 ( .A1(n95), .A2(n89), .ZN(n90) );
  NAND2_X1 U108 ( .A1(B[27]), .A2(A[27]), .ZN(n89) );
  INV_X1 U109 ( .A(n87), .ZN(n95) );
  NOR2_X1 U110 ( .A1(B[27]), .A2(A[27]), .ZN(n87) );
  XOR2_X1 U111 ( .A(n91), .B(n96), .Z(SUM[26]) );
  NOR2_X1 U112 ( .A1(n93), .A2(n94), .ZN(n96) );
  NOR2_X1 U113 ( .A1(B[26]), .A2(A[26]), .ZN(n94) );
  AND2_X1 U114 ( .A1(B[26]), .A2(A[26]), .ZN(n93) );
  OAI21_X1 U115 ( .B1(n97), .B2(n98), .A(n99), .ZN(n91) );
  XOR2_X1 U116 ( .A(n100), .B(n98), .Z(SUM[25]) );
  AOI21_X1 U117 ( .B1(n101), .B2(n102), .A(n103), .ZN(n98) );
  INV_X1 U118 ( .A(n104), .ZN(n101) );
  NAND2_X1 U119 ( .A1(n105), .A2(n99), .ZN(n100) );
  NAND2_X1 U120 ( .A1(B[25]), .A2(A[25]), .ZN(n99) );
  INV_X1 U121 ( .A(n97), .ZN(n105) );
  NOR2_X1 U122 ( .A1(B[25]), .A2(A[25]), .ZN(n97) );
  XOR2_X1 U123 ( .A(n102), .B(n106), .Z(SUM[24]) );
  NOR2_X1 U124 ( .A1(n103), .A2(n104), .ZN(n106) );
  NOR2_X1 U125 ( .A1(B[24]), .A2(A[24]), .ZN(n104) );
  AND2_X1 U126 ( .A1(B[24]), .A2(A[24]), .ZN(n103) );
  OAI21_X1 U127 ( .B1(n107), .B2(n108), .A(n109), .ZN(n102) );
  XOR2_X1 U128 ( .A(n108), .B(n110), .Z(SUM[23]) );
  NAND2_X1 U129 ( .A1(n111), .A2(n109), .ZN(n110) );
  NAND2_X1 U130 ( .A1(B[23]), .A2(A[23]), .ZN(n109) );
  INV_X1 U131 ( .A(n107), .ZN(n111) );
  NOR2_X1 U132 ( .A1(B[23]), .A2(A[23]), .ZN(n107) );
  INV_X1 U133 ( .A(n112), .ZN(SUM[22]) );
  OAI21_X1 U134 ( .B1(B[22]), .B2(A[22]), .A(n108), .ZN(n112) );
  NAND2_X1 U135 ( .A1(B[22]), .A2(A[22]), .ZN(n108) );
endmodule


module iir_filter_DW02_mult_3 ( A, B, TC, PRODUCT );
  input [23:0] A;
  input [23:0] B;
  output [47:0] PRODUCT;
  input TC;
  wire   ab_23__23_, ab_23__22_, ab_23__21_, ab_23__20_, ab_23__19_,
         ab_23__18_, ab_23__17_, ab_23__16_, ab_23__15_, ab_23__14_,
         ab_23__13_, ab_23__12_, ab_23__11_, ab_23__10_, ab_23__9_, ab_23__8_,
         ab_23__7_, ab_23__6_, ab_23__5_, ab_23__4_, ab_23__3_, ab_23__2_,
         ab_23__1_, ab_23__0_, ab_22__23_, ab_22__22_, ab_22__21_, ab_22__20_,
         ab_22__19_, ab_22__18_, ab_22__17_, ab_22__16_, ab_22__15_,
         ab_22__14_, ab_22__13_, ab_22__12_, ab_22__11_, ab_22__10_, ab_22__9_,
         ab_22__8_, ab_22__7_, ab_22__6_, ab_22__5_, ab_22__4_, ab_22__3_,
         ab_22__2_, ab_22__1_, ab_22__0_, ab_21__23_, ab_21__22_, ab_21__21_,
         ab_21__20_, ab_21__19_, ab_21__18_, ab_21__17_, ab_21__16_,
         ab_21__15_, ab_21__14_, ab_21__13_, ab_21__12_, ab_21__11_,
         ab_21__10_, ab_21__9_, ab_21__8_, ab_21__7_, ab_21__6_, ab_21__5_,
         ab_21__4_, ab_21__3_, ab_21__2_, ab_21__1_, ab_21__0_, ab_20__23_,
         ab_20__22_, ab_20__21_, ab_20__20_, ab_20__19_, ab_20__18_,
         ab_20__17_, ab_20__16_, ab_20__15_, ab_20__14_, ab_20__13_,
         ab_20__12_, ab_20__11_, ab_20__10_, ab_20__9_, ab_20__8_, ab_20__7_,
         ab_20__6_, ab_20__5_, ab_20__4_, ab_20__3_, ab_20__2_, ab_20__1_,
         ab_20__0_, ab_19__23_, ab_19__22_, ab_19__21_, ab_19__20_, ab_19__19_,
         ab_19__18_, ab_19__17_, ab_19__16_, ab_19__15_, ab_19__14_,
         ab_19__13_, ab_19__12_, ab_19__11_, ab_19__10_, ab_19__9_, ab_19__8_,
         ab_19__7_, ab_19__6_, ab_19__5_, ab_19__4_, ab_19__3_, ab_19__2_,
         ab_19__1_, ab_19__0_, ab_18__23_, ab_18__22_, ab_18__21_, ab_18__20_,
         ab_18__19_, ab_18__18_, ab_18__17_, ab_18__16_, ab_18__15_,
         ab_18__14_, ab_18__13_, ab_18__12_, ab_18__11_, ab_18__10_, ab_18__9_,
         ab_18__8_, ab_18__7_, ab_18__6_, ab_18__5_, ab_18__4_, ab_18__3_,
         ab_18__2_, ab_18__1_, ab_18__0_, ab_17__23_, ab_17__22_, ab_17__21_,
         ab_17__20_, ab_17__19_, ab_17__18_, ab_17__17_, ab_17__16_,
         ab_17__15_, ab_17__14_, ab_17__13_, ab_17__12_, ab_17__11_,
         ab_17__10_, ab_17__9_, ab_17__8_, ab_17__7_, ab_17__6_, ab_17__5_,
         ab_17__4_, ab_17__3_, ab_17__2_, ab_17__1_, ab_17__0_, ab_16__23_,
         ab_16__22_, ab_16__21_, ab_16__20_, ab_16__19_, ab_16__18_,
         ab_16__17_, ab_16__16_, ab_16__15_, ab_16__14_, ab_16__13_,
         ab_16__12_, ab_16__11_, ab_16__10_, ab_16__9_, ab_16__8_, ab_16__7_,
         ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_, ab_16__1_,
         ab_16__0_, ab_15__23_, ab_15__22_, ab_15__21_, ab_15__20_, ab_15__19_,
         ab_15__18_, ab_15__17_, ab_15__16_, ab_15__15_, ab_15__14_,
         ab_15__13_, ab_15__12_, ab_15__11_, ab_15__10_, ab_15__9_, ab_15__8_,
         ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_, ab_15__3_, ab_15__2_,
         ab_15__1_, ab_15__0_, ab_14__23_, ab_14__22_, ab_14__21_, ab_14__20_,
         ab_14__19_, ab_14__18_, ab_14__17_, ab_14__16_, ab_14__15_,
         ab_14__14_, ab_14__13_, ab_14__12_, ab_14__11_, ab_14__10_, ab_14__9_,
         ab_14__8_, ab_14__7_, ab_14__6_, ab_14__5_, ab_14__4_, ab_14__3_,
         ab_14__2_, ab_14__1_, ab_14__0_, ab_13__23_, ab_13__22_, ab_13__21_,
         ab_13__20_, ab_13__19_, ab_13__18_, ab_13__17_, ab_13__16_,
         ab_13__15_, ab_13__14_, ab_13__13_, ab_13__12_, ab_13__11_,
         ab_13__10_, ab_13__9_, ab_13__8_, ab_13__7_, ab_13__6_, ab_13__5_,
         ab_13__4_, ab_13__3_, ab_13__2_, ab_13__1_, ab_13__0_, ab_12__23_,
         ab_12__22_, ab_12__21_, ab_12__20_, ab_12__19_, ab_12__18_,
         ab_12__17_, ab_12__16_, ab_12__15_, ab_12__14_, ab_12__13_,
         ab_12__12_, ab_12__11_, ab_12__10_, ab_12__9_, ab_12__8_, ab_12__7_,
         ab_12__6_, ab_12__5_, ab_12__4_, ab_12__3_, ab_12__2_, ab_12__1_,
         ab_12__0_, ab_11__23_, ab_11__22_, ab_11__21_, ab_11__20_, ab_11__19_,
         ab_11__18_, ab_11__17_, ab_11__16_, ab_11__15_, ab_11__14_,
         ab_11__13_, ab_11__12_, ab_11__11_, ab_11__10_, ab_11__9_, ab_11__8_,
         ab_11__7_, ab_11__6_, ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_,
         ab_11__1_, ab_11__0_, ab_10__23_, ab_10__22_, ab_10__21_, ab_10__20_,
         ab_10__19_, ab_10__18_, ab_10__17_, ab_10__16_, ab_10__15_,
         ab_10__14_, ab_10__13_, ab_10__12_, ab_10__11_, ab_10__10_, ab_10__9_,
         ab_10__8_, ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_,
         ab_10__2_, ab_10__1_, ab_10__0_, ab_9__23_, ab_9__22_, ab_9__21_,
         ab_9__20_, ab_9__19_, ab_9__18_, ab_9__17_, ab_9__16_, ab_9__15_,
         ab_9__14_, ab_9__13_, ab_9__12_, ab_9__11_, ab_9__10_, ab_9__9_,
         ab_9__8_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_,
         ab_9__1_, ab_9__0_, ab_8__23_, ab_8__22_, ab_8__21_, ab_8__20_,
         ab_8__19_, ab_8__18_, ab_8__17_, ab_8__16_, ab_8__15_, ab_8__14_,
         ab_8__13_, ab_8__12_, ab_8__11_, ab_8__10_, ab_8__9_, ab_8__8_,
         ab_8__7_, ab_8__6_, ab_8__5_, ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_,
         ab_8__0_, ab_7__23_, ab_7__22_, ab_7__21_, ab_7__20_, ab_7__19_,
         ab_7__18_, ab_7__17_, ab_7__16_, ab_7__15_, ab_7__14_, ab_7__13_,
         ab_7__12_, ab_7__11_, ab_7__10_, ab_7__9_, ab_7__8_, ab_7__7_,
         ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_,
         ab_6__23_, ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_, ab_6__18_,
         ab_6__17_, ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_, ab_6__12_,
         ab_6__11_, ab_6__10_, ab_6__9_, ab_6__8_, ab_6__7_, ab_6__6_,
         ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_, ab_5__23_,
         ab_5__22_, ab_5__21_, ab_5__20_, ab_5__19_, ab_5__18_, ab_5__17_,
         ab_5__16_, ab_5__15_, ab_5__14_, ab_5__13_, ab_5__12_, ab_5__11_,
         ab_5__10_, ab_5__9_, ab_5__8_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_,
         ab_5__3_, ab_5__2_, ab_5__1_, ab_5__0_, ab_4__23_, ab_4__22_,
         ab_4__21_, ab_4__20_, ab_4__19_, ab_4__18_, ab_4__17_, ab_4__16_,
         ab_4__15_, ab_4__14_, ab_4__13_, ab_4__12_, ab_4__11_, ab_4__10_,
         ab_4__9_, ab_4__8_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_,
         ab_4__2_, ab_4__1_, ab_4__0_, ab_3__23_, ab_3__22_, ab_3__21_,
         ab_3__20_, ab_3__19_, ab_3__18_, ab_3__17_, ab_3__16_, ab_3__15_,
         ab_3__14_, ab_3__13_, ab_3__12_, ab_3__11_, ab_3__10_, ab_3__9_,
         ab_3__8_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_, ab_3__2_,
         ab_3__1_, ab_3__0_, ab_2__23_, ab_2__22_, ab_2__21_, ab_2__20_,
         ab_2__19_, ab_2__18_, ab_2__17_, ab_2__16_, ab_2__15_, ab_2__14_,
         ab_2__13_, ab_2__12_, ab_2__11_, ab_2__10_, ab_2__9_, ab_2__8_,
         ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_,
         ab_2__0_, ab_1__23_, ab_1__22_, ab_1__21_, ab_1__20_, ab_1__19_,
         ab_1__18_, ab_1__17_, ab_1__16_, ab_1__15_, ab_1__14_, ab_1__13_,
         ab_1__12_, ab_1__11_, ab_1__10_, ab_1__9_, ab_1__8_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_0__23_,
         ab_0__22_, ab_0__21_, ab_0__20_, ab_0__19_, ab_0__18_, ab_0__17_,
         ab_0__16_, ab_0__15_, ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_,
         ab_0__10_, ab_0__9_, ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_23__23_, CARRYB_23__22_, CARRYB_23__21_,
         CARRYB_23__20_, CARRYB_23__19_, CARRYB_23__18_, CARRYB_23__17_,
         CARRYB_23__16_, CARRYB_23__15_, CARRYB_23__14_, CARRYB_23__13_,
         CARRYB_23__12_, CARRYB_23__11_, CARRYB_23__10_, CARRYB_23__9_,
         CARRYB_23__8_, CARRYB_23__7_, CARRYB_23__6_, CARRYB_23__5_,
         CARRYB_23__4_, CARRYB_23__3_, CARRYB_23__2_, CARRYB_23__1_,
         CARRYB_23__0_, CARRYB_22__22_, CARRYB_22__21_, CARRYB_22__20_,
         CARRYB_22__19_, CARRYB_22__18_, CARRYB_22__17_, CARRYB_22__16_,
         CARRYB_22__15_, CARRYB_22__14_, CARRYB_22__13_, CARRYB_22__12_,
         CARRYB_22__11_, CARRYB_22__10_, CARRYB_22__9_, CARRYB_22__8_,
         CARRYB_22__7_, CARRYB_22__6_, CARRYB_22__5_, CARRYB_22__4_,
         CARRYB_22__3_, CARRYB_22__2_, CARRYB_22__1_, CARRYB_22__0_,
         CARRYB_21__22_, CARRYB_21__21_, CARRYB_21__20_, CARRYB_21__19_,
         CARRYB_21__18_, CARRYB_21__17_, CARRYB_21__16_, CARRYB_21__15_,
         CARRYB_21__14_, CARRYB_21__13_, CARRYB_21__12_, CARRYB_21__11_,
         CARRYB_21__10_, CARRYB_21__9_, CARRYB_21__8_, CARRYB_21__7_,
         CARRYB_21__6_, CARRYB_21__5_, CARRYB_21__4_, CARRYB_21__3_,
         CARRYB_21__2_, CARRYB_21__1_, CARRYB_21__0_, CARRYB_20__22_,
         CARRYB_20__21_, CARRYB_20__20_, CARRYB_20__19_, CARRYB_20__18_,
         CARRYB_20__17_, CARRYB_20__16_, CARRYB_20__15_, CARRYB_20__14_,
         CARRYB_20__13_, CARRYB_20__12_, CARRYB_20__11_, CARRYB_20__10_,
         CARRYB_20__9_, CARRYB_20__8_, CARRYB_20__7_, CARRYB_20__6_,
         CARRYB_20__5_, CARRYB_20__4_, CARRYB_20__3_, CARRYB_20__2_,
         CARRYB_20__1_, CARRYB_20__0_, CARRYB_19__22_, CARRYB_19__21_,
         CARRYB_19__20_, CARRYB_19__19_, CARRYB_19__18_, CARRYB_19__17_,
         CARRYB_19__16_, CARRYB_19__15_, CARRYB_19__14_, CARRYB_19__13_,
         CARRYB_19__12_, CARRYB_19__11_, CARRYB_19__10_, CARRYB_19__9_,
         CARRYB_19__8_, CARRYB_19__7_, CARRYB_19__6_, CARRYB_19__5_,
         CARRYB_19__4_, CARRYB_19__3_, CARRYB_19__2_, CARRYB_19__1_,
         CARRYB_19__0_, CARRYB_18__22_, CARRYB_18__21_, CARRYB_18__20_,
         CARRYB_18__19_, CARRYB_18__18_, CARRYB_18__17_, CARRYB_18__16_,
         CARRYB_18__15_, CARRYB_18__14_, CARRYB_18__13_, CARRYB_18__12_,
         CARRYB_18__11_, CARRYB_18__10_, CARRYB_18__9_, CARRYB_18__8_,
         CARRYB_18__7_, CARRYB_18__6_, CARRYB_18__5_, CARRYB_18__4_,
         CARRYB_18__3_, CARRYB_18__2_, CARRYB_18__1_, CARRYB_18__0_,
         CARRYB_17__22_, CARRYB_17__21_, CARRYB_17__20_, CARRYB_17__19_,
         CARRYB_17__18_, CARRYB_17__17_, CARRYB_17__16_, CARRYB_17__15_,
         CARRYB_17__14_, CARRYB_17__13_, CARRYB_17__12_, CARRYB_17__11_,
         CARRYB_17__10_, CARRYB_17__9_, CARRYB_17__8_, CARRYB_17__7_,
         CARRYB_17__6_, CARRYB_17__5_, CARRYB_17__4_, CARRYB_17__3_,
         CARRYB_17__2_, CARRYB_17__1_, CARRYB_17__0_, CARRYB_16__22_,
         CARRYB_16__21_, CARRYB_16__20_, CARRYB_16__19_, CARRYB_16__18_,
         CARRYB_16__17_, CARRYB_16__16_, CARRYB_16__15_, CARRYB_16__14_,
         CARRYB_16__13_, CARRYB_16__12_, CARRYB_16__11_, CARRYB_16__10_,
         CARRYB_16__9_, CARRYB_16__8_, CARRYB_16__7_, CARRYB_16__6_,
         CARRYB_16__5_, CARRYB_16__4_, CARRYB_16__3_, CARRYB_16__2_,
         CARRYB_16__1_, CARRYB_16__0_, CARRYB_15__22_, CARRYB_15__21_,
         CARRYB_15__20_, CARRYB_15__19_, CARRYB_15__18_, CARRYB_15__17_,
         CARRYB_15__16_, CARRYB_15__15_, CARRYB_15__14_, CARRYB_15__13_,
         CARRYB_15__12_, CARRYB_15__11_, CARRYB_15__10_, CARRYB_15__9_,
         CARRYB_15__8_, CARRYB_15__7_, CARRYB_15__6_, CARRYB_15__5_,
         CARRYB_15__4_, CARRYB_15__3_, CARRYB_15__2_, CARRYB_15__1_,
         CARRYB_15__0_, CARRYB_14__22_, CARRYB_14__21_, CARRYB_14__20_,
         CARRYB_14__19_, CARRYB_14__18_, CARRYB_14__17_, CARRYB_14__16_,
         CARRYB_14__15_, CARRYB_14__14_, CARRYB_14__13_, CARRYB_14__12_,
         CARRYB_14__11_, CARRYB_14__10_, CARRYB_14__9_, CARRYB_14__8_,
         CARRYB_14__7_, CARRYB_14__6_, CARRYB_14__5_, CARRYB_14__4_,
         CARRYB_14__3_, CARRYB_14__2_, CARRYB_14__1_, CARRYB_14__0_,
         CARRYB_13__22_, CARRYB_13__21_, CARRYB_13__20_, CARRYB_13__19_,
         CARRYB_13__18_, CARRYB_13__17_, CARRYB_13__16_, CARRYB_13__15_,
         CARRYB_13__14_, CARRYB_13__13_, CARRYB_13__12_, CARRYB_13__11_,
         CARRYB_13__10_, CARRYB_13__9_, CARRYB_13__8_, CARRYB_13__7_,
         CARRYB_13__6_, CARRYB_13__5_, CARRYB_13__4_, CARRYB_13__3_,
         CARRYB_13__2_, CARRYB_13__1_, CARRYB_13__0_, CARRYB_12__22_,
         CARRYB_12__21_, CARRYB_12__20_, CARRYB_12__19_, CARRYB_12__18_,
         CARRYB_12__17_, CARRYB_12__16_, CARRYB_12__15_, CARRYB_12__14_,
         CARRYB_12__13_, CARRYB_12__12_, CARRYB_12__11_, CARRYB_12__10_,
         CARRYB_12__9_, CARRYB_12__8_, CARRYB_12__7_, CARRYB_12__6_,
         CARRYB_12__5_, CARRYB_12__4_, CARRYB_12__3_, CARRYB_12__2_,
         CARRYB_12__1_, CARRYB_12__0_, CARRYB_11__22_, CARRYB_11__21_,
         CARRYB_11__20_, CARRYB_11__19_, CARRYB_11__18_, CARRYB_11__17_,
         CARRYB_11__16_, CARRYB_11__15_, CARRYB_11__14_, CARRYB_11__13_,
         CARRYB_11__12_, CARRYB_11__11_, CARRYB_11__10_, CARRYB_11__9_,
         CARRYB_11__8_, CARRYB_11__7_, CARRYB_11__6_, CARRYB_11__5_,
         CARRYB_11__4_, CARRYB_11__3_, CARRYB_11__2_, CARRYB_11__1_,
         CARRYB_11__0_, CARRYB_10__22_, CARRYB_10__21_, CARRYB_10__20_,
         CARRYB_10__19_, CARRYB_10__18_, CARRYB_10__17_, CARRYB_10__16_,
         CARRYB_10__15_, CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_,
         CARRYB_10__11_, CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_,
         CARRYB_10__7_, CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_,
         CARRYB_10__3_, CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_,
         CARRYB_9__22_, CARRYB_9__21_, CARRYB_9__20_, CARRYB_9__19_,
         CARRYB_9__18_, CARRYB_9__17_, CARRYB_9__16_, CARRYB_9__15_,
         CARRYB_9__14_, CARRYB_9__13_, CARRYB_9__12_, CARRYB_9__11_,
         CARRYB_9__10_, CARRYB_9__9_, CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_,
         CARRYB_9__5_, CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_,
         CARRYB_9__0_, CARRYB_8__22_, CARRYB_8__21_, CARRYB_8__20_,
         CARRYB_8__19_, CARRYB_8__18_, CARRYB_8__17_, CARRYB_8__16_,
         CARRYB_8__15_, CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_,
         CARRYB_8__11_, CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_,
         CARRYB_8__7_, CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_,
         CARRYB_8__2_, CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__22_,
         CARRYB_7__21_, CARRYB_7__20_, CARRYB_7__19_, CARRYB_7__18_,
         CARRYB_7__17_, CARRYB_7__16_, CARRYB_7__15_, CARRYB_7__14_,
         CARRYB_7__13_, CARRYB_7__12_, CARRYB_7__11_, CARRYB_7__10_,
         CARRYB_7__9_, CARRYB_7__8_, CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_,
         CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_,
         CARRYB_6__22_, CARRYB_6__21_, CARRYB_6__20_, CARRYB_6__19_,
         CARRYB_6__18_, CARRYB_6__17_, CARRYB_6__16_, CARRYB_6__15_,
         CARRYB_6__14_, CARRYB_6__13_, CARRYB_6__12_, CARRYB_6__11_,
         CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_, CARRYB_6__7_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__22_, CARRYB_5__21_, CARRYB_5__20_,
         CARRYB_5__19_, CARRYB_5__18_, CARRYB_5__17_, CARRYB_5__16_,
         CARRYB_5__15_, CARRYB_5__14_, CARRYB_5__13_, CARRYB_5__12_,
         CARRYB_5__11_, CARRYB_5__10_, CARRYB_5__9_, CARRYB_5__8_,
         CARRYB_5__7_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__22_,
         CARRYB_4__21_, CARRYB_4__20_, CARRYB_4__19_, CARRYB_4__18_,
         CARRYB_4__17_, CARRYB_4__16_, CARRYB_4__15_, CARRYB_4__14_,
         CARRYB_4__13_, CARRYB_4__12_, CARRYB_4__11_, CARRYB_4__10_,
         CARRYB_4__9_, CARRYB_4__8_, CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__22_, CARRYB_3__21_, CARRYB_3__20_, CARRYB_3__19_,
         CARRYB_3__18_, CARRYB_3__17_, CARRYB_3__16_, CARRYB_3__15_,
         CARRYB_3__14_, CARRYB_3__13_, CARRYB_3__12_, CARRYB_3__11_,
         CARRYB_3__10_, CARRYB_3__9_, CARRYB_3__8_, CARRYB_3__7_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__22_, CARRYB_2__21_, CARRYB_2__20_,
         CARRYB_2__19_, CARRYB_2__18_, CARRYB_2__17_, CARRYB_2__16_,
         CARRYB_2__15_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__22_,
         CARRYB_1__21_, CARRYB_1__20_, CARRYB_1__19_, CARRYB_1__18_,
         CARRYB_1__17_, CARRYB_1__16_, CARRYB_1__15_, CARRYB_1__14_,
         CARRYB_1__13_, CARRYB_1__12_, CARRYB_1__11_, CARRYB_1__10_,
         CARRYB_1__9_, CARRYB_1__8_, CARRYB_1__7_, CARRYB_1__6_, CARRYB_1__5_,
         CARRYB_1__4_, CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_,
         SUMB_23__23_, SUMB_23__22_, SUMB_23__21_, SUMB_23__20_, SUMB_23__19_,
         SUMB_23__18_, SUMB_23__17_, SUMB_23__16_, SUMB_23__15_, SUMB_23__14_,
         SUMB_23__13_, SUMB_23__12_, SUMB_23__11_, SUMB_23__10_, SUMB_23__9_,
         SUMB_23__8_, SUMB_23__7_, SUMB_23__6_, SUMB_23__5_, SUMB_23__4_,
         SUMB_23__3_, SUMB_23__2_, SUMB_23__1_, SUMB_23__0_, SUMB_22__22_,
         SUMB_22__21_, SUMB_22__20_, SUMB_22__19_, SUMB_22__18_, SUMB_22__17_,
         SUMB_22__16_, SUMB_22__15_, SUMB_22__14_, SUMB_22__13_, SUMB_22__12_,
         SUMB_22__11_, SUMB_22__10_, SUMB_22__9_, SUMB_22__8_, SUMB_22__7_,
         SUMB_22__6_, SUMB_22__5_, SUMB_22__4_, SUMB_22__3_, SUMB_22__2_,
         SUMB_22__1_, SUMB_21__22_, SUMB_21__21_, SUMB_21__20_, SUMB_21__19_,
         SUMB_21__18_, SUMB_21__17_, SUMB_21__16_, SUMB_21__15_, SUMB_21__14_,
         SUMB_21__13_, SUMB_21__12_, SUMB_21__11_, SUMB_21__10_, SUMB_21__9_,
         SUMB_21__8_, SUMB_21__7_, SUMB_21__6_, SUMB_21__5_, SUMB_21__4_,
         SUMB_21__3_, SUMB_21__2_, SUMB_21__1_, SUMB_20__22_, SUMB_20__21_,
         SUMB_20__20_, SUMB_20__19_, SUMB_20__18_, SUMB_20__17_, SUMB_20__16_,
         SUMB_20__15_, SUMB_20__14_, SUMB_20__13_, SUMB_20__12_, SUMB_20__11_,
         SUMB_20__10_, SUMB_20__9_, SUMB_20__8_, SUMB_20__7_, SUMB_20__6_,
         SUMB_20__5_, SUMB_20__4_, SUMB_20__3_, SUMB_20__2_, SUMB_20__1_,
         SUMB_19__22_, SUMB_19__21_, SUMB_19__20_, SUMB_19__19_, SUMB_19__18_,
         SUMB_19__17_, SUMB_19__16_, SUMB_19__15_, SUMB_19__14_, SUMB_19__13_,
         SUMB_19__12_, SUMB_19__11_, SUMB_19__10_, SUMB_19__9_, SUMB_19__8_,
         SUMB_19__7_, SUMB_19__6_, SUMB_19__5_, SUMB_19__4_, SUMB_19__3_,
         SUMB_19__2_, SUMB_19__1_, SUMB_18__22_, SUMB_18__21_, SUMB_18__20_,
         SUMB_18__19_, SUMB_18__18_, SUMB_18__17_, SUMB_18__16_, SUMB_18__15_,
         SUMB_18__14_, SUMB_18__13_, SUMB_18__12_, SUMB_18__11_, SUMB_18__10_,
         SUMB_18__9_, SUMB_18__8_, SUMB_18__7_, SUMB_18__6_, SUMB_18__5_,
         SUMB_18__4_, SUMB_18__3_, SUMB_18__2_, SUMB_18__1_, SUMB_17__22_,
         SUMB_17__21_, SUMB_17__20_, SUMB_17__19_, SUMB_17__18_, SUMB_17__17_,
         SUMB_17__16_, SUMB_17__15_, SUMB_17__14_, SUMB_17__13_, SUMB_17__12_,
         SUMB_17__11_, SUMB_17__10_, SUMB_17__9_, SUMB_17__8_, SUMB_17__7_,
         SUMB_17__6_, SUMB_17__5_, SUMB_17__4_, SUMB_17__3_, SUMB_17__2_,
         SUMB_17__1_, SUMB_16__22_, SUMB_16__21_, SUMB_16__20_, SUMB_16__19_,
         SUMB_16__18_, SUMB_16__17_, SUMB_16__16_, SUMB_16__15_, SUMB_16__14_,
         SUMB_16__13_, SUMB_16__12_, SUMB_16__11_, SUMB_16__10_, SUMB_16__9_,
         SUMB_16__8_, SUMB_16__7_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_,
         SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, SUMB_15__22_, SUMB_15__21_,
         SUMB_15__20_, SUMB_15__19_, SUMB_15__18_, SUMB_15__17_, SUMB_15__16_,
         SUMB_15__15_, SUMB_15__14_, SUMB_15__13_, SUMB_15__12_, SUMB_15__11_,
         SUMB_15__10_, SUMB_15__9_, SUMB_15__8_, SUMB_15__7_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_14__22_, SUMB_14__21_, SUMB_14__20_, SUMB_14__19_, SUMB_14__18_,
         SUMB_14__17_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_, SUMB_14__13_,
         SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_, SUMB_14__8_,
         SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_,
         SUMB_14__2_, SUMB_14__1_, SUMB_13__22_, SUMB_13__21_, SUMB_13__20_,
         SUMB_13__19_, SUMB_13__18_, SUMB_13__17_, SUMB_13__16_, SUMB_13__15_,
         SUMB_13__14_, SUMB_13__13_, SUMB_13__12_, SUMB_13__11_, SUMB_13__10_,
         SUMB_13__9_, SUMB_13__8_, SUMB_13__7_, SUMB_13__6_, SUMB_13__5_,
         SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_, SUMB_12__22_,
         SUMB_12__21_, SUMB_12__20_, SUMB_12__19_, SUMB_12__18_, SUMB_12__17_,
         SUMB_12__16_, SUMB_12__15_, SUMB_12__14_, SUMB_12__13_, SUMB_12__12_,
         SUMB_12__11_, SUMB_12__10_, SUMB_12__9_, SUMB_12__8_, SUMB_12__7_,
         SUMB_12__6_, SUMB_12__5_, SUMB_12__4_, SUMB_12__3_, SUMB_12__2_,
         SUMB_12__1_, SUMB_11__22_, SUMB_11__21_, SUMB_11__20_, SUMB_11__19_,
         SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_, SUMB_11__14_,
         SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_, SUMB_11__9_,
         SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_, SUMB_11__4_,
         SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__22_, SUMB_10__21_,
         SUMB_10__20_, SUMB_10__19_, SUMB_10__18_, SUMB_10__17_, SUMB_10__16_,
         SUMB_10__15_, SUMB_10__14_, SUMB_10__13_, SUMB_10__12_, SUMB_10__11_,
         SUMB_10__10_, SUMB_10__9_, SUMB_10__8_, SUMB_10__7_, SUMB_10__6_,
         SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_,
         SUMB_9__22_, SUMB_9__21_, SUMB_9__20_, SUMB_9__19_, SUMB_9__18_,
         SUMB_9__17_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_, SUMB_9__13_,
         SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_, SUMB_9__8_,
         SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_,
         SUMB_9__2_, SUMB_9__1_, SUMB_8__22_, SUMB_8__21_, SUMB_8__20_,
         SUMB_8__19_, SUMB_8__18_, SUMB_8__17_, SUMB_8__16_, SUMB_8__15_,
         SUMB_8__14_, SUMB_8__13_, SUMB_8__12_, SUMB_8__11_, SUMB_8__10_,
         SUMB_8__9_, SUMB_8__8_, SUMB_8__7_, SUMB_8__6_, SUMB_8__5_,
         SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_, SUMB_7__22_,
         SUMB_7__21_, SUMB_7__20_, SUMB_7__19_, SUMB_7__18_, SUMB_7__17_,
         SUMB_7__16_, SUMB_7__15_, SUMB_7__14_, SUMB_7__13_, SUMB_7__12_,
         SUMB_7__11_, SUMB_7__10_, SUMB_7__9_, SUMB_7__8_, SUMB_7__7_,
         SUMB_7__6_, SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_,
         SUMB_7__1_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_, SUMB_6__19_,
         SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_, SUMB_6__14_,
         SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_, SUMB_6__9_,
         SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_,
         SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__22_, SUMB_5__21_,
         SUMB_5__20_, SUMB_5__19_, SUMB_5__18_, SUMB_5__17_, SUMB_5__16_,
         SUMB_5__15_, SUMB_5__14_, SUMB_5__13_, SUMB_5__12_, SUMB_5__11_,
         SUMB_5__10_, SUMB_5__9_, SUMB_5__8_, SUMB_5__7_, SUMB_5__6_,
         SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_,
         SUMB_4__22_, SUMB_4__21_, SUMB_4__20_, SUMB_4__19_, SUMB_4__18_,
         SUMB_4__17_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_, SUMB_4__13_,
         SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_, SUMB_4__8_,
         SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_,
         SUMB_4__2_, SUMB_4__1_, SUMB_3__22_, SUMB_3__21_, SUMB_3__20_,
         SUMB_3__19_, SUMB_3__18_, SUMB_3__17_, SUMB_3__16_, SUMB_3__15_,
         SUMB_3__14_, SUMB_3__13_, SUMB_3__12_, SUMB_3__11_, SUMB_3__10_,
         SUMB_3__9_, SUMB_3__8_, SUMB_3__7_, SUMB_3__6_, SUMB_3__5_,
         SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_, SUMB_2__22_,
         SUMB_2__21_, SUMB_2__20_, SUMB_2__19_, SUMB_2__18_, SUMB_2__17_,
         SUMB_2__16_, SUMB_2__15_, SUMB_2__14_, SUMB_2__13_, SUMB_2__12_,
         SUMB_2__11_, SUMB_2__10_, SUMB_2__9_, SUMB_2__8_, SUMB_2__7_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__22_, SUMB_1__21_, SUMB_1__20_, SUMB_1__19_,
         SUMB_1__18_, SUMB_1__17_, SUMB_1__16_, SUMB_1__15_, SUMB_1__14_,
         SUMB_1__13_, SUMB_1__12_, SUMB_1__11_, SUMB_1__10_, SUMB_1__9_,
         SUMB_1__8_, SUMB_1__7_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_,
         SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, QA, QB, A1_45_, A1_44_, A1_43_,
         A1_42_, A1_41_, A1_40_, A1_39_, A1_38_, A1_37_, A1_36_, A1_35_,
         A1_34_, A1_33_, A1_32_, A1_31_, A1_30_, A1_29_, A1_28_, A1_27_,
         A1_26_, A1_25_, A1_24_, A1_23_, A1_22_, A1_21_, A1_20_, A1_19_,
         A1_18_, A1_17_, A1_16_, A1_15_, A1_14_, A1_13_, A1_12_, A1_11_,
         A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_,
         A1_0_, A2_45_, A2_44_, A2_43_, A2_42_, A2_41_, A2_40_, A2_39_, A2_38_,
         A2_37_, A2_36_, A2_35_, A2_34_, A2_33_, A2_32_, A2_31_, A2_30_,
         A2_29_, A2_28_, A2_27_, A2_26_, A2_25_, A2_24_, A2_23_, A2_22_, n1,
         n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21;

  FA_X1 S14_23_0 ( .A(A[23]), .B(B[23]), .CI(SUMB_23__0_), .CO(A2_22_), .S(
        A1_21_) );
  FA_X1 S4_0 ( .A(ab_23__0_), .B(CARRYB_22__0_), .CI(SUMB_22__1_), .CO(
        CARRYB_23__0_), .S(SUMB_23__0_) );
  FA_X1 S4_1 ( .A(ab_23__1_), .B(CARRYB_22__1_), .CI(SUMB_22__2_), .CO(
        CARRYB_23__1_), .S(SUMB_23__1_) );
  FA_X1 S4_2 ( .A(ab_23__2_), .B(CARRYB_22__2_), .CI(SUMB_22__3_), .CO(
        CARRYB_23__2_), .S(SUMB_23__2_) );
  FA_X1 S4_3 ( .A(ab_23__3_), .B(CARRYB_22__3_), .CI(SUMB_22__4_), .CO(
        CARRYB_23__3_), .S(SUMB_23__3_) );
  FA_X1 S4_4 ( .A(ab_23__4_), .B(CARRYB_22__4_), .CI(SUMB_22__5_), .CO(
        CARRYB_23__4_), .S(SUMB_23__4_) );
  FA_X1 S4_5 ( .A(ab_23__5_), .B(CARRYB_22__5_), .CI(SUMB_22__6_), .CO(
        CARRYB_23__5_), .S(SUMB_23__5_) );
  FA_X1 S4_6 ( .A(ab_23__6_), .B(CARRYB_22__6_), .CI(SUMB_22__7_), .CO(
        CARRYB_23__6_), .S(SUMB_23__6_) );
  FA_X1 S4_7 ( .A(ab_23__7_), .B(CARRYB_22__7_), .CI(SUMB_22__8_), .CO(
        CARRYB_23__7_), .S(SUMB_23__7_) );
  FA_X1 S4_8 ( .A(ab_23__8_), .B(CARRYB_22__8_), .CI(SUMB_22__9_), .CO(
        CARRYB_23__8_), .S(SUMB_23__8_) );
  FA_X1 S4_9 ( .A(ab_23__9_), .B(CARRYB_22__9_), .CI(SUMB_22__10_), .CO(
        CARRYB_23__9_), .S(SUMB_23__9_) );
  FA_X1 S4_10 ( .A(ab_23__10_), .B(CARRYB_22__10_), .CI(SUMB_22__11_), .CO(
        CARRYB_23__10_), .S(SUMB_23__10_) );
  FA_X1 S4_11 ( .A(ab_23__11_), .B(CARRYB_22__11_), .CI(SUMB_22__12_), .CO(
        CARRYB_23__11_), .S(SUMB_23__11_) );
  FA_X1 S4_12 ( .A(ab_23__12_), .B(CARRYB_22__12_), .CI(SUMB_22__13_), .CO(
        CARRYB_23__12_), .S(SUMB_23__12_) );
  FA_X1 S4_13 ( .A(ab_23__13_), .B(CARRYB_22__13_), .CI(SUMB_22__14_), .CO(
        CARRYB_23__13_), .S(SUMB_23__13_) );
  FA_X1 S4_14 ( .A(ab_23__14_), .B(CARRYB_22__14_), .CI(SUMB_22__15_), .CO(
        CARRYB_23__14_), .S(SUMB_23__14_) );
  FA_X1 S4_15 ( .A(ab_23__15_), .B(CARRYB_22__15_), .CI(SUMB_22__16_), .CO(
        CARRYB_23__15_), .S(SUMB_23__15_) );
  FA_X1 S4_16 ( .A(ab_23__16_), .B(CARRYB_22__16_), .CI(SUMB_22__17_), .CO(
        CARRYB_23__16_), .S(SUMB_23__16_) );
  FA_X1 S4_17 ( .A(ab_23__17_), .B(CARRYB_22__17_), .CI(SUMB_22__18_), .CO(
        CARRYB_23__17_), .S(SUMB_23__17_) );
  FA_X1 S4_18 ( .A(ab_23__18_), .B(CARRYB_22__18_), .CI(SUMB_22__19_), .CO(
        CARRYB_23__18_), .S(SUMB_23__18_) );
  FA_X1 S4_19 ( .A(ab_23__19_), .B(CARRYB_22__19_), .CI(SUMB_22__20_), .CO(
        CARRYB_23__19_), .S(SUMB_23__19_) );
  FA_X1 S4_20 ( .A(ab_23__20_), .B(CARRYB_22__20_), .CI(SUMB_22__21_), .CO(
        CARRYB_23__20_), .S(SUMB_23__20_) );
  FA_X1 S4_21 ( .A(ab_23__21_), .B(CARRYB_22__21_), .CI(SUMB_22__22_), .CO(
        CARRYB_23__21_), .S(SUMB_23__21_) );
  FA_X1 S5_22 ( .A(ab_23__22_), .B(CARRYB_22__22_), .CI(ab_22__23_), .CO(
        CARRYB_23__22_), .S(SUMB_23__22_) );
  FA_X1 S14_23 ( .A(n3), .B(n1), .CI(ab_23__23_), .CO(CARRYB_23__23_), .S(
        SUMB_23__23_) );
  FA_X1 S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), .CO(
        CARRYB_22__0_), .S(A1_20_) );
  FA_X1 S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), .CO(
        CARRYB_22__1_), .S(SUMB_22__1_) );
  FA_X1 S2_22_2 ( .A(ab_22__2_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), .CO(
        CARRYB_22__2_), .S(SUMB_22__2_) );
  FA_X1 S2_22_3 ( .A(ab_22__3_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), .CO(
        CARRYB_22__3_), .S(SUMB_22__3_) );
  FA_X1 S2_22_4 ( .A(ab_22__4_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), .CO(
        CARRYB_22__4_), .S(SUMB_22__4_) );
  FA_X1 S2_22_5 ( .A(ab_22__5_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), .CO(
        CARRYB_22__5_), .S(SUMB_22__5_) );
  FA_X1 S2_22_6 ( .A(ab_22__6_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), .CO(
        CARRYB_22__6_), .S(SUMB_22__6_) );
  FA_X1 S2_22_7 ( .A(ab_22__7_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), .CO(
        CARRYB_22__7_), .S(SUMB_22__7_) );
  FA_X1 S2_22_8 ( .A(ab_22__8_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), .CO(
        CARRYB_22__8_), .S(SUMB_22__8_) );
  FA_X1 S2_22_9 ( .A(ab_22__9_), .B(CARRYB_21__9_), .CI(SUMB_21__10_), .CO(
        CARRYB_22__9_), .S(SUMB_22__9_) );
  FA_X1 S2_22_10 ( .A(ab_22__10_), .B(CARRYB_21__10_), .CI(SUMB_21__11_), .CO(
        CARRYB_22__10_), .S(SUMB_22__10_) );
  FA_X1 S2_22_11 ( .A(ab_22__11_), .B(CARRYB_21__11_), .CI(SUMB_21__12_), .CO(
        CARRYB_22__11_), .S(SUMB_22__11_) );
  FA_X1 S2_22_12 ( .A(ab_22__12_), .B(CARRYB_21__12_), .CI(SUMB_21__13_), .CO(
        CARRYB_22__12_), .S(SUMB_22__12_) );
  FA_X1 S2_22_13 ( .A(ab_22__13_), .B(CARRYB_21__13_), .CI(SUMB_21__14_), .CO(
        CARRYB_22__13_), .S(SUMB_22__13_) );
  FA_X1 S2_22_14 ( .A(ab_22__14_), .B(CARRYB_21__14_), .CI(SUMB_21__15_), .CO(
        CARRYB_22__14_), .S(SUMB_22__14_) );
  FA_X1 S2_22_15 ( .A(ab_22__15_), .B(CARRYB_21__15_), .CI(SUMB_21__16_), .CO(
        CARRYB_22__15_), .S(SUMB_22__15_) );
  FA_X1 S2_22_16 ( .A(ab_22__16_), .B(CARRYB_21__16_), .CI(SUMB_21__17_), .CO(
        CARRYB_22__16_), .S(SUMB_22__16_) );
  FA_X1 S2_22_17 ( .A(ab_22__17_), .B(CARRYB_21__17_), .CI(SUMB_21__18_), .CO(
        CARRYB_22__17_), .S(SUMB_22__17_) );
  FA_X1 S2_22_18 ( .A(ab_22__18_), .B(CARRYB_21__18_), .CI(SUMB_21__19_), .CO(
        CARRYB_22__18_), .S(SUMB_22__18_) );
  FA_X1 S2_22_19 ( .A(ab_22__19_), .B(CARRYB_21__19_), .CI(SUMB_21__20_), .CO(
        CARRYB_22__19_), .S(SUMB_22__19_) );
  FA_X1 S2_22_20 ( .A(ab_22__20_), .B(CARRYB_21__20_), .CI(SUMB_21__21_), .CO(
        CARRYB_22__20_), .S(SUMB_22__20_) );
  FA_X1 S2_22_21 ( .A(ab_22__21_), .B(CARRYB_21__21_), .CI(SUMB_21__22_), .CO(
        CARRYB_22__21_), .S(SUMB_22__21_) );
  FA_X1 S3_22_22 ( .A(ab_22__22_), .B(CARRYB_21__22_), .CI(ab_21__23_), .CO(
        CARRYB_22__22_), .S(SUMB_22__22_) );
  FA_X1 S1_21_0 ( .A(ab_21__0_), .B(CARRYB_20__0_), .CI(SUMB_20__1_), .CO(
        CARRYB_21__0_), .S(A1_19_) );
  FA_X1 S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), .CO(
        CARRYB_21__1_), .S(SUMB_21__1_) );
  FA_X1 S2_21_2 ( .A(ab_21__2_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), .CO(
        CARRYB_21__2_), .S(SUMB_21__2_) );
  FA_X1 S2_21_3 ( .A(ab_21__3_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), .CO(
        CARRYB_21__3_), .S(SUMB_21__3_) );
  FA_X1 S2_21_4 ( .A(ab_21__4_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), .CO(
        CARRYB_21__4_), .S(SUMB_21__4_) );
  FA_X1 S2_21_5 ( .A(ab_21__5_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), .CO(
        CARRYB_21__5_), .S(SUMB_21__5_) );
  FA_X1 S2_21_6 ( .A(ab_21__6_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), .CO(
        CARRYB_21__6_), .S(SUMB_21__6_) );
  FA_X1 S2_21_7 ( .A(ab_21__7_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), .CO(
        CARRYB_21__7_), .S(SUMB_21__7_) );
  FA_X1 S2_21_8 ( .A(ab_21__8_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), .CO(
        CARRYB_21__8_), .S(SUMB_21__8_) );
  FA_X1 S2_21_9 ( .A(ab_21__9_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), .CO(
        CARRYB_21__9_), .S(SUMB_21__9_) );
  FA_X1 S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .CI(SUMB_20__11_), .CO(
        CARRYB_21__10_), .S(SUMB_21__10_) );
  FA_X1 S2_21_11 ( .A(ab_21__11_), .B(CARRYB_20__11_), .CI(SUMB_20__12_), .CO(
        CARRYB_21__11_), .S(SUMB_21__11_) );
  FA_X1 S2_21_12 ( .A(ab_21__12_), .B(CARRYB_20__12_), .CI(SUMB_20__13_), .CO(
        CARRYB_21__12_), .S(SUMB_21__12_) );
  FA_X1 S2_21_13 ( .A(ab_21__13_), .B(CARRYB_20__13_), .CI(SUMB_20__14_), .CO(
        CARRYB_21__13_), .S(SUMB_21__13_) );
  FA_X1 S2_21_14 ( .A(ab_21__14_), .B(CARRYB_20__14_), .CI(SUMB_20__15_), .CO(
        CARRYB_21__14_), .S(SUMB_21__14_) );
  FA_X1 S2_21_15 ( .A(ab_21__15_), .B(CARRYB_20__15_), .CI(SUMB_20__16_), .CO(
        CARRYB_21__15_), .S(SUMB_21__15_) );
  FA_X1 S2_21_16 ( .A(ab_21__16_), .B(CARRYB_20__16_), .CI(SUMB_20__17_), .CO(
        CARRYB_21__16_), .S(SUMB_21__16_) );
  FA_X1 S2_21_17 ( .A(ab_21__17_), .B(CARRYB_20__17_), .CI(SUMB_20__18_), .CO(
        CARRYB_21__17_), .S(SUMB_21__17_) );
  FA_X1 S2_21_18 ( .A(ab_21__18_), .B(CARRYB_20__18_), .CI(SUMB_20__19_), .CO(
        CARRYB_21__18_), .S(SUMB_21__18_) );
  FA_X1 S2_21_19 ( .A(ab_21__19_), .B(CARRYB_20__19_), .CI(SUMB_20__20_), .CO(
        CARRYB_21__19_), .S(SUMB_21__19_) );
  FA_X1 S2_21_20 ( .A(ab_21__20_), .B(CARRYB_20__20_), .CI(SUMB_20__21_), .CO(
        CARRYB_21__20_), .S(SUMB_21__20_) );
  FA_X1 S2_21_21 ( .A(ab_21__21_), .B(CARRYB_20__21_), .CI(SUMB_20__22_), .CO(
        CARRYB_21__21_), .S(SUMB_21__21_) );
  FA_X1 S3_21_22 ( .A(ab_21__22_), .B(CARRYB_20__22_), .CI(ab_20__23_), .CO(
        CARRYB_21__22_), .S(SUMB_21__22_) );
  FA_X1 S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), .CO(
        CARRYB_20__0_), .S(A1_18_) );
  FA_X1 S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), .CO(
        CARRYB_20__1_), .S(SUMB_20__1_) );
  FA_X1 S2_20_2 ( .A(ab_20__2_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), .CO(
        CARRYB_20__2_), .S(SUMB_20__2_) );
  FA_X1 S2_20_3 ( .A(ab_20__3_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), .CO(
        CARRYB_20__3_), .S(SUMB_20__3_) );
  FA_X1 S2_20_4 ( .A(ab_20__4_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), .CO(
        CARRYB_20__4_), .S(SUMB_20__4_) );
  FA_X1 S2_20_5 ( .A(ab_20__5_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), .CO(
        CARRYB_20__5_), .S(SUMB_20__5_) );
  FA_X1 S2_20_6 ( .A(ab_20__6_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), .CO(
        CARRYB_20__6_), .S(SUMB_20__6_) );
  FA_X1 S2_20_7 ( .A(ab_20__7_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), .CO(
        CARRYB_20__7_), .S(SUMB_20__7_) );
  FA_X1 S2_20_8 ( .A(ab_20__8_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), .CO(
        CARRYB_20__8_), .S(SUMB_20__8_) );
  FA_X1 S2_20_9 ( .A(ab_20__9_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), .CO(
        CARRYB_20__9_), .S(SUMB_20__9_) );
  FA_X1 S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), .CO(
        CARRYB_20__10_), .S(SUMB_20__10_) );
  FA_X1 S2_20_11 ( .A(ab_20__11_), .B(CARRYB_19__11_), .CI(SUMB_19__12_), .CO(
        CARRYB_20__11_), .S(SUMB_20__11_) );
  FA_X1 S2_20_12 ( .A(ab_20__12_), .B(CARRYB_19__12_), .CI(SUMB_19__13_), .CO(
        CARRYB_20__12_), .S(SUMB_20__12_) );
  FA_X1 S2_20_13 ( .A(ab_20__13_), .B(CARRYB_19__13_), .CI(SUMB_19__14_), .CO(
        CARRYB_20__13_), .S(SUMB_20__13_) );
  FA_X1 S2_20_14 ( .A(ab_20__14_), .B(CARRYB_19__14_), .CI(SUMB_19__15_), .CO(
        CARRYB_20__14_), .S(SUMB_20__14_) );
  FA_X1 S2_20_15 ( .A(ab_20__15_), .B(CARRYB_19__15_), .CI(SUMB_19__16_), .CO(
        CARRYB_20__15_), .S(SUMB_20__15_) );
  FA_X1 S2_20_16 ( .A(ab_20__16_), .B(CARRYB_19__16_), .CI(SUMB_19__17_), .CO(
        CARRYB_20__16_), .S(SUMB_20__16_) );
  FA_X1 S2_20_17 ( .A(ab_20__17_), .B(CARRYB_19__17_), .CI(SUMB_19__18_), .CO(
        CARRYB_20__17_), .S(SUMB_20__17_) );
  FA_X1 S2_20_18 ( .A(ab_20__18_), .B(CARRYB_19__18_), .CI(SUMB_19__19_), .CO(
        CARRYB_20__18_), .S(SUMB_20__18_) );
  FA_X1 S2_20_19 ( .A(ab_20__19_), .B(CARRYB_19__19_), .CI(SUMB_19__20_), .CO(
        CARRYB_20__19_), .S(SUMB_20__19_) );
  FA_X1 S2_20_20 ( .A(ab_20__20_), .B(CARRYB_19__20_), .CI(SUMB_19__21_), .CO(
        CARRYB_20__20_), .S(SUMB_20__20_) );
  FA_X1 S2_20_21 ( .A(ab_20__21_), .B(CARRYB_19__21_), .CI(SUMB_19__22_), .CO(
        CARRYB_20__21_), .S(SUMB_20__21_) );
  FA_X1 S3_20_22 ( .A(ab_20__22_), .B(CARRYB_19__22_), .CI(ab_19__23_), .CO(
        CARRYB_20__22_), .S(SUMB_20__22_) );
  FA_X1 S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), .CO(
        CARRYB_19__0_), .S(A1_17_) );
  FA_X1 S2_19_1 ( .A(ab_19__1_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), .CO(
        CARRYB_19__1_), .S(SUMB_19__1_) );
  FA_X1 S2_19_2 ( .A(ab_19__2_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), .CO(
        CARRYB_19__2_), .S(SUMB_19__2_) );
  FA_X1 S2_19_3 ( .A(ab_19__3_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), .CO(
        CARRYB_19__3_), .S(SUMB_19__3_) );
  FA_X1 S2_19_4 ( .A(ab_19__4_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), .CO(
        CARRYB_19__4_), .S(SUMB_19__4_) );
  FA_X1 S2_19_5 ( .A(ab_19__5_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), .CO(
        CARRYB_19__5_), .S(SUMB_19__5_) );
  FA_X1 S2_19_6 ( .A(ab_19__6_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), .CO(
        CARRYB_19__6_), .S(SUMB_19__6_) );
  FA_X1 S2_19_7 ( .A(ab_19__7_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), .CO(
        CARRYB_19__7_), .S(SUMB_19__7_) );
  FA_X1 S2_19_8 ( .A(ab_19__8_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), .CO(
        CARRYB_19__8_), .S(SUMB_19__8_) );
  FA_X1 S2_19_9 ( .A(ab_19__9_), .B(CARRYB_18__9_), .CI(SUMB_18__10_), .CO(
        CARRYB_19__9_), .S(SUMB_19__9_) );
  FA_X1 S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), .CO(
        CARRYB_19__10_), .S(SUMB_19__10_) );
  FA_X1 S2_19_11 ( .A(ab_19__11_), .B(CARRYB_18__11_), .CI(SUMB_18__12_), .CO(
        CARRYB_19__11_), .S(SUMB_19__11_) );
  FA_X1 S2_19_12 ( .A(ab_19__12_), .B(CARRYB_18__12_), .CI(SUMB_18__13_), .CO(
        CARRYB_19__12_), .S(SUMB_19__12_) );
  FA_X1 S2_19_13 ( .A(ab_19__13_), .B(CARRYB_18__13_), .CI(SUMB_18__14_), .CO(
        CARRYB_19__13_), .S(SUMB_19__13_) );
  FA_X1 S2_19_14 ( .A(ab_19__14_), .B(CARRYB_18__14_), .CI(SUMB_18__15_), .CO(
        CARRYB_19__14_), .S(SUMB_19__14_) );
  FA_X1 S2_19_15 ( .A(ab_19__15_), .B(CARRYB_18__15_), .CI(SUMB_18__16_), .CO(
        CARRYB_19__15_), .S(SUMB_19__15_) );
  FA_X1 S2_19_16 ( .A(ab_19__16_), .B(CARRYB_18__16_), .CI(SUMB_18__17_), .CO(
        CARRYB_19__16_), .S(SUMB_19__16_) );
  FA_X1 S2_19_17 ( .A(ab_19__17_), .B(CARRYB_18__17_), .CI(SUMB_18__18_), .CO(
        CARRYB_19__17_), .S(SUMB_19__17_) );
  FA_X1 S2_19_18 ( .A(ab_19__18_), .B(CARRYB_18__18_), .CI(SUMB_18__19_), .CO(
        CARRYB_19__18_), .S(SUMB_19__18_) );
  FA_X1 S2_19_19 ( .A(ab_19__19_), .B(CARRYB_18__19_), .CI(SUMB_18__20_), .CO(
        CARRYB_19__19_), .S(SUMB_19__19_) );
  FA_X1 S2_19_20 ( .A(ab_19__20_), .B(CARRYB_18__20_), .CI(SUMB_18__21_), .CO(
        CARRYB_19__20_), .S(SUMB_19__20_) );
  FA_X1 S2_19_21 ( .A(ab_19__21_), .B(CARRYB_18__21_), .CI(SUMB_18__22_), .CO(
        CARRYB_19__21_), .S(SUMB_19__21_) );
  FA_X1 S3_19_22 ( .A(ab_19__22_), .B(CARRYB_18__22_), .CI(ab_18__23_), .CO(
        CARRYB_19__22_), .S(SUMB_19__22_) );
  FA_X1 S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), .CO(
        CARRYB_18__0_), .S(A1_16_) );
  FA_X1 S2_18_1 ( .A(ab_18__1_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), .CO(
        CARRYB_18__1_), .S(SUMB_18__1_) );
  FA_X1 S2_18_2 ( .A(ab_18__2_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), .CO(
        CARRYB_18__2_), .S(SUMB_18__2_) );
  FA_X1 S2_18_3 ( .A(ab_18__3_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), .CO(
        CARRYB_18__3_), .S(SUMB_18__3_) );
  FA_X1 S2_18_4 ( .A(ab_18__4_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), .CO(
        CARRYB_18__4_), .S(SUMB_18__4_) );
  FA_X1 S2_18_5 ( .A(ab_18__5_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), .CO(
        CARRYB_18__5_), .S(SUMB_18__5_) );
  FA_X1 S2_18_6 ( .A(ab_18__6_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), .CO(
        CARRYB_18__6_), .S(SUMB_18__6_) );
  FA_X1 S2_18_7 ( .A(ab_18__7_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), .CO(
        CARRYB_18__7_), .S(SUMB_18__7_) );
  FA_X1 S2_18_8 ( .A(ab_18__8_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), .CO(
        CARRYB_18__8_), .S(SUMB_18__8_) );
  FA_X1 S2_18_9 ( .A(ab_18__9_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), .CO(
        CARRYB_18__9_), .S(SUMB_18__9_) );
  FA_X1 S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), .CO(
        CARRYB_18__10_), .S(SUMB_18__10_) );
  FA_X1 S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), .CO(
        CARRYB_18__11_), .S(SUMB_18__11_) );
  FA_X1 S2_18_12 ( .A(ab_18__12_), .B(CARRYB_17__12_), .CI(SUMB_17__13_), .CO(
        CARRYB_18__12_), .S(SUMB_18__12_) );
  FA_X1 S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .CI(SUMB_17__14_), .CO(
        CARRYB_18__13_), .S(SUMB_18__13_) );
  FA_X1 S2_18_14 ( .A(ab_18__14_), .B(CARRYB_17__14_), .CI(SUMB_17__15_), .CO(
        CARRYB_18__14_), .S(SUMB_18__14_) );
  FA_X1 S2_18_15 ( .A(ab_18__15_), .B(CARRYB_17__15_), .CI(SUMB_17__16_), .CO(
        CARRYB_18__15_), .S(SUMB_18__15_) );
  FA_X1 S2_18_16 ( .A(ab_18__16_), .B(CARRYB_17__16_), .CI(SUMB_17__17_), .CO(
        CARRYB_18__16_), .S(SUMB_18__16_) );
  FA_X1 S2_18_17 ( .A(ab_18__17_), .B(CARRYB_17__17_), .CI(SUMB_17__18_), .CO(
        CARRYB_18__17_), .S(SUMB_18__17_) );
  FA_X1 S2_18_18 ( .A(ab_18__18_), .B(CARRYB_17__18_), .CI(SUMB_17__19_), .CO(
        CARRYB_18__18_), .S(SUMB_18__18_) );
  FA_X1 S2_18_19 ( .A(ab_18__19_), .B(CARRYB_17__19_), .CI(SUMB_17__20_), .CO(
        CARRYB_18__19_), .S(SUMB_18__19_) );
  FA_X1 S2_18_20 ( .A(ab_18__20_), .B(CARRYB_17__20_), .CI(SUMB_17__21_), .CO(
        CARRYB_18__20_), .S(SUMB_18__20_) );
  FA_X1 S2_18_21 ( .A(ab_18__21_), .B(CARRYB_17__21_), .CI(SUMB_17__22_), .CO(
        CARRYB_18__21_), .S(SUMB_18__21_) );
  FA_X1 S3_18_22 ( .A(ab_18__22_), .B(CARRYB_17__22_), .CI(ab_17__23_), .CO(
        CARRYB_18__22_), .S(SUMB_18__22_) );
  FA_X1 S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), .CO(
        CARRYB_17__0_), .S(A1_15_) );
  FA_X1 S2_17_1 ( .A(ab_17__1_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), .CO(
        CARRYB_17__1_), .S(SUMB_17__1_) );
  FA_X1 S2_17_2 ( .A(ab_17__2_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), .CO(
        CARRYB_17__2_), .S(SUMB_17__2_) );
  FA_X1 S2_17_3 ( .A(ab_17__3_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), .CO(
        CARRYB_17__3_), .S(SUMB_17__3_) );
  FA_X1 S2_17_4 ( .A(ab_17__4_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), .CO(
        CARRYB_17__4_), .S(SUMB_17__4_) );
  FA_X1 S2_17_5 ( .A(ab_17__5_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), .CO(
        CARRYB_17__5_), .S(SUMB_17__5_) );
  FA_X1 S2_17_6 ( .A(ab_17__6_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), .CO(
        CARRYB_17__6_), .S(SUMB_17__6_) );
  FA_X1 S2_17_7 ( .A(ab_17__7_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), .CO(
        CARRYB_17__7_), .S(SUMB_17__7_) );
  FA_X1 S2_17_8 ( .A(ab_17__8_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), .CO(
        CARRYB_17__8_), .S(SUMB_17__8_) );
  FA_X1 S2_17_9 ( .A(ab_17__9_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), .CO(
        CARRYB_17__9_), .S(SUMB_17__9_) );
  FA_X1 S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), .CO(
        CARRYB_17__10_), .S(SUMB_17__10_) );
  FA_X1 S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), .CO(
        CARRYB_17__11_), .S(SUMB_17__11_) );
  FA_X1 S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), .CO(
        CARRYB_17__12_), .S(SUMB_17__12_) );
  FA_X1 S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), .CO(
        CARRYB_17__13_), .S(SUMB_17__13_) );
  FA_X1 S2_17_14 ( .A(ab_17__14_), .B(CARRYB_16__14_), .CI(SUMB_16__15_), .CO(
        CARRYB_17__14_), .S(SUMB_17__14_) );
  FA_X1 S2_17_15 ( .A(ab_17__15_), .B(CARRYB_16__15_), .CI(SUMB_16__16_), .CO(
        CARRYB_17__15_), .S(SUMB_17__15_) );
  FA_X1 S2_17_16 ( .A(ab_17__16_), .B(CARRYB_16__16_), .CI(SUMB_16__17_), .CO(
        CARRYB_17__16_), .S(SUMB_17__16_) );
  FA_X1 S2_17_17 ( .A(ab_17__17_), .B(CARRYB_16__17_), .CI(SUMB_16__18_), .CO(
        CARRYB_17__17_), .S(SUMB_17__17_) );
  FA_X1 S2_17_18 ( .A(ab_17__18_), .B(CARRYB_16__18_), .CI(SUMB_16__19_), .CO(
        CARRYB_17__18_), .S(SUMB_17__18_) );
  FA_X1 S2_17_19 ( .A(ab_17__19_), .B(CARRYB_16__19_), .CI(SUMB_16__20_), .CO(
        CARRYB_17__19_), .S(SUMB_17__19_) );
  FA_X1 S2_17_20 ( .A(ab_17__20_), .B(CARRYB_16__20_), .CI(SUMB_16__21_), .CO(
        CARRYB_17__20_), .S(SUMB_17__20_) );
  FA_X1 S2_17_21 ( .A(ab_17__21_), .B(CARRYB_16__21_), .CI(SUMB_16__22_), .CO(
        CARRYB_17__21_), .S(SUMB_17__21_) );
  FA_X1 S3_17_22 ( .A(ab_17__22_), .B(CARRYB_16__22_), .CI(ab_16__23_), .CO(
        CARRYB_17__22_), .S(SUMB_17__22_) );
  FA_X1 S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(A1_14_) );
  FA_X1 S2_16_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  FA_X1 S2_16_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  FA_X1 S2_16_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  FA_X1 S2_16_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  FA_X1 S2_16_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  FA_X1 S2_16_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  FA_X1 S2_16_7 ( .A(ab_16__7_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), .CO(
        CARRYB_16__7_), .S(SUMB_16__7_) );
  FA_X1 S2_16_8 ( .A(ab_16__8_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), .CO(
        CARRYB_16__8_), .S(SUMB_16__8_) );
  FA_X1 S2_16_9 ( .A(ab_16__9_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), .CO(
        CARRYB_16__9_), .S(SUMB_16__9_) );
  FA_X1 S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), .CO(
        CARRYB_16__10_), .S(SUMB_16__10_) );
  FA_X1 S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), .CO(
        CARRYB_16__11_), .S(SUMB_16__11_) );
  FA_X1 S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), .CO(
        CARRYB_16__12_), .S(SUMB_16__12_) );
  FA_X1 S2_16_13 ( .A(ab_16__13_), .B(CARRYB_15__13_), .CI(SUMB_15__14_), .CO(
        CARRYB_16__13_), .S(SUMB_16__13_) );
  FA_X1 S2_16_14 ( .A(ab_16__14_), .B(CARRYB_15__14_), .CI(SUMB_15__15_), .CO(
        CARRYB_16__14_), .S(SUMB_16__14_) );
  FA_X1 S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .CI(SUMB_15__16_), .CO(
        CARRYB_16__15_), .S(SUMB_16__15_) );
  FA_X1 S2_16_16 ( .A(ab_16__16_), .B(CARRYB_15__16_), .CI(SUMB_15__17_), .CO(
        CARRYB_16__16_), .S(SUMB_16__16_) );
  FA_X1 S2_16_17 ( .A(ab_16__17_), .B(CARRYB_15__17_), .CI(SUMB_15__18_), .CO(
        CARRYB_16__17_), .S(SUMB_16__17_) );
  FA_X1 S2_16_18 ( .A(ab_16__18_), .B(CARRYB_15__18_), .CI(SUMB_15__19_), .CO(
        CARRYB_16__18_), .S(SUMB_16__18_) );
  FA_X1 S2_16_19 ( .A(ab_16__19_), .B(CARRYB_15__19_), .CI(SUMB_15__20_), .CO(
        CARRYB_16__19_), .S(SUMB_16__19_) );
  FA_X1 S2_16_20 ( .A(ab_16__20_), .B(CARRYB_15__20_), .CI(SUMB_15__21_), .CO(
        CARRYB_16__20_), .S(SUMB_16__20_) );
  FA_X1 S2_16_21 ( .A(ab_16__21_), .B(CARRYB_15__21_), .CI(SUMB_15__22_), .CO(
        CARRYB_16__21_), .S(SUMB_16__21_) );
  FA_X1 S3_16_22 ( .A(ab_16__22_), .B(CARRYB_15__22_), .CI(ab_15__23_), .CO(
        CARRYB_16__22_), .S(SUMB_16__22_) );
  FA_X1 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  FA_X1 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  FA_X1 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  FA_X1 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  FA_X1 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  FA_X1 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  FA_X1 S2_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  FA_X1 S2_15_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), .CO(
        CARRYB_15__7_), .S(SUMB_15__7_) );
  FA_X1 S2_15_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), .CO(
        CARRYB_15__8_), .S(SUMB_15__8_) );
  FA_X1 S2_15_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), .CO(
        CARRYB_15__9_), .S(SUMB_15__9_) );
  FA_X1 S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), .CO(
        CARRYB_15__10_), .S(SUMB_15__10_) );
  FA_X1 S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), .CO(
        CARRYB_15__11_), .S(SUMB_15__11_) );
  FA_X1 S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), .CO(
        CARRYB_15__12_), .S(SUMB_15__12_) );
  FA_X1 S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), .CO(
        CARRYB_15__13_), .S(SUMB_15__13_) );
  FA_X1 S2_15_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), .CO(
        CARRYB_15__14_), .S(SUMB_15__14_) );
  FA_X1 S2_15_15 ( .A(ab_15__15_), .B(CARRYB_14__15_), .CI(SUMB_14__16_), .CO(
        CARRYB_15__15_), .S(SUMB_15__15_) );
  FA_X1 S2_15_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .CI(SUMB_14__17_), .CO(
        CARRYB_15__16_), .S(SUMB_15__16_) );
  FA_X1 S2_15_17 ( .A(ab_15__17_), .B(CARRYB_14__17_), .CI(SUMB_14__18_), .CO(
        CARRYB_15__17_), .S(SUMB_15__17_) );
  FA_X1 S2_15_18 ( .A(ab_15__18_), .B(CARRYB_14__18_), .CI(SUMB_14__19_), .CO(
        CARRYB_15__18_), .S(SUMB_15__18_) );
  FA_X1 S2_15_19 ( .A(ab_15__19_), .B(CARRYB_14__19_), .CI(SUMB_14__20_), .CO(
        CARRYB_15__19_), .S(SUMB_15__19_) );
  FA_X1 S2_15_20 ( .A(ab_15__20_), .B(CARRYB_14__20_), .CI(SUMB_14__21_), .CO(
        CARRYB_15__20_), .S(SUMB_15__20_) );
  FA_X1 S2_15_21 ( .A(ab_15__21_), .B(CARRYB_14__21_), .CI(SUMB_14__22_), .CO(
        CARRYB_15__21_), .S(SUMB_15__21_) );
  FA_X1 S3_15_22 ( .A(ab_15__22_), .B(CARRYB_14__22_), .CI(ab_14__23_), .CO(
        CARRYB_15__22_), .S(SUMB_15__22_) );
  FA_X1 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  FA_X1 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  FA_X1 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  FA_X1 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  FA_X1 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  FA_X1 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  FA_X1 S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  FA_X1 S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), .CO(
        CARRYB_14__7_), .S(SUMB_14__7_) );
  FA_X1 S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), .CO(
        CARRYB_14__8_), .S(SUMB_14__8_) );
  FA_X1 S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), .CO(
        CARRYB_14__9_), .S(SUMB_14__9_) );
  FA_X1 S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), .CO(
        CARRYB_14__10_), .S(SUMB_14__10_) );
  FA_X1 S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), .CO(
        CARRYB_14__11_), .S(SUMB_14__11_) );
  FA_X1 S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), .CO(
        CARRYB_14__12_), .S(SUMB_14__12_) );
  FA_X1 S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), .CO(
        CARRYB_14__13_), .S(SUMB_14__13_) );
  FA_X1 S2_14_14 ( .A(ab_14__14_), .B(CARRYB_13__14_), .CI(SUMB_13__15_), .CO(
        CARRYB_14__14_), .S(SUMB_14__14_) );
  FA_X1 S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), .CO(
        CARRYB_14__15_), .S(SUMB_14__15_) );
  FA_X1 S2_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), .CO(
        CARRYB_14__16_), .S(SUMB_14__16_) );
  FA_X1 S2_14_17 ( .A(ab_14__17_), .B(CARRYB_13__17_), .CI(SUMB_13__18_), .CO(
        CARRYB_14__17_), .S(SUMB_14__17_) );
  FA_X1 S2_14_18 ( .A(ab_14__18_), .B(CARRYB_13__18_), .CI(SUMB_13__19_), .CO(
        CARRYB_14__18_), .S(SUMB_14__18_) );
  FA_X1 S2_14_19 ( .A(ab_14__19_), .B(CARRYB_13__19_), .CI(SUMB_13__20_), .CO(
        CARRYB_14__19_), .S(SUMB_14__19_) );
  FA_X1 S2_14_20 ( .A(ab_14__20_), .B(CARRYB_13__20_), .CI(SUMB_13__21_), .CO(
        CARRYB_14__20_), .S(SUMB_14__20_) );
  FA_X1 S2_14_21 ( .A(ab_14__21_), .B(CARRYB_13__21_), .CI(SUMB_13__22_), .CO(
        CARRYB_14__21_), .S(SUMB_14__21_) );
  FA_X1 S3_14_22 ( .A(ab_14__22_), .B(CARRYB_13__22_), .CI(ab_13__23_), .CO(
        CARRYB_14__22_), .S(SUMB_14__22_) );
  FA_X1 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  FA_X1 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  FA_X1 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  FA_X1 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  FA_X1 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  FA_X1 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  FA_X1 S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  FA_X1 S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), .CO(
        CARRYB_13__7_), .S(SUMB_13__7_) );
  FA_X1 S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), .CO(
        CARRYB_13__8_), .S(SUMB_13__8_) );
  FA_X1 S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), .CO(
        CARRYB_13__9_), .S(SUMB_13__9_) );
  FA_X1 S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), .CO(
        CARRYB_13__10_), .S(SUMB_13__10_) );
  FA_X1 S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), .CO(
        CARRYB_13__11_), .S(SUMB_13__11_) );
  FA_X1 S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), .CO(
        CARRYB_13__12_), .S(SUMB_13__12_) );
  FA_X1 S2_13_13 ( .A(ab_13__13_), .B(CARRYB_12__13_), .CI(SUMB_12__14_), .CO(
        CARRYB_13__13_), .S(SUMB_13__13_) );
  FA_X1 S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), .CO(
        CARRYB_13__14_), .S(SUMB_13__14_) );
  FA_X1 S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), .CO(
        CARRYB_13__15_), .S(SUMB_13__15_) );
  FA_X1 S2_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), .CO(
        CARRYB_13__16_), .S(SUMB_13__16_) );
  FA_X1 S2_13_17 ( .A(ab_13__17_), .B(CARRYB_12__17_), .CI(SUMB_12__18_), .CO(
        CARRYB_13__17_), .S(SUMB_13__17_) );
  FA_X1 S2_13_18 ( .A(ab_13__18_), .B(CARRYB_12__18_), .CI(SUMB_12__19_), .CO(
        CARRYB_13__18_), .S(SUMB_13__18_) );
  FA_X1 S2_13_19 ( .A(ab_13__19_), .B(CARRYB_12__19_), .CI(SUMB_12__20_), .CO(
        CARRYB_13__19_), .S(SUMB_13__19_) );
  FA_X1 S2_13_20 ( .A(ab_13__20_), .B(CARRYB_12__20_), .CI(SUMB_12__21_), .CO(
        CARRYB_13__20_), .S(SUMB_13__20_) );
  FA_X1 S2_13_21 ( .A(ab_13__21_), .B(CARRYB_12__21_), .CI(SUMB_12__22_), .CO(
        CARRYB_13__21_), .S(SUMB_13__21_) );
  FA_X1 S3_13_22 ( .A(ab_13__22_), .B(CARRYB_12__22_), .CI(ab_12__23_), .CO(
        CARRYB_13__22_), .S(SUMB_13__22_) );
  FA_X1 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  FA_X1 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  FA_X1 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  FA_X1 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  FA_X1 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  FA_X1 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  FA_X1 S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  FA_X1 S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), .CO(
        CARRYB_12__7_), .S(SUMB_12__7_) );
  FA_X1 S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), .CO(
        CARRYB_12__8_), .S(SUMB_12__8_) );
  FA_X1 S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), .CO(
        CARRYB_12__9_), .S(SUMB_12__9_) );
  FA_X1 S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), .CO(
        CARRYB_12__10_), .S(SUMB_12__10_) );
  FA_X1 S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), .CO(
        CARRYB_12__11_), .S(SUMB_12__11_) );
  FA_X1 S2_12_12 ( .A(ab_12__12_), .B(CARRYB_11__12_), .CI(SUMB_11__13_), .CO(
        CARRYB_12__12_), .S(SUMB_12__12_) );
  FA_X1 S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), .CO(
        CARRYB_12__13_), .S(SUMB_12__13_) );
  FA_X1 S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), .CO(
        CARRYB_12__14_), .S(SUMB_12__14_) );
  FA_X1 S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), .CO(
        CARRYB_12__15_), .S(SUMB_12__15_) );
  FA_X1 S2_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), .CO(
        CARRYB_12__16_), .S(SUMB_12__16_) );
  FA_X1 S2_12_17 ( .A(ab_12__17_), .B(CARRYB_11__17_), .CI(SUMB_11__18_), .CO(
        CARRYB_12__17_), .S(SUMB_12__17_) );
  FA_X1 S2_12_18 ( .A(ab_12__18_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), .CO(
        CARRYB_12__18_), .S(SUMB_12__18_) );
  FA_X1 S2_12_19 ( .A(ab_12__19_), .B(CARRYB_11__19_), .CI(SUMB_11__20_), .CO(
        CARRYB_12__19_), .S(SUMB_12__19_) );
  FA_X1 S2_12_20 ( .A(ab_12__20_), .B(CARRYB_11__20_), .CI(SUMB_11__21_), .CO(
        CARRYB_12__20_), .S(SUMB_12__20_) );
  FA_X1 S2_12_21 ( .A(ab_12__21_), .B(CARRYB_11__21_), .CI(SUMB_11__22_), .CO(
        CARRYB_12__21_), .S(SUMB_12__21_) );
  FA_X1 S3_12_22 ( .A(ab_12__22_), .B(CARRYB_11__22_), .CI(ab_11__23_), .CO(
        CARRYB_12__22_), .S(SUMB_12__22_) );
  FA_X1 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  FA_X1 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  FA_X1 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  FA_X1 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  FA_X1 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  FA_X1 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  FA_X1 S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  FA_X1 S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), .CO(
        CARRYB_11__7_), .S(SUMB_11__7_) );
  FA_X1 S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), .CO(
        CARRYB_11__8_), .S(SUMB_11__8_) );
  FA_X1 S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), .CO(
        CARRYB_11__9_), .S(SUMB_11__9_) );
  FA_X1 S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), .CO(
        CARRYB_11__10_), .S(SUMB_11__10_) );
  FA_X1 S2_11_11 ( .A(ab_11__11_), .B(CARRYB_10__11_), .CI(SUMB_10__12_), .CO(
        CARRYB_11__11_), .S(SUMB_11__11_) );
  FA_X1 S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), .CO(
        CARRYB_11__12_), .S(SUMB_11__12_) );
  FA_X1 S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), .CO(
        CARRYB_11__13_), .S(SUMB_11__13_) );
  FA_X1 S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), .CO(
        CARRYB_11__14_), .S(SUMB_11__14_) );
  FA_X1 S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), .CO(
        CARRYB_11__15_), .S(SUMB_11__15_) );
  FA_X1 S2_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(SUMB_10__17_), .CO(
        CARRYB_11__16_), .S(SUMB_11__16_) );
  FA_X1 S2_11_17 ( .A(ab_11__17_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), .CO(
        CARRYB_11__17_), .S(SUMB_11__17_) );
  FA_X1 S2_11_18 ( .A(ab_11__18_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), .CO(
        CARRYB_11__18_), .S(SUMB_11__18_) );
  FA_X1 S2_11_19 ( .A(ab_11__19_), .B(CARRYB_10__19_), .CI(SUMB_10__20_), .CO(
        CARRYB_11__19_), .S(SUMB_11__19_) );
  FA_X1 S2_11_20 ( .A(ab_11__20_), .B(CARRYB_10__20_), .CI(SUMB_10__21_), .CO(
        CARRYB_11__20_), .S(SUMB_11__20_) );
  FA_X1 S2_11_21 ( .A(ab_11__21_), .B(CARRYB_10__21_), .CI(SUMB_10__22_), .CO(
        CARRYB_11__21_), .S(SUMB_11__21_) );
  FA_X1 S3_11_22 ( .A(ab_11__22_), .B(CARRYB_10__22_), .CI(ab_10__23_), .CO(
        CARRYB_11__22_), .S(SUMB_11__22_) );
  FA_X1 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  FA_X1 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  FA_X1 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  FA_X1 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  FA_X1 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  FA_X1 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  FA_X1 S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  FA_X1 S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  FA_X1 S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  FA_X1 S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  FA_X1 S2_10_10 ( .A(ab_10__10_), .B(CARRYB_9__10_), .CI(SUMB_9__11_), .CO(
        CARRYB_10__10_), .S(SUMB_10__10_) );
  FA_X1 S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), .CO(
        CARRYB_10__11_), .S(SUMB_10__11_) );
  FA_X1 S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), .CO(
        CARRYB_10__12_), .S(SUMB_10__12_) );
  FA_X1 S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), .CO(
        CARRYB_10__13_), .S(SUMB_10__13_) );
  FA_X1 S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), .CO(
        CARRYB_10__14_), .S(SUMB_10__14_) );
  FA_X1 S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), .CO(
        CARRYB_10__15_), .S(SUMB_10__15_) );
  FA_X1 S2_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), .CO(
        CARRYB_10__16_), .S(SUMB_10__16_) );
  FA_X1 S2_10_17 ( .A(ab_10__17_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), .CO(
        CARRYB_10__17_), .S(SUMB_10__17_) );
  FA_X1 S2_10_18 ( .A(ab_10__18_), .B(CARRYB_9__18_), .CI(SUMB_9__19_), .CO(
        CARRYB_10__18_), .S(SUMB_10__18_) );
  FA_X1 S2_10_19 ( .A(ab_10__19_), .B(CARRYB_9__19_), .CI(SUMB_9__20_), .CO(
        CARRYB_10__19_), .S(SUMB_10__19_) );
  FA_X1 S2_10_20 ( .A(ab_10__20_), .B(CARRYB_9__20_), .CI(SUMB_9__21_), .CO(
        CARRYB_10__20_), .S(SUMB_10__20_) );
  FA_X1 S2_10_21 ( .A(ab_10__21_), .B(CARRYB_9__21_), .CI(SUMB_9__22_), .CO(
        CARRYB_10__21_), .S(SUMB_10__21_) );
  FA_X1 S3_10_22 ( .A(ab_10__22_), .B(CARRYB_9__22_), .CI(ab_9__23_), .CO(
        CARRYB_10__22_), .S(SUMB_10__22_) );
  FA_X1 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  FA_X1 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  FA_X1 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  FA_X1 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  FA_X1 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  FA_X1 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  FA_X1 S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  FA_X1 S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  FA_X1 S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  FA_X1 S2_9_9 ( .A(ab_9__9_), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  FA_X1 S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), .CO(
        CARRYB_9__10_), .S(SUMB_9__10_) );
  FA_X1 S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), .CO(
        CARRYB_9__11_), .S(SUMB_9__11_) );
  FA_X1 S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), .CO(
        CARRYB_9__12_), .S(SUMB_9__12_) );
  FA_X1 S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), .CO(
        CARRYB_9__13_), .S(SUMB_9__13_) );
  FA_X1 S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), .CO(
        CARRYB_9__14_), .S(SUMB_9__14_) );
  FA_X1 S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), .CO(
        CARRYB_9__15_), .S(SUMB_9__15_) );
  FA_X1 S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), .CO(
        CARRYB_9__16_), .S(SUMB_9__16_) );
  FA_X1 S2_9_17 ( .A(ab_9__17_), .B(CARRYB_8__17_), .CI(SUMB_8__18_), .CO(
        CARRYB_9__17_), .S(SUMB_9__17_) );
  FA_X1 S2_9_18 ( .A(ab_9__18_), .B(CARRYB_8__18_), .CI(SUMB_8__19_), .CO(
        CARRYB_9__18_), .S(SUMB_9__18_) );
  FA_X1 S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), .CO(
        CARRYB_9__19_), .S(SUMB_9__19_) );
  FA_X1 S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(SUMB_8__21_), .CO(
        CARRYB_9__20_), .S(SUMB_9__20_) );
  FA_X1 S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), .CO(
        CARRYB_9__21_), .S(SUMB_9__21_) );
  FA_X1 S3_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .CI(ab_8__23_), .CO(
        CARRYB_9__22_), .S(SUMB_9__22_) );
  FA_X1 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  FA_X1 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  FA_X1 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  FA_X1 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  FA_X1 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  FA_X1 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  FA_X1 S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  FA_X1 S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  FA_X1 S2_8_8 ( .A(ab_8__8_), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  FA_X1 S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  FA_X1 S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), .CO(
        CARRYB_8__10_), .S(SUMB_8__10_) );
  FA_X1 S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), .CO(
        CARRYB_8__11_), .S(SUMB_8__11_) );
  FA_X1 S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), .CO(
        CARRYB_8__12_), .S(SUMB_8__12_) );
  FA_X1 S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), .CO(
        CARRYB_8__13_), .S(SUMB_8__13_) );
  FA_X1 S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), .CO(
        CARRYB_8__14_), .S(SUMB_8__14_) );
  FA_X1 S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), .CO(
        CARRYB_8__15_), .S(SUMB_8__15_) );
  FA_X1 S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), .CO(
        CARRYB_8__16_), .S(SUMB_8__16_) );
  FA_X1 S2_8_17 ( .A(ab_8__17_), .B(CARRYB_7__17_), .CI(SUMB_7__18_), .CO(
        CARRYB_8__17_), .S(SUMB_8__17_) );
  FA_X1 S2_8_18 ( .A(ab_8__18_), .B(CARRYB_7__18_), .CI(SUMB_7__19_), .CO(
        CARRYB_8__18_), .S(SUMB_8__18_) );
  FA_X1 S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), .CO(
        CARRYB_8__19_), .S(SUMB_8__19_) );
  FA_X1 S2_8_20 ( .A(ab_8__20_), .B(CARRYB_7__20_), .CI(SUMB_7__21_), .CO(
        CARRYB_8__20_), .S(SUMB_8__20_) );
  FA_X1 S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), .CO(
        CARRYB_8__21_), .S(SUMB_8__21_) );
  FA_X1 S3_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(ab_7__23_), .CO(
        CARRYB_8__22_), .S(SUMB_8__22_) );
  FA_X1 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(A1_5_) );
  FA_X1 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S2_7_7 ( .A(ab_7__7_), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  FA_X1 S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  FA_X1 S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  FA_X1 S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), .CO(
        CARRYB_7__10_), .S(SUMB_7__10_) );
  FA_X1 S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), .CO(
        CARRYB_7__11_), .S(SUMB_7__11_) );
  FA_X1 S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), .CO(
        CARRYB_7__12_), .S(SUMB_7__12_) );
  FA_X1 S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), .CO(
        CARRYB_7__13_), .S(SUMB_7__13_) );
  FA_X1 S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), .CO(
        CARRYB_7__14_), .S(SUMB_7__14_) );
  FA_X1 S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), .CO(
        CARRYB_7__15_), .S(SUMB_7__15_) );
  FA_X1 S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), .CO(
        CARRYB_7__16_), .S(SUMB_7__16_) );
  FA_X1 S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), .CO(
        CARRYB_7__17_), .S(SUMB_7__17_) );
  FA_X1 S2_7_18 ( .A(ab_7__18_), .B(CARRYB_6__18_), .CI(SUMB_6__19_), .CO(
        CARRYB_7__18_), .S(SUMB_7__18_) );
  FA_X1 S2_7_19 ( .A(ab_7__19_), .B(CARRYB_6__19_), .CI(SUMB_6__20_), .CO(
        CARRYB_7__19_), .S(SUMB_7__19_) );
  FA_X1 S2_7_20 ( .A(ab_7__20_), .B(CARRYB_6__20_), .CI(SUMB_6__21_), .CO(
        CARRYB_7__20_), .S(SUMB_7__20_) );
  FA_X1 S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), .CO(
        CARRYB_7__21_), .S(SUMB_7__21_) );
  FA_X1 S3_7_22 ( .A(ab_7__22_), .B(CARRYB_6__22_), .CI(ab_6__23_), .CO(
        CARRYB_7__22_), .S(SUMB_7__22_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S2_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  FA_X1 S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  FA_X1 S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  FA_X1 S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), .CO(
        CARRYB_6__10_), .S(SUMB_6__10_) );
  FA_X1 S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), .CO(
        CARRYB_6__11_), .S(SUMB_6__11_) );
  FA_X1 S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), .CO(
        CARRYB_6__12_), .S(SUMB_6__12_) );
  FA_X1 S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), .CO(
        CARRYB_6__13_), .S(SUMB_6__13_) );
  FA_X1 S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), .CO(
        CARRYB_6__14_), .S(SUMB_6__14_) );
  FA_X1 S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), .CO(
        CARRYB_6__15_), .S(SUMB_6__15_) );
  FA_X1 S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), .CO(
        CARRYB_6__16_), .S(SUMB_6__16_) );
  FA_X1 S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), .CO(
        CARRYB_6__17_), .S(SUMB_6__17_) );
  FA_X1 S2_6_18 ( .A(ab_6__18_), .B(CARRYB_5__18_), .CI(SUMB_5__19_), .CO(
        CARRYB_6__18_), .S(SUMB_6__18_) );
  FA_X1 S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), .CO(
        CARRYB_6__19_), .S(SUMB_6__19_) );
  FA_X1 S2_6_20 ( .A(ab_6__20_), .B(CARRYB_5__20_), .CI(SUMB_5__21_), .CO(
        CARRYB_6__20_), .S(SUMB_6__20_) );
  FA_X1 S2_6_21 ( .A(ab_6__21_), .B(CARRYB_5__21_), .CI(SUMB_5__22_), .CO(
        CARRYB_6__21_), .S(SUMB_6__21_) );
  FA_X1 S3_6_22 ( .A(ab_6__22_), .B(CARRYB_5__22_), .CI(ab_5__23_), .CO(
        CARRYB_6__22_), .S(SUMB_6__22_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  FA_X1 S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  FA_X1 S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  FA_X1 S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), .CO(
        CARRYB_5__10_), .S(SUMB_5__10_) );
  FA_X1 S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), .CO(
        CARRYB_5__11_), .S(SUMB_5__11_) );
  FA_X1 S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), .CO(
        CARRYB_5__12_), .S(SUMB_5__12_) );
  FA_X1 S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), .CO(
        CARRYB_5__13_), .S(SUMB_5__13_) );
  FA_X1 S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), .CO(
        CARRYB_5__14_), .S(SUMB_5__14_) );
  FA_X1 S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), .CO(
        CARRYB_5__15_), .S(SUMB_5__15_) );
  FA_X1 S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), .CO(
        CARRYB_5__16_), .S(SUMB_5__16_) );
  FA_X1 S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), .CO(
        CARRYB_5__17_), .S(SUMB_5__17_) );
  FA_X1 S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), .CO(
        CARRYB_5__18_), .S(SUMB_5__18_) );
  FA_X1 S2_5_19 ( .A(ab_5__19_), .B(CARRYB_4__19_), .CI(SUMB_4__20_), .CO(
        CARRYB_5__19_), .S(SUMB_5__19_) );
  FA_X1 S2_5_20 ( .A(ab_5__20_), .B(CARRYB_4__20_), .CI(SUMB_4__21_), .CO(
        CARRYB_5__20_), .S(SUMB_5__20_) );
  FA_X1 S2_5_21 ( .A(ab_5__21_), .B(CARRYB_4__21_), .CI(SUMB_4__22_), .CO(
        CARRYB_5__21_), .S(SUMB_5__21_) );
  FA_X1 S3_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(ab_4__23_), .CO(
        CARRYB_5__22_), .S(SUMB_5__22_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  FA_X1 S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  FA_X1 S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  FA_X1 S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), .CO(
        CARRYB_4__10_), .S(SUMB_4__10_) );
  FA_X1 S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), .CO(
        CARRYB_4__11_), .S(SUMB_4__11_) );
  FA_X1 S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), .CO(
        CARRYB_4__12_), .S(SUMB_4__12_) );
  FA_X1 S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), .CO(
        CARRYB_4__13_), .S(SUMB_4__13_) );
  FA_X1 S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), .CO(
        CARRYB_4__14_), .S(SUMB_4__14_) );
  FA_X1 S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), .CO(
        CARRYB_4__15_), .S(SUMB_4__15_) );
  FA_X1 S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), .CO(
        CARRYB_4__16_), .S(SUMB_4__16_) );
  FA_X1 S2_4_17 ( .A(ab_4__17_), .B(CARRYB_3__17_), .CI(SUMB_3__18_), .CO(
        CARRYB_4__17_), .S(SUMB_4__17_) );
  FA_X1 S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), .CO(
        CARRYB_4__18_), .S(SUMB_4__18_) );
  FA_X1 S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), .CO(
        CARRYB_4__19_), .S(SUMB_4__19_) );
  FA_X1 S2_4_20 ( .A(ab_4__20_), .B(CARRYB_3__20_), .CI(SUMB_3__21_), .CO(
        CARRYB_4__20_), .S(SUMB_4__20_) );
  FA_X1 S2_4_21 ( .A(ab_4__21_), .B(CARRYB_3__21_), .CI(SUMB_3__22_), .CO(
        CARRYB_4__21_), .S(SUMB_4__21_) );
  FA_X1 S3_4_22 ( .A(ab_4__22_), .B(CARRYB_3__22_), .CI(ab_3__23_), .CO(
        CARRYB_4__22_), .S(SUMB_4__22_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  FA_X1 S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  FA_X1 S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  FA_X1 S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), .CO(
        CARRYB_3__10_), .S(SUMB_3__10_) );
  FA_X1 S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), .CO(
        CARRYB_3__11_), .S(SUMB_3__11_) );
  FA_X1 S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), .CO(
        CARRYB_3__12_), .S(SUMB_3__12_) );
  FA_X1 S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), .CO(
        CARRYB_3__13_), .S(SUMB_3__13_) );
  FA_X1 S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), .CO(
        CARRYB_3__14_), .S(SUMB_3__14_) );
  FA_X1 S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), .CO(
        CARRYB_3__15_), .S(SUMB_3__15_) );
  FA_X1 S2_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(SUMB_2__17_), .CO(
        CARRYB_3__16_), .S(SUMB_3__16_) );
  FA_X1 S2_3_17 ( .A(ab_3__17_), .B(CARRYB_2__17_), .CI(SUMB_2__18_), .CO(
        CARRYB_3__17_), .S(SUMB_3__17_) );
  FA_X1 S2_3_18 ( .A(ab_3__18_), .B(CARRYB_2__18_), .CI(SUMB_2__19_), .CO(
        CARRYB_3__18_), .S(SUMB_3__18_) );
  FA_X1 S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), .CO(
        CARRYB_3__19_), .S(SUMB_3__19_) );
  FA_X1 S2_3_20 ( .A(ab_3__20_), .B(CARRYB_2__20_), .CI(SUMB_2__21_), .CO(
        CARRYB_3__20_), .S(SUMB_3__20_) );
  FA_X1 S2_3_21 ( .A(ab_3__21_), .B(CARRYB_2__21_), .CI(SUMB_2__22_), .CO(
        CARRYB_3__21_), .S(SUMB_3__21_) );
  FA_X1 S3_3_22 ( .A(ab_3__22_), .B(CARRYB_2__22_), .CI(ab_2__23_), .CO(
        CARRYB_3__22_), .S(SUMB_3__22_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S2_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(SUMB_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  FA_X1 S2_2_7 ( .A(ab_2__7_), .B(CARRYB_1__7_), .CI(SUMB_1__8_), .CO(
        CARRYB_2__7_), .S(SUMB_2__7_) );
  FA_X1 S2_2_8 ( .A(ab_2__8_), .B(CARRYB_1__8_), .CI(SUMB_1__9_), .CO(
        CARRYB_2__8_), .S(SUMB_2__8_) );
  FA_X1 S2_2_9 ( .A(ab_2__9_), .B(CARRYB_1__9_), .CI(SUMB_1__10_), .CO(
        CARRYB_2__9_), .S(SUMB_2__9_) );
  FA_X1 S2_2_10 ( .A(ab_2__10_), .B(CARRYB_1__10_), .CI(SUMB_1__11_), .CO(
        CARRYB_2__10_), .S(SUMB_2__10_) );
  FA_X1 S2_2_11 ( .A(ab_2__11_), .B(CARRYB_1__11_), .CI(SUMB_1__12_), .CO(
        CARRYB_2__11_), .S(SUMB_2__11_) );
  FA_X1 S2_2_12 ( .A(ab_2__12_), .B(CARRYB_1__12_), .CI(SUMB_1__13_), .CO(
        CARRYB_2__12_), .S(SUMB_2__12_) );
  FA_X1 S2_2_13 ( .A(ab_2__13_), .B(CARRYB_1__13_), .CI(SUMB_1__14_), .CO(
        CARRYB_2__13_), .S(SUMB_2__13_) );
  FA_X1 S2_2_14 ( .A(ab_2__14_), .B(CARRYB_1__14_), .CI(SUMB_1__15_), .CO(
        CARRYB_2__14_), .S(SUMB_2__14_) );
  FA_X1 S2_2_15 ( .A(ab_2__15_), .B(CARRYB_1__15_), .CI(SUMB_1__16_), .CO(
        CARRYB_2__15_), .S(SUMB_2__15_) );
  FA_X1 S2_2_16 ( .A(ab_2__16_), .B(CARRYB_1__16_), .CI(SUMB_1__17_), .CO(
        CARRYB_2__16_), .S(SUMB_2__16_) );
  FA_X1 S2_2_17 ( .A(ab_2__17_), .B(CARRYB_1__17_), .CI(SUMB_1__18_), .CO(
        CARRYB_2__17_), .S(SUMB_2__17_) );
  FA_X1 S2_2_18 ( .A(ab_2__18_), .B(CARRYB_1__18_), .CI(SUMB_1__19_), .CO(
        CARRYB_2__18_), .S(SUMB_2__18_) );
  FA_X1 S2_2_19 ( .A(ab_2__19_), .B(CARRYB_1__19_), .CI(SUMB_1__20_), .CO(
        CARRYB_2__19_), .S(SUMB_2__19_) );
  FA_X1 S2_2_20 ( .A(ab_2__20_), .B(CARRYB_1__20_), .CI(SUMB_1__21_), .CO(
        CARRYB_2__20_), .S(SUMB_2__20_) );
  FA_X1 S2_2_21 ( .A(ab_2__21_), .B(CARRYB_1__21_), .CI(SUMB_1__22_), .CO(
        CARRYB_2__21_), .S(SUMB_2__21_) );
  FA_X1 S3_2_22 ( .A(ab_2__22_), .B(CARRYB_1__22_), .CI(ab_1__23_), .CO(
        CARRYB_2__22_), .S(SUMB_2__22_) );
  iir_filter_DW01_add_7 FS_1 ( .A({A1_45_, A1_44_, A1_43_, A1_42_, A1_41_, 
        A1_40_, A1_39_, A1_38_, A1_37_, A1_36_, A1_35_, A1_34_, A1_33_, A1_32_, 
        A1_31_, A1_30_, A1_29_, A1_28_, A1_27_, A1_26_, A1_25_, A1_24_, A1_23_, 
        A1_22_, A1_21_, A1_20_, A1_19_, A1_18_, A1_17_, A1_16_, A1_15_, A1_14_, 
        A1_13_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, A1_5_, 
        A1_4_, A1_3_, A1_2_, A1_1_, A1_0_}), .B({A2_45_, A2_44_, A2_43_, 
        A2_42_, A2_41_, A2_40_, A2_39_, A2_38_, A2_37_, A2_36_, A2_35_, A2_34_, 
        A2_33_, A2_32_, A2_31_, A2_30_, A2_29_, A2_28_, A2_27_, A2_26_, A2_25_, 
        A2_24_, A2_23_, A2_22_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({PRODUCT[47], SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, PRODUCT[44:22], SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21}) );
  BUF_X1 U2 ( .A(QB), .Z(n1) );
  BUF_X1 U3 ( .A(QB), .Z(n2) );
  BUF_X1 U4 ( .A(QA), .Z(n3) );
  BUF_X1 U5 ( .A(QA), .Z(n4) );
  INV_X1 U6 ( .A(A[2]), .ZN(n36) );
  INV_X1 U7 ( .A(A[3]), .ZN(n35) );
  INV_X1 U8 ( .A(A[4]), .ZN(n34) );
  INV_X1 U9 ( .A(A[5]), .ZN(n33) );
  INV_X1 U10 ( .A(A[6]), .ZN(n32) );
  INV_X1 U11 ( .A(B[1]), .ZN(n18) );
  INV_X1 U12 ( .A(A[1]), .ZN(n40) );
  INV_X1 U13 ( .A(B[0]), .ZN(n29) );
  INV_X1 U14 ( .A(A[0]), .ZN(n51) );
  INV_X1 U15 ( .A(B[22]), .ZN(n15) );
  INV_X1 U16 ( .A(B[21]), .ZN(n16) );
  INV_X1 U17 ( .A(B[20]), .ZN(n17) );
  INV_X1 U18 ( .A(B[19]), .ZN(n19) );
  INV_X1 U19 ( .A(B[18]), .ZN(n20) );
  INV_X1 U20 ( .A(B[17]), .ZN(n21) );
  INV_X1 U21 ( .A(B[16]), .ZN(n22) );
  INV_X1 U22 ( .A(B[15]), .ZN(n23) );
  INV_X1 U23 ( .A(B[14]), .ZN(n24) );
  INV_X1 U24 ( .A(B[13]), .ZN(n25) );
  INV_X1 U25 ( .A(B[12]), .ZN(n26) );
  INV_X1 U26 ( .A(B[11]), .ZN(n27) );
  INV_X1 U27 ( .A(B[10]), .ZN(n28) );
  INV_X1 U28 ( .A(B[9]), .ZN(n7) );
  INV_X1 U29 ( .A(B[8]), .ZN(n8) );
  INV_X1 U30 ( .A(B[7]), .ZN(n9) );
  INV_X1 U31 ( .A(B[6]), .ZN(n10) );
  INV_X1 U32 ( .A(B[5]), .ZN(n11) );
  INV_X1 U33 ( .A(B[4]), .ZN(n12) );
  INV_X1 U34 ( .A(B[3]), .ZN(n13) );
  INV_X1 U35 ( .A(B[2]), .ZN(n14) );
  INV_X1 U36 ( .A(A[7]), .ZN(n31) );
  INV_X1 U37 ( .A(A[8]), .ZN(n30) );
  INV_X1 U38 ( .A(A[10]), .ZN(n50) );
  INV_X1 U39 ( .A(A[11]), .ZN(n49) );
  INV_X1 U40 ( .A(A[12]), .ZN(n48) );
  INV_X1 U41 ( .A(A[13]), .ZN(n47) );
  INV_X1 U42 ( .A(A[14]), .ZN(n46) );
  INV_X1 U43 ( .A(A[9]), .ZN(n6) );
  INV_X1 U44 ( .A(A[22]), .ZN(n37) );
  INV_X1 U45 ( .A(A[15]), .ZN(n45) );
  INV_X1 U46 ( .A(A[16]), .ZN(n44) );
  INV_X1 U47 ( .A(A[17]), .ZN(n43) );
  INV_X1 U48 ( .A(A[18]), .ZN(n42) );
  INV_X1 U49 ( .A(A[19]), .ZN(n41) );
  INV_X1 U50 ( .A(A[20]), .ZN(n39) );
  INV_X1 U51 ( .A(A[21]), .ZN(n38) );
  AND2_X1 U52 ( .A1(SUMB_23__23_), .A2(CARRYB_23__22_), .ZN(A2_45_) );
  XOR2_X1 U53 ( .A(CARRYB_23__22_), .B(SUMB_23__23_), .Z(A1_44_) );
  AND2_X1 U54 ( .A1(SUMB_23__22_), .A2(CARRYB_23__21_), .ZN(A2_44_) );
  XOR2_X1 U55 ( .A(CARRYB_23__21_), .B(SUMB_23__22_), .Z(A1_43_) );
  AND2_X1 U56 ( .A1(SUMB_23__21_), .A2(CARRYB_23__20_), .ZN(A2_43_) );
  XOR2_X1 U57 ( .A(CARRYB_23__20_), .B(SUMB_23__21_), .Z(A1_42_) );
  AND2_X1 U58 ( .A1(SUMB_23__20_), .A2(CARRYB_23__19_), .ZN(A2_42_) );
  XOR2_X1 U59 ( .A(CARRYB_23__19_), .B(SUMB_23__20_), .Z(A1_41_) );
  AND2_X1 U60 ( .A1(SUMB_23__19_), .A2(CARRYB_23__18_), .ZN(A2_41_) );
  XOR2_X1 U61 ( .A(CARRYB_23__18_), .B(SUMB_23__19_), .Z(A1_40_) );
  AND2_X1 U62 ( .A1(SUMB_23__18_), .A2(CARRYB_23__17_), .ZN(A2_40_) );
  XOR2_X1 U63 ( .A(CARRYB_23__17_), .B(SUMB_23__18_), .Z(A1_39_) );
  AND2_X1 U64 ( .A1(SUMB_23__17_), .A2(CARRYB_23__16_), .ZN(A2_39_) );
  XOR2_X1 U65 ( .A(CARRYB_23__16_), .B(SUMB_23__17_), .Z(A1_38_) );
  AND2_X1 U66 ( .A1(SUMB_23__16_), .A2(CARRYB_23__15_), .ZN(A2_38_) );
  XOR2_X1 U67 ( .A(CARRYB_23__15_), .B(SUMB_23__16_), .Z(A1_37_) );
  AND2_X1 U68 ( .A1(SUMB_23__15_), .A2(CARRYB_23__14_), .ZN(A2_37_) );
  XOR2_X1 U69 ( .A(CARRYB_23__14_), .B(SUMB_23__15_), .Z(A1_36_) );
  AND2_X1 U70 ( .A1(SUMB_23__14_), .A2(CARRYB_23__13_), .ZN(A2_36_) );
  XOR2_X1 U71 ( .A(CARRYB_23__13_), .B(SUMB_23__14_), .Z(A1_35_) );
  AND2_X1 U72 ( .A1(SUMB_23__13_), .A2(CARRYB_23__12_), .ZN(A2_35_) );
  XOR2_X1 U73 ( .A(CARRYB_23__12_), .B(SUMB_23__13_), .Z(A1_34_) );
  AND2_X1 U74 ( .A1(SUMB_23__12_), .A2(CARRYB_23__11_), .ZN(A2_34_) );
  XOR2_X1 U75 ( .A(CARRYB_23__11_), .B(SUMB_23__12_), .Z(A1_33_) );
  AND2_X1 U76 ( .A1(SUMB_23__11_), .A2(CARRYB_23__10_), .ZN(A2_33_) );
  XOR2_X1 U77 ( .A(CARRYB_23__10_), .B(SUMB_23__11_), .Z(A1_32_) );
  AND2_X1 U78 ( .A1(SUMB_23__10_), .A2(CARRYB_23__9_), .ZN(A2_32_) );
  XOR2_X1 U79 ( .A(CARRYB_23__9_), .B(SUMB_23__10_), .Z(A1_31_) );
  AND2_X1 U80 ( .A1(SUMB_23__9_), .A2(CARRYB_23__8_), .ZN(A2_31_) );
  XOR2_X1 U81 ( .A(CARRYB_23__8_), .B(SUMB_23__9_), .Z(A1_30_) );
  AND2_X1 U82 ( .A1(SUMB_23__8_), .A2(CARRYB_23__7_), .ZN(A2_30_) );
  XOR2_X1 U83 ( .A(CARRYB_23__7_), .B(SUMB_23__8_), .Z(A1_29_) );
  AND2_X1 U84 ( .A1(SUMB_23__7_), .A2(CARRYB_23__6_), .ZN(A2_29_) );
  XOR2_X1 U85 ( .A(CARRYB_23__6_), .B(SUMB_23__7_), .Z(A1_28_) );
  AND2_X1 U86 ( .A1(SUMB_23__6_), .A2(CARRYB_23__5_), .ZN(A2_28_) );
  XOR2_X1 U87 ( .A(CARRYB_23__5_), .B(SUMB_23__6_), .Z(A1_27_) );
  AND2_X1 U88 ( .A1(SUMB_23__5_), .A2(CARRYB_23__4_), .ZN(A2_27_) );
  XOR2_X1 U89 ( .A(CARRYB_23__4_), .B(SUMB_23__5_), .Z(A1_26_) );
  AND2_X1 U90 ( .A1(SUMB_23__4_), .A2(CARRYB_23__3_), .ZN(A2_26_) );
  XOR2_X1 U91 ( .A(CARRYB_23__3_), .B(SUMB_23__4_), .Z(A1_25_) );
  AND2_X1 U92 ( .A1(SUMB_23__3_), .A2(CARRYB_23__2_), .ZN(A2_25_) );
  XOR2_X1 U93 ( .A(CARRYB_23__2_), .B(SUMB_23__3_), .Z(A1_24_) );
  AND2_X1 U94 ( .A1(SUMB_23__2_), .A2(CARRYB_23__1_), .ZN(A2_24_) );
  XOR2_X1 U95 ( .A(CARRYB_23__1_), .B(SUMB_23__2_), .Z(A1_23_) );
  AND2_X1 U96 ( .A1(SUMB_23__1_), .A2(CARRYB_23__0_), .ZN(A2_23_) );
  XOR2_X1 U97 ( .A(CARRYB_23__0_), .B(SUMB_23__1_), .Z(A1_22_) );
  AND2_X1 U98 ( .A1(ab_1__22_), .A2(ab_0__23_), .ZN(CARRYB_1__22_) );
  XOR2_X1 U99 ( .A(ab_1__22_), .B(ab_0__23_), .Z(SUMB_1__22_) );
  AND2_X1 U100 ( .A1(ab_1__21_), .A2(ab_0__22_), .ZN(CARRYB_1__21_) );
  XOR2_X1 U101 ( .A(ab_1__21_), .B(ab_0__22_), .Z(SUMB_1__21_) );
  AND2_X1 U102 ( .A1(ab_1__20_), .A2(ab_0__21_), .ZN(CARRYB_1__20_) );
  XOR2_X1 U103 ( .A(ab_1__20_), .B(ab_0__21_), .Z(SUMB_1__20_) );
  AND2_X1 U104 ( .A1(ab_1__19_), .A2(ab_0__20_), .ZN(CARRYB_1__19_) );
  XOR2_X1 U105 ( .A(ab_1__19_), .B(ab_0__20_), .Z(SUMB_1__19_) );
  AND2_X1 U106 ( .A1(ab_1__18_), .A2(ab_0__19_), .ZN(CARRYB_1__18_) );
  XOR2_X1 U107 ( .A(ab_1__18_), .B(ab_0__19_), .Z(SUMB_1__18_) );
  AND2_X1 U108 ( .A1(ab_1__17_), .A2(ab_0__18_), .ZN(CARRYB_1__17_) );
  XOR2_X1 U109 ( .A(ab_1__17_), .B(ab_0__18_), .Z(SUMB_1__17_) );
  AND2_X1 U110 ( .A1(ab_1__16_), .A2(ab_0__17_), .ZN(CARRYB_1__16_) );
  XOR2_X1 U111 ( .A(ab_1__16_), .B(ab_0__17_), .Z(SUMB_1__16_) );
  AND2_X1 U112 ( .A1(ab_1__15_), .A2(ab_0__16_), .ZN(CARRYB_1__15_) );
  XOR2_X1 U113 ( .A(ab_1__15_), .B(ab_0__16_), .Z(SUMB_1__15_) );
  AND2_X1 U114 ( .A1(ab_1__14_), .A2(ab_0__15_), .ZN(CARRYB_1__14_) );
  XOR2_X1 U115 ( .A(ab_1__14_), .B(ab_0__15_), .Z(SUMB_1__14_) );
  AND2_X1 U116 ( .A1(ab_1__13_), .A2(ab_0__14_), .ZN(CARRYB_1__13_) );
  XOR2_X1 U117 ( .A(ab_1__13_), .B(ab_0__14_), .Z(SUMB_1__13_) );
  AND2_X1 U118 ( .A1(ab_1__12_), .A2(ab_0__13_), .ZN(CARRYB_1__12_) );
  XOR2_X1 U119 ( .A(ab_1__12_), .B(ab_0__13_), .Z(SUMB_1__12_) );
  AND2_X1 U120 ( .A1(ab_1__11_), .A2(ab_0__12_), .ZN(CARRYB_1__11_) );
  XOR2_X1 U121 ( .A(ab_1__11_), .B(ab_0__12_), .Z(SUMB_1__11_) );
  AND2_X1 U122 ( .A1(ab_1__10_), .A2(ab_0__11_), .ZN(CARRYB_1__10_) );
  XOR2_X1 U123 ( .A(ab_1__10_), .B(ab_0__11_), .Z(SUMB_1__10_) );
  AND2_X1 U124 ( .A1(ab_1__9_), .A2(ab_0__10_), .ZN(CARRYB_1__9_) );
  XOR2_X1 U125 ( .A(ab_1__9_), .B(ab_0__10_), .Z(SUMB_1__9_) );
  AND2_X1 U126 ( .A1(ab_1__8_), .A2(ab_0__9_), .ZN(CARRYB_1__8_) );
  XOR2_X1 U127 ( .A(ab_1__8_), .B(ab_0__9_), .Z(SUMB_1__8_) );
  AND2_X1 U128 ( .A1(ab_1__7_), .A2(ab_0__8_), .ZN(CARRYB_1__7_) );
  XOR2_X1 U129 ( .A(ab_1__7_), .B(ab_0__8_), .Z(SUMB_1__7_) );
  AND2_X1 U130 ( .A1(ab_1__6_), .A2(ab_0__7_), .ZN(CARRYB_1__6_) );
  XOR2_X1 U131 ( .A(ab_1__6_), .B(ab_0__7_), .Z(SUMB_1__6_) );
  AND2_X1 U132 ( .A1(ab_1__5_), .A2(ab_0__6_), .ZN(CARRYB_1__5_) );
  XOR2_X1 U133 ( .A(ab_1__5_), .B(ab_0__6_), .Z(SUMB_1__5_) );
  AND2_X1 U134 ( .A1(ab_1__4_), .A2(ab_0__5_), .ZN(CARRYB_1__4_) );
  XOR2_X1 U135 ( .A(ab_1__4_), .B(ab_0__5_), .Z(SUMB_1__4_) );
  AND2_X1 U136 ( .A1(ab_1__3_), .A2(ab_0__4_), .ZN(CARRYB_1__3_) );
  XOR2_X1 U137 ( .A(ab_1__3_), .B(ab_0__4_), .Z(SUMB_1__3_) );
  AND2_X1 U138 ( .A1(ab_1__2_), .A2(ab_0__3_), .ZN(CARRYB_1__2_) );
  XOR2_X1 U139 ( .A(ab_1__2_), .B(ab_0__3_), .Z(SUMB_1__2_) );
  AND2_X1 U140 ( .A1(ab_1__1_), .A2(ab_0__2_), .ZN(CARRYB_1__1_) );
  XOR2_X1 U141 ( .A(ab_1__1_), .B(ab_0__2_), .Z(SUMB_1__1_) );
  NOR2_X1 U142 ( .A1(n6), .A2(n7), .ZN(ab_9__9_) );
  NOR2_X1 U143 ( .A1(n6), .A2(n8), .ZN(ab_9__8_) );
  NOR2_X1 U144 ( .A1(n6), .A2(n9), .ZN(ab_9__7_) );
  NOR2_X1 U145 ( .A1(n6), .A2(n10), .ZN(ab_9__6_) );
  NOR2_X1 U146 ( .A1(n6), .A2(n11), .ZN(ab_9__5_) );
  NOR2_X1 U147 ( .A1(n6), .A2(n12), .ZN(ab_9__4_) );
  NOR2_X1 U148 ( .A1(n6), .A2(n13), .ZN(ab_9__3_) );
  NOR2_X1 U149 ( .A1(n6), .A2(n14), .ZN(ab_9__2_) );
  NOR2_X1 U150 ( .A1(A[9]), .A2(n1), .ZN(ab_9__23_) );
  NOR2_X1 U151 ( .A1(n6), .A2(n15), .ZN(ab_9__22_) );
  NOR2_X1 U152 ( .A1(n6), .A2(n16), .ZN(ab_9__21_) );
  NOR2_X1 U153 ( .A1(n6), .A2(n17), .ZN(ab_9__20_) );
  NOR2_X1 U154 ( .A1(n6), .A2(n18), .ZN(ab_9__1_) );
  NOR2_X1 U155 ( .A1(n6), .A2(n19), .ZN(ab_9__19_) );
  NOR2_X1 U156 ( .A1(n6), .A2(n20), .ZN(ab_9__18_) );
  NOR2_X1 U157 ( .A1(n6), .A2(n21), .ZN(ab_9__17_) );
  NOR2_X1 U158 ( .A1(n6), .A2(n22), .ZN(ab_9__16_) );
  NOR2_X1 U159 ( .A1(n6), .A2(n23), .ZN(ab_9__15_) );
  NOR2_X1 U160 ( .A1(n6), .A2(n24), .ZN(ab_9__14_) );
  NOR2_X1 U161 ( .A1(n6), .A2(n25), .ZN(ab_9__13_) );
  NOR2_X1 U162 ( .A1(n6), .A2(n26), .ZN(ab_9__12_) );
  NOR2_X1 U163 ( .A1(n6), .A2(n27), .ZN(ab_9__11_) );
  NOR2_X1 U164 ( .A1(n6), .A2(n28), .ZN(ab_9__10_) );
  NOR2_X1 U165 ( .A1(n6), .A2(n29), .ZN(ab_9__0_) );
  NOR2_X1 U166 ( .A1(n7), .A2(n30), .ZN(ab_8__9_) );
  NOR2_X1 U167 ( .A1(n8), .A2(n30), .ZN(ab_8__8_) );
  NOR2_X1 U168 ( .A1(n9), .A2(n30), .ZN(ab_8__7_) );
  NOR2_X1 U169 ( .A1(n10), .A2(n30), .ZN(ab_8__6_) );
  NOR2_X1 U170 ( .A1(n11), .A2(n30), .ZN(ab_8__5_) );
  NOR2_X1 U171 ( .A1(n12), .A2(n30), .ZN(ab_8__4_) );
  NOR2_X1 U172 ( .A1(n13), .A2(n30), .ZN(ab_8__3_) );
  NOR2_X1 U173 ( .A1(n14), .A2(n30), .ZN(ab_8__2_) );
  NOR2_X1 U174 ( .A1(A[8]), .A2(n1), .ZN(ab_8__23_) );
  NOR2_X1 U175 ( .A1(n15), .A2(n30), .ZN(ab_8__22_) );
  NOR2_X1 U176 ( .A1(n16), .A2(n30), .ZN(ab_8__21_) );
  NOR2_X1 U177 ( .A1(n17), .A2(n30), .ZN(ab_8__20_) );
  NOR2_X1 U178 ( .A1(n18), .A2(n30), .ZN(ab_8__1_) );
  NOR2_X1 U179 ( .A1(n19), .A2(n30), .ZN(ab_8__19_) );
  NOR2_X1 U180 ( .A1(n20), .A2(n30), .ZN(ab_8__18_) );
  NOR2_X1 U181 ( .A1(n21), .A2(n30), .ZN(ab_8__17_) );
  NOR2_X1 U182 ( .A1(n22), .A2(n30), .ZN(ab_8__16_) );
  NOR2_X1 U183 ( .A1(n23), .A2(n30), .ZN(ab_8__15_) );
  NOR2_X1 U184 ( .A1(n24), .A2(n30), .ZN(ab_8__14_) );
  NOR2_X1 U185 ( .A1(n25), .A2(n30), .ZN(ab_8__13_) );
  NOR2_X1 U186 ( .A1(n26), .A2(n30), .ZN(ab_8__12_) );
  NOR2_X1 U187 ( .A1(n27), .A2(n30), .ZN(ab_8__11_) );
  NOR2_X1 U188 ( .A1(n28), .A2(n30), .ZN(ab_8__10_) );
  NOR2_X1 U189 ( .A1(n29), .A2(n30), .ZN(ab_8__0_) );
  NOR2_X1 U190 ( .A1(n7), .A2(n31), .ZN(ab_7__9_) );
  NOR2_X1 U191 ( .A1(n8), .A2(n31), .ZN(ab_7__8_) );
  NOR2_X1 U192 ( .A1(n9), .A2(n31), .ZN(ab_7__7_) );
  NOR2_X1 U193 ( .A1(n10), .A2(n31), .ZN(ab_7__6_) );
  NOR2_X1 U194 ( .A1(n11), .A2(n31), .ZN(ab_7__5_) );
  NOR2_X1 U195 ( .A1(n12), .A2(n31), .ZN(ab_7__4_) );
  NOR2_X1 U196 ( .A1(n13), .A2(n31), .ZN(ab_7__3_) );
  NOR2_X1 U197 ( .A1(n14), .A2(n31), .ZN(ab_7__2_) );
  NOR2_X1 U198 ( .A1(A[7]), .A2(n1), .ZN(ab_7__23_) );
  NOR2_X1 U199 ( .A1(n15), .A2(n31), .ZN(ab_7__22_) );
  NOR2_X1 U200 ( .A1(n16), .A2(n31), .ZN(ab_7__21_) );
  NOR2_X1 U201 ( .A1(n17), .A2(n31), .ZN(ab_7__20_) );
  NOR2_X1 U202 ( .A1(n18), .A2(n31), .ZN(ab_7__1_) );
  NOR2_X1 U203 ( .A1(n19), .A2(n31), .ZN(ab_7__19_) );
  NOR2_X1 U204 ( .A1(n20), .A2(n31), .ZN(ab_7__18_) );
  NOR2_X1 U205 ( .A1(n21), .A2(n31), .ZN(ab_7__17_) );
  NOR2_X1 U206 ( .A1(n22), .A2(n31), .ZN(ab_7__16_) );
  NOR2_X1 U207 ( .A1(n23), .A2(n31), .ZN(ab_7__15_) );
  NOR2_X1 U208 ( .A1(n24), .A2(n31), .ZN(ab_7__14_) );
  NOR2_X1 U209 ( .A1(n25), .A2(n31), .ZN(ab_7__13_) );
  NOR2_X1 U210 ( .A1(n26), .A2(n31), .ZN(ab_7__12_) );
  NOR2_X1 U211 ( .A1(n27), .A2(n31), .ZN(ab_7__11_) );
  NOR2_X1 U212 ( .A1(n28), .A2(n31), .ZN(ab_7__10_) );
  NOR2_X1 U213 ( .A1(n29), .A2(n31), .ZN(ab_7__0_) );
  NOR2_X1 U214 ( .A1(n7), .A2(n32), .ZN(ab_6__9_) );
  NOR2_X1 U215 ( .A1(n8), .A2(n32), .ZN(ab_6__8_) );
  NOR2_X1 U216 ( .A1(n9), .A2(n32), .ZN(ab_6__7_) );
  NOR2_X1 U217 ( .A1(n10), .A2(n32), .ZN(ab_6__6_) );
  NOR2_X1 U218 ( .A1(n11), .A2(n32), .ZN(ab_6__5_) );
  NOR2_X1 U219 ( .A1(n12), .A2(n32), .ZN(ab_6__4_) );
  NOR2_X1 U220 ( .A1(n13), .A2(n32), .ZN(ab_6__3_) );
  NOR2_X1 U221 ( .A1(n14), .A2(n32), .ZN(ab_6__2_) );
  NOR2_X1 U222 ( .A1(A[6]), .A2(n1), .ZN(ab_6__23_) );
  NOR2_X1 U223 ( .A1(n15), .A2(n32), .ZN(ab_6__22_) );
  NOR2_X1 U224 ( .A1(n16), .A2(n32), .ZN(ab_6__21_) );
  NOR2_X1 U225 ( .A1(n17), .A2(n32), .ZN(ab_6__20_) );
  NOR2_X1 U226 ( .A1(n18), .A2(n32), .ZN(ab_6__1_) );
  NOR2_X1 U227 ( .A1(n19), .A2(n32), .ZN(ab_6__19_) );
  NOR2_X1 U228 ( .A1(n20), .A2(n32), .ZN(ab_6__18_) );
  NOR2_X1 U229 ( .A1(n21), .A2(n32), .ZN(ab_6__17_) );
  NOR2_X1 U230 ( .A1(n22), .A2(n32), .ZN(ab_6__16_) );
  NOR2_X1 U231 ( .A1(n23), .A2(n32), .ZN(ab_6__15_) );
  NOR2_X1 U232 ( .A1(n24), .A2(n32), .ZN(ab_6__14_) );
  NOR2_X1 U233 ( .A1(n25), .A2(n32), .ZN(ab_6__13_) );
  NOR2_X1 U234 ( .A1(n26), .A2(n32), .ZN(ab_6__12_) );
  NOR2_X1 U235 ( .A1(n27), .A2(n32), .ZN(ab_6__11_) );
  NOR2_X1 U236 ( .A1(n28), .A2(n32), .ZN(ab_6__10_) );
  NOR2_X1 U237 ( .A1(n29), .A2(n32), .ZN(ab_6__0_) );
  NOR2_X1 U238 ( .A1(n7), .A2(n33), .ZN(ab_5__9_) );
  NOR2_X1 U239 ( .A1(n8), .A2(n33), .ZN(ab_5__8_) );
  NOR2_X1 U240 ( .A1(n9), .A2(n33), .ZN(ab_5__7_) );
  NOR2_X1 U241 ( .A1(n10), .A2(n33), .ZN(ab_5__6_) );
  NOR2_X1 U242 ( .A1(n11), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U243 ( .A1(n12), .A2(n33), .ZN(ab_5__4_) );
  NOR2_X1 U244 ( .A1(n13), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U245 ( .A1(n14), .A2(n33), .ZN(ab_5__2_) );
  NOR2_X1 U246 ( .A1(A[5]), .A2(n1), .ZN(ab_5__23_) );
  NOR2_X1 U247 ( .A1(n15), .A2(n33), .ZN(ab_5__22_) );
  NOR2_X1 U248 ( .A1(n16), .A2(n33), .ZN(ab_5__21_) );
  NOR2_X1 U249 ( .A1(n17), .A2(n33), .ZN(ab_5__20_) );
  NOR2_X1 U250 ( .A1(n18), .A2(n33), .ZN(ab_5__1_) );
  NOR2_X1 U251 ( .A1(n19), .A2(n33), .ZN(ab_5__19_) );
  NOR2_X1 U252 ( .A1(n20), .A2(n33), .ZN(ab_5__18_) );
  NOR2_X1 U253 ( .A1(n21), .A2(n33), .ZN(ab_5__17_) );
  NOR2_X1 U254 ( .A1(n22), .A2(n33), .ZN(ab_5__16_) );
  NOR2_X1 U255 ( .A1(n23), .A2(n33), .ZN(ab_5__15_) );
  NOR2_X1 U256 ( .A1(n24), .A2(n33), .ZN(ab_5__14_) );
  NOR2_X1 U257 ( .A1(n25), .A2(n33), .ZN(ab_5__13_) );
  NOR2_X1 U258 ( .A1(n26), .A2(n33), .ZN(ab_5__12_) );
  NOR2_X1 U259 ( .A1(n27), .A2(n33), .ZN(ab_5__11_) );
  NOR2_X1 U260 ( .A1(n28), .A2(n33), .ZN(ab_5__10_) );
  NOR2_X1 U261 ( .A1(n29), .A2(n33), .ZN(ab_5__0_) );
  NOR2_X1 U262 ( .A1(n7), .A2(n34), .ZN(ab_4__9_) );
  NOR2_X1 U263 ( .A1(n8), .A2(n34), .ZN(ab_4__8_) );
  NOR2_X1 U264 ( .A1(n9), .A2(n34), .ZN(ab_4__7_) );
  NOR2_X1 U265 ( .A1(n10), .A2(n34), .ZN(ab_4__6_) );
  NOR2_X1 U266 ( .A1(n11), .A2(n34), .ZN(ab_4__5_) );
  NOR2_X1 U267 ( .A1(n12), .A2(n34), .ZN(ab_4__4_) );
  NOR2_X1 U268 ( .A1(n13), .A2(n34), .ZN(ab_4__3_) );
  NOR2_X1 U269 ( .A1(n14), .A2(n34), .ZN(ab_4__2_) );
  NOR2_X1 U270 ( .A1(A[4]), .A2(n1), .ZN(ab_4__23_) );
  NOR2_X1 U271 ( .A1(n15), .A2(n34), .ZN(ab_4__22_) );
  NOR2_X1 U272 ( .A1(n16), .A2(n34), .ZN(ab_4__21_) );
  NOR2_X1 U273 ( .A1(n17), .A2(n34), .ZN(ab_4__20_) );
  NOR2_X1 U274 ( .A1(n18), .A2(n34), .ZN(ab_4__1_) );
  NOR2_X1 U275 ( .A1(n19), .A2(n34), .ZN(ab_4__19_) );
  NOR2_X1 U276 ( .A1(n20), .A2(n34), .ZN(ab_4__18_) );
  NOR2_X1 U277 ( .A1(n21), .A2(n34), .ZN(ab_4__17_) );
  NOR2_X1 U278 ( .A1(n22), .A2(n34), .ZN(ab_4__16_) );
  NOR2_X1 U279 ( .A1(n23), .A2(n34), .ZN(ab_4__15_) );
  NOR2_X1 U280 ( .A1(n24), .A2(n34), .ZN(ab_4__14_) );
  NOR2_X1 U281 ( .A1(n25), .A2(n34), .ZN(ab_4__13_) );
  NOR2_X1 U282 ( .A1(n26), .A2(n34), .ZN(ab_4__12_) );
  NOR2_X1 U283 ( .A1(n27), .A2(n34), .ZN(ab_4__11_) );
  NOR2_X1 U284 ( .A1(n28), .A2(n34), .ZN(ab_4__10_) );
  NOR2_X1 U285 ( .A1(n29), .A2(n34), .ZN(ab_4__0_) );
  NOR2_X1 U286 ( .A1(n7), .A2(n35), .ZN(ab_3__9_) );
  NOR2_X1 U287 ( .A1(n8), .A2(n35), .ZN(ab_3__8_) );
  NOR2_X1 U288 ( .A1(n9), .A2(n35), .ZN(ab_3__7_) );
  NOR2_X1 U289 ( .A1(n10), .A2(n35), .ZN(ab_3__6_) );
  NOR2_X1 U290 ( .A1(n11), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U291 ( .A1(n12), .A2(n35), .ZN(ab_3__4_) );
  NOR2_X1 U292 ( .A1(n13), .A2(n35), .ZN(ab_3__3_) );
  NOR2_X1 U293 ( .A1(n14), .A2(n35), .ZN(ab_3__2_) );
  NOR2_X1 U294 ( .A1(A[3]), .A2(n1), .ZN(ab_3__23_) );
  NOR2_X1 U295 ( .A1(n15), .A2(n35), .ZN(ab_3__22_) );
  NOR2_X1 U296 ( .A1(n16), .A2(n35), .ZN(ab_3__21_) );
  NOR2_X1 U297 ( .A1(n17), .A2(n35), .ZN(ab_3__20_) );
  NOR2_X1 U298 ( .A1(n18), .A2(n35), .ZN(ab_3__1_) );
  NOR2_X1 U299 ( .A1(n19), .A2(n35), .ZN(ab_3__19_) );
  NOR2_X1 U300 ( .A1(n20), .A2(n35), .ZN(ab_3__18_) );
  NOR2_X1 U301 ( .A1(n21), .A2(n35), .ZN(ab_3__17_) );
  NOR2_X1 U302 ( .A1(n22), .A2(n35), .ZN(ab_3__16_) );
  NOR2_X1 U303 ( .A1(n23), .A2(n35), .ZN(ab_3__15_) );
  NOR2_X1 U304 ( .A1(n24), .A2(n35), .ZN(ab_3__14_) );
  NOR2_X1 U305 ( .A1(n25), .A2(n35), .ZN(ab_3__13_) );
  NOR2_X1 U306 ( .A1(n26), .A2(n35), .ZN(ab_3__12_) );
  NOR2_X1 U307 ( .A1(n27), .A2(n35), .ZN(ab_3__11_) );
  NOR2_X1 U308 ( .A1(n28), .A2(n35), .ZN(ab_3__10_) );
  NOR2_X1 U309 ( .A1(n29), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U310 ( .A1(n7), .A2(n36), .ZN(ab_2__9_) );
  NOR2_X1 U311 ( .A1(n8), .A2(n36), .ZN(ab_2__8_) );
  NOR2_X1 U312 ( .A1(n9), .A2(n36), .ZN(ab_2__7_) );
  NOR2_X1 U313 ( .A1(n10), .A2(n36), .ZN(ab_2__6_) );
  NOR2_X1 U314 ( .A1(n11), .A2(n36), .ZN(ab_2__5_) );
  NOR2_X1 U315 ( .A1(n12), .A2(n36), .ZN(ab_2__4_) );
  NOR2_X1 U316 ( .A1(n13), .A2(n36), .ZN(ab_2__3_) );
  NOR2_X1 U317 ( .A1(n14), .A2(n36), .ZN(ab_2__2_) );
  NOR2_X1 U318 ( .A1(A[2]), .A2(n1), .ZN(ab_2__23_) );
  NOR2_X1 U319 ( .A1(n15), .A2(n36), .ZN(ab_2__22_) );
  NOR2_X1 U320 ( .A1(n16), .A2(n36), .ZN(ab_2__21_) );
  NOR2_X1 U321 ( .A1(n17), .A2(n36), .ZN(ab_2__20_) );
  NOR2_X1 U322 ( .A1(n18), .A2(n36), .ZN(ab_2__1_) );
  NOR2_X1 U323 ( .A1(n19), .A2(n36), .ZN(ab_2__19_) );
  NOR2_X1 U324 ( .A1(n20), .A2(n36), .ZN(ab_2__18_) );
  NOR2_X1 U325 ( .A1(n21), .A2(n36), .ZN(ab_2__17_) );
  NOR2_X1 U326 ( .A1(n22), .A2(n36), .ZN(ab_2__16_) );
  NOR2_X1 U327 ( .A1(n23), .A2(n36), .ZN(ab_2__15_) );
  NOR2_X1 U328 ( .A1(n24), .A2(n36), .ZN(ab_2__14_) );
  NOR2_X1 U329 ( .A1(n25), .A2(n36), .ZN(ab_2__13_) );
  NOR2_X1 U330 ( .A1(n26), .A2(n36), .ZN(ab_2__12_) );
  NOR2_X1 U331 ( .A1(n27), .A2(n36), .ZN(ab_2__11_) );
  NOR2_X1 U332 ( .A1(n28), .A2(n36), .ZN(ab_2__10_) );
  NOR2_X1 U333 ( .A1(n29), .A2(n36), .ZN(ab_2__0_) );
  NOR2_X1 U334 ( .A1(B[9]), .A2(n4), .ZN(ab_23__9_) );
  NOR2_X1 U335 ( .A1(B[8]), .A2(n4), .ZN(ab_23__8_) );
  NOR2_X1 U336 ( .A1(B[7]), .A2(n4), .ZN(ab_23__7_) );
  NOR2_X1 U337 ( .A1(B[6]), .A2(n4), .ZN(ab_23__6_) );
  NOR2_X1 U338 ( .A1(B[5]), .A2(n3), .ZN(ab_23__5_) );
  NOR2_X1 U339 ( .A1(B[4]), .A2(n3), .ZN(ab_23__4_) );
  NOR2_X1 U340 ( .A1(B[3]), .A2(n3), .ZN(ab_23__3_) );
  NOR2_X1 U341 ( .A1(B[2]), .A2(n3), .ZN(ab_23__2_) );
  NOR2_X1 U342 ( .A1(n1), .A2(n3), .ZN(ab_23__23_) );
  NOR2_X1 U343 ( .A1(B[22]), .A2(n3), .ZN(ab_23__22_) );
  NOR2_X1 U344 ( .A1(B[21]), .A2(n3), .ZN(ab_23__21_) );
  NOR2_X1 U345 ( .A1(B[20]), .A2(n3), .ZN(ab_23__20_) );
  NOR2_X1 U346 ( .A1(B[1]), .A2(n3), .ZN(ab_23__1_) );
  NOR2_X1 U347 ( .A1(B[19]), .A2(n3), .ZN(ab_23__19_) );
  NOR2_X1 U348 ( .A1(B[18]), .A2(n3), .ZN(ab_23__18_) );
  NOR2_X1 U349 ( .A1(B[17]), .A2(n3), .ZN(ab_23__17_) );
  NOR2_X1 U350 ( .A1(B[16]), .A2(n3), .ZN(ab_23__16_) );
  NOR2_X1 U351 ( .A1(B[15]), .A2(n3), .ZN(ab_23__15_) );
  NOR2_X1 U352 ( .A1(B[14]), .A2(n3), .ZN(ab_23__14_) );
  NOR2_X1 U353 ( .A1(B[13]), .A2(n3), .ZN(ab_23__13_) );
  NOR2_X1 U354 ( .A1(B[12]), .A2(n3), .ZN(ab_23__12_) );
  NOR2_X1 U355 ( .A1(B[11]), .A2(n3), .ZN(ab_23__11_) );
  NOR2_X1 U356 ( .A1(B[10]), .A2(n3), .ZN(ab_23__10_) );
  NOR2_X1 U357 ( .A1(B[0]), .A2(n3), .ZN(ab_23__0_) );
  NOR2_X1 U358 ( .A1(n7), .A2(n37), .ZN(ab_22__9_) );
  NOR2_X1 U359 ( .A1(n8), .A2(n37), .ZN(ab_22__8_) );
  NOR2_X1 U360 ( .A1(n9), .A2(n37), .ZN(ab_22__7_) );
  NOR2_X1 U361 ( .A1(n10), .A2(n37), .ZN(ab_22__6_) );
  NOR2_X1 U362 ( .A1(n11), .A2(n37), .ZN(ab_22__5_) );
  NOR2_X1 U363 ( .A1(n12), .A2(n37), .ZN(ab_22__4_) );
  NOR2_X1 U364 ( .A1(n13), .A2(n37), .ZN(ab_22__3_) );
  NOR2_X1 U365 ( .A1(n14), .A2(n37), .ZN(ab_22__2_) );
  NOR2_X1 U366 ( .A1(A[22]), .A2(n1), .ZN(ab_22__23_) );
  NOR2_X1 U367 ( .A1(n15), .A2(n37), .ZN(ab_22__22_) );
  NOR2_X1 U368 ( .A1(n16), .A2(n37), .ZN(ab_22__21_) );
  NOR2_X1 U369 ( .A1(n17), .A2(n37), .ZN(ab_22__20_) );
  NOR2_X1 U370 ( .A1(n18), .A2(n37), .ZN(ab_22__1_) );
  NOR2_X1 U371 ( .A1(n19), .A2(n37), .ZN(ab_22__19_) );
  NOR2_X1 U372 ( .A1(n20), .A2(n37), .ZN(ab_22__18_) );
  NOR2_X1 U373 ( .A1(n21), .A2(n37), .ZN(ab_22__17_) );
  NOR2_X1 U374 ( .A1(n22), .A2(n37), .ZN(ab_22__16_) );
  NOR2_X1 U375 ( .A1(n23), .A2(n37), .ZN(ab_22__15_) );
  NOR2_X1 U376 ( .A1(n24), .A2(n37), .ZN(ab_22__14_) );
  NOR2_X1 U377 ( .A1(n25), .A2(n37), .ZN(ab_22__13_) );
  NOR2_X1 U378 ( .A1(n26), .A2(n37), .ZN(ab_22__12_) );
  NOR2_X1 U379 ( .A1(n27), .A2(n37), .ZN(ab_22__11_) );
  NOR2_X1 U380 ( .A1(n28), .A2(n37), .ZN(ab_22__10_) );
  NOR2_X1 U381 ( .A1(n29), .A2(n37), .ZN(ab_22__0_) );
  NOR2_X1 U382 ( .A1(n7), .A2(n38), .ZN(ab_21__9_) );
  NOR2_X1 U383 ( .A1(n8), .A2(n38), .ZN(ab_21__8_) );
  NOR2_X1 U384 ( .A1(n9), .A2(n38), .ZN(ab_21__7_) );
  NOR2_X1 U385 ( .A1(n10), .A2(n38), .ZN(ab_21__6_) );
  NOR2_X1 U386 ( .A1(n11), .A2(n38), .ZN(ab_21__5_) );
  NOR2_X1 U387 ( .A1(n12), .A2(n38), .ZN(ab_21__4_) );
  NOR2_X1 U388 ( .A1(n13), .A2(n38), .ZN(ab_21__3_) );
  NOR2_X1 U389 ( .A1(n14), .A2(n38), .ZN(ab_21__2_) );
  NOR2_X1 U390 ( .A1(A[21]), .A2(n1), .ZN(ab_21__23_) );
  NOR2_X1 U391 ( .A1(n15), .A2(n38), .ZN(ab_21__22_) );
  NOR2_X1 U392 ( .A1(n16), .A2(n38), .ZN(ab_21__21_) );
  NOR2_X1 U393 ( .A1(n17), .A2(n38), .ZN(ab_21__20_) );
  NOR2_X1 U394 ( .A1(n18), .A2(n38), .ZN(ab_21__1_) );
  NOR2_X1 U395 ( .A1(n19), .A2(n38), .ZN(ab_21__19_) );
  NOR2_X1 U396 ( .A1(n20), .A2(n38), .ZN(ab_21__18_) );
  NOR2_X1 U397 ( .A1(n21), .A2(n38), .ZN(ab_21__17_) );
  NOR2_X1 U398 ( .A1(n22), .A2(n38), .ZN(ab_21__16_) );
  NOR2_X1 U399 ( .A1(n23), .A2(n38), .ZN(ab_21__15_) );
  NOR2_X1 U400 ( .A1(n24), .A2(n38), .ZN(ab_21__14_) );
  NOR2_X1 U401 ( .A1(n25), .A2(n38), .ZN(ab_21__13_) );
  NOR2_X1 U402 ( .A1(n26), .A2(n38), .ZN(ab_21__12_) );
  NOR2_X1 U403 ( .A1(n27), .A2(n38), .ZN(ab_21__11_) );
  NOR2_X1 U404 ( .A1(n28), .A2(n38), .ZN(ab_21__10_) );
  NOR2_X1 U405 ( .A1(n29), .A2(n38), .ZN(ab_21__0_) );
  NOR2_X1 U406 ( .A1(n7), .A2(n39), .ZN(ab_20__9_) );
  NOR2_X1 U407 ( .A1(n8), .A2(n39), .ZN(ab_20__8_) );
  NOR2_X1 U408 ( .A1(n9), .A2(n39), .ZN(ab_20__7_) );
  NOR2_X1 U409 ( .A1(n10), .A2(n39), .ZN(ab_20__6_) );
  NOR2_X1 U410 ( .A1(n11), .A2(n39), .ZN(ab_20__5_) );
  NOR2_X1 U411 ( .A1(n12), .A2(n39), .ZN(ab_20__4_) );
  NOR2_X1 U412 ( .A1(n13), .A2(n39), .ZN(ab_20__3_) );
  NOR2_X1 U413 ( .A1(n14), .A2(n39), .ZN(ab_20__2_) );
  NOR2_X1 U414 ( .A1(A[20]), .A2(n1), .ZN(ab_20__23_) );
  NOR2_X1 U415 ( .A1(n15), .A2(n39), .ZN(ab_20__22_) );
  NOR2_X1 U416 ( .A1(n16), .A2(n39), .ZN(ab_20__21_) );
  NOR2_X1 U417 ( .A1(n17), .A2(n39), .ZN(ab_20__20_) );
  NOR2_X1 U418 ( .A1(n18), .A2(n39), .ZN(ab_20__1_) );
  NOR2_X1 U419 ( .A1(n19), .A2(n39), .ZN(ab_20__19_) );
  NOR2_X1 U420 ( .A1(n20), .A2(n39), .ZN(ab_20__18_) );
  NOR2_X1 U421 ( .A1(n21), .A2(n39), .ZN(ab_20__17_) );
  NOR2_X1 U422 ( .A1(n22), .A2(n39), .ZN(ab_20__16_) );
  NOR2_X1 U423 ( .A1(n23), .A2(n39), .ZN(ab_20__15_) );
  NOR2_X1 U424 ( .A1(n24), .A2(n39), .ZN(ab_20__14_) );
  NOR2_X1 U425 ( .A1(n25), .A2(n39), .ZN(ab_20__13_) );
  NOR2_X1 U426 ( .A1(n26), .A2(n39), .ZN(ab_20__12_) );
  NOR2_X1 U427 ( .A1(n27), .A2(n39), .ZN(ab_20__11_) );
  NOR2_X1 U428 ( .A1(n28), .A2(n39), .ZN(ab_20__10_) );
  NOR2_X1 U429 ( .A1(n29), .A2(n39), .ZN(ab_20__0_) );
  NOR2_X1 U430 ( .A1(n7), .A2(n40), .ZN(ab_1__9_) );
  NOR2_X1 U431 ( .A1(n8), .A2(n40), .ZN(ab_1__8_) );
  NOR2_X1 U432 ( .A1(n9), .A2(n40), .ZN(ab_1__7_) );
  NOR2_X1 U433 ( .A1(n10), .A2(n40), .ZN(ab_1__6_) );
  NOR2_X1 U434 ( .A1(n11), .A2(n40), .ZN(ab_1__5_) );
  NOR2_X1 U435 ( .A1(n12), .A2(n40), .ZN(ab_1__4_) );
  NOR2_X1 U436 ( .A1(n13), .A2(n40), .ZN(ab_1__3_) );
  NOR2_X1 U437 ( .A1(n14), .A2(n40), .ZN(ab_1__2_) );
  NOR2_X1 U438 ( .A1(A[1]), .A2(n1), .ZN(ab_1__23_) );
  NOR2_X1 U439 ( .A1(n15), .A2(n40), .ZN(ab_1__22_) );
  NOR2_X1 U440 ( .A1(n16), .A2(n40), .ZN(ab_1__21_) );
  NOR2_X1 U441 ( .A1(n17), .A2(n40), .ZN(ab_1__20_) );
  NOR2_X1 U442 ( .A1(n19), .A2(n40), .ZN(ab_1__19_) );
  NOR2_X1 U443 ( .A1(n20), .A2(n40), .ZN(ab_1__18_) );
  NOR2_X1 U444 ( .A1(n21), .A2(n40), .ZN(ab_1__17_) );
  NOR2_X1 U445 ( .A1(n22), .A2(n40), .ZN(ab_1__16_) );
  NOR2_X1 U446 ( .A1(n23), .A2(n40), .ZN(ab_1__15_) );
  NOR2_X1 U447 ( .A1(n24), .A2(n40), .ZN(ab_1__14_) );
  NOR2_X1 U448 ( .A1(n25), .A2(n40), .ZN(ab_1__13_) );
  NOR2_X1 U449 ( .A1(n26), .A2(n40), .ZN(ab_1__12_) );
  NOR2_X1 U450 ( .A1(n27), .A2(n40), .ZN(ab_1__11_) );
  NOR2_X1 U451 ( .A1(n28), .A2(n40), .ZN(ab_1__10_) );
  NOR2_X1 U452 ( .A1(n7), .A2(n41), .ZN(ab_19__9_) );
  NOR2_X1 U453 ( .A1(n8), .A2(n41), .ZN(ab_19__8_) );
  NOR2_X1 U454 ( .A1(n9), .A2(n41), .ZN(ab_19__7_) );
  NOR2_X1 U455 ( .A1(n10), .A2(n41), .ZN(ab_19__6_) );
  NOR2_X1 U456 ( .A1(n11), .A2(n41), .ZN(ab_19__5_) );
  NOR2_X1 U457 ( .A1(n12), .A2(n41), .ZN(ab_19__4_) );
  NOR2_X1 U458 ( .A1(n13), .A2(n41), .ZN(ab_19__3_) );
  NOR2_X1 U459 ( .A1(n14), .A2(n41), .ZN(ab_19__2_) );
  NOR2_X1 U460 ( .A1(A[19]), .A2(n1), .ZN(ab_19__23_) );
  NOR2_X1 U461 ( .A1(n15), .A2(n41), .ZN(ab_19__22_) );
  NOR2_X1 U462 ( .A1(n16), .A2(n41), .ZN(ab_19__21_) );
  NOR2_X1 U463 ( .A1(n17), .A2(n41), .ZN(ab_19__20_) );
  NOR2_X1 U464 ( .A1(n18), .A2(n41), .ZN(ab_19__1_) );
  NOR2_X1 U465 ( .A1(n19), .A2(n41), .ZN(ab_19__19_) );
  NOR2_X1 U466 ( .A1(n20), .A2(n41), .ZN(ab_19__18_) );
  NOR2_X1 U467 ( .A1(n21), .A2(n41), .ZN(ab_19__17_) );
  NOR2_X1 U468 ( .A1(n22), .A2(n41), .ZN(ab_19__16_) );
  NOR2_X1 U469 ( .A1(n23), .A2(n41), .ZN(ab_19__15_) );
  NOR2_X1 U470 ( .A1(n24), .A2(n41), .ZN(ab_19__14_) );
  NOR2_X1 U471 ( .A1(n25), .A2(n41), .ZN(ab_19__13_) );
  NOR2_X1 U472 ( .A1(n26), .A2(n41), .ZN(ab_19__12_) );
  NOR2_X1 U473 ( .A1(n27), .A2(n41), .ZN(ab_19__11_) );
  NOR2_X1 U474 ( .A1(n28), .A2(n41), .ZN(ab_19__10_) );
  NOR2_X1 U475 ( .A1(n29), .A2(n41), .ZN(ab_19__0_) );
  NOR2_X1 U476 ( .A1(n7), .A2(n42), .ZN(ab_18__9_) );
  NOR2_X1 U477 ( .A1(n8), .A2(n42), .ZN(ab_18__8_) );
  NOR2_X1 U478 ( .A1(n9), .A2(n42), .ZN(ab_18__7_) );
  NOR2_X1 U479 ( .A1(n10), .A2(n42), .ZN(ab_18__6_) );
  NOR2_X1 U480 ( .A1(n11), .A2(n42), .ZN(ab_18__5_) );
  NOR2_X1 U481 ( .A1(n12), .A2(n42), .ZN(ab_18__4_) );
  NOR2_X1 U482 ( .A1(n13), .A2(n42), .ZN(ab_18__3_) );
  NOR2_X1 U483 ( .A1(n14), .A2(n42), .ZN(ab_18__2_) );
  NOR2_X1 U484 ( .A1(A[18]), .A2(n1), .ZN(ab_18__23_) );
  NOR2_X1 U485 ( .A1(n15), .A2(n42), .ZN(ab_18__22_) );
  NOR2_X1 U486 ( .A1(n16), .A2(n42), .ZN(ab_18__21_) );
  NOR2_X1 U487 ( .A1(n17), .A2(n42), .ZN(ab_18__20_) );
  NOR2_X1 U488 ( .A1(n18), .A2(n42), .ZN(ab_18__1_) );
  NOR2_X1 U489 ( .A1(n19), .A2(n42), .ZN(ab_18__19_) );
  NOR2_X1 U490 ( .A1(n20), .A2(n42), .ZN(ab_18__18_) );
  NOR2_X1 U491 ( .A1(n21), .A2(n42), .ZN(ab_18__17_) );
  NOR2_X1 U492 ( .A1(n22), .A2(n42), .ZN(ab_18__16_) );
  NOR2_X1 U493 ( .A1(n23), .A2(n42), .ZN(ab_18__15_) );
  NOR2_X1 U494 ( .A1(n24), .A2(n42), .ZN(ab_18__14_) );
  NOR2_X1 U495 ( .A1(n25), .A2(n42), .ZN(ab_18__13_) );
  NOR2_X1 U496 ( .A1(n26), .A2(n42), .ZN(ab_18__12_) );
  NOR2_X1 U497 ( .A1(n27), .A2(n42), .ZN(ab_18__11_) );
  NOR2_X1 U498 ( .A1(n28), .A2(n42), .ZN(ab_18__10_) );
  NOR2_X1 U499 ( .A1(n29), .A2(n42), .ZN(ab_18__0_) );
  NOR2_X1 U500 ( .A1(n7), .A2(n43), .ZN(ab_17__9_) );
  NOR2_X1 U501 ( .A1(n8), .A2(n43), .ZN(ab_17__8_) );
  NOR2_X1 U502 ( .A1(n9), .A2(n43), .ZN(ab_17__7_) );
  NOR2_X1 U503 ( .A1(n10), .A2(n43), .ZN(ab_17__6_) );
  NOR2_X1 U504 ( .A1(n11), .A2(n43), .ZN(ab_17__5_) );
  NOR2_X1 U505 ( .A1(n12), .A2(n43), .ZN(ab_17__4_) );
  NOR2_X1 U506 ( .A1(n13), .A2(n43), .ZN(ab_17__3_) );
  NOR2_X1 U507 ( .A1(n14), .A2(n43), .ZN(ab_17__2_) );
  NOR2_X1 U508 ( .A1(A[17]), .A2(n1), .ZN(ab_17__23_) );
  NOR2_X1 U509 ( .A1(n15), .A2(n43), .ZN(ab_17__22_) );
  NOR2_X1 U510 ( .A1(n16), .A2(n43), .ZN(ab_17__21_) );
  NOR2_X1 U511 ( .A1(n17), .A2(n43), .ZN(ab_17__20_) );
  NOR2_X1 U512 ( .A1(n18), .A2(n43), .ZN(ab_17__1_) );
  NOR2_X1 U513 ( .A1(n19), .A2(n43), .ZN(ab_17__19_) );
  NOR2_X1 U514 ( .A1(n20), .A2(n43), .ZN(ab_17__18_) );
  NOR2_X1 U515 ( .A1(n21), .A2(n43), .ZN(ab_17__17_) );
  NOR2_X1 U516 ( .A1(n22), .A2(n43), .ZN(ab_17__16_) );
  NOR2_X1 U517 ( .A1(n23), .A2(n43), .ZN(ab_17__15_) );
  NOR2_X1 U518 ( .A1(n24), .A2(n43), .ZN(ab_17__14_) );
  NOR2_X1 U519 ( .A1(n25), .A2(n43), .ZN(ab_17__13_) );
  NOR2_X1 U520 ( .A1(n26), .A2(n43), .ZN(ab_17__12_) );
  NOR2_X1 U521 ( .A1(n27), .A2(n43), .ZN(ab_17__11_) );
  NOR2_X1 U522 ( .A1(n28), .A2(n43), .ZN(ab_17__10_) );
  NOR2_X1 U523 ( .A1(n29), .A2(n43), .ZN(ab_17__0_) );
  NOR2_X1 U524 ( .A1(n7), .A2(n44), .ZN(ab_16__9_) );
  NOR2_X1 U525 ( .A1(n8), .A2(n44), .ZN(ab_16__8_) );
  NOR2_X1 U526 ( .A1(n9), .A2(n44), .ZN(ab_16__7_) );
  NOR2_X1 U527 ( .A1(n10), .A2(n44), .ZN(ab_16__6_) );
  NOR2_X1 U528 ( .A1(n11), .A2(n44), .ZN(ab_16__5_) );
  NOR2_X1 U529 ( .A1(n12), .A2(n44), .ZN(ab_16__4_) );
  NOR2_X1 U530 ( .A1(n13), .A2(n44), .ZN(ab_16__3_) );
  NOR2_X1 U531 ( .A1(n14), .A2(n44), .ZN(ab_16__2_) );
  NOR2_X1 U532 ( .A1(A[16]), .A2(n1), .ZN(ab_16__23_) );
  NOR2_X1 U533 ( .A1(n15), .A2(n44), .ZN(ab_16__22_) );
  NOR2_X1 U534 ( .A1(n16), .A2(n44), .ZN(ab_16__21_) );
  NOR2_X1 U535 ( .A1(n17), .A2(n44), .ZN(ab_16__20_) );
  NOR2_X1 U536 ( .A1(n18), .A2(n44), .ZN(ab_16__1_) );
  NOR2_X1 U537 ( .A1(n19), .A2(n44), .ZN(ab_16__19_) );
  NOR2_X1 U538 ( .A1(n20), .A2(n44), .ZN(ab_16__18_) );
  NOR2_X1 U539 ( .A1(n21), .A2(n44), .ZN(ab_16__17_) );
  NOR2_X1 U540 ( .A1(n22), .A2(n44), .ZN(ab_16__16_) );
  NOR2_X1 U541 ( .A1(n23), .A2(n44), .ZN(ab_16__15_) );
  NOR2_X1 U542 ( .A1(n24), .A2(n44), .ZN(ab_16__14_) );
  NOR2_X1 U543 ( .A1(n25), .A2(n44), .ZN(ab_16__13_) );
  NOR2_X1 U544 ( .A1(n26), .A2(n44), .ZN(ab_16__12_) );
  NOR2_X1 U545 ( .A1(n27), .A2(n44), .ZN(ab_16__11_) );
  NOR2_X1 U546 ( .A1(n28), .A2(n44), .ZN(ab_16__10_) );
  NOR2_X1 U547 ( .A1(n29), .A2(n44), .ZN(ab_16__0_) );
  NOR2_X1 U548 ( .A1(n7), .A2(n45), .ZN(ab_15__9_) );
  NOR2_X1 U549 ( .A1(n8), .A2(n45), .ZN(ab_15__8_) );
  NOR2_X1 U550 ( .A1(n9), .A2(n45), .ZN(ab_15__7_) );
  NOR2_X1 U551 ( .A1(n10), .A2(n45), .ZN(ab_15__6_) );
  NOR2_X1 U552 ( .A1(n11), .A2(n45), .ZN(ab_15__5_) );
  NOR2_X1 U553 ( .A1(n12), .A2(n45), .ZN(ab_15__4_) );
  NOR2_X1 U554 ( .A1(n13), .A2(n45), .ZN(ab_15__3_) );
  NOR2_X1 U555 ( .A1(n14), .A2(n45), .ZN(ab_15__2_) );
  NOR2_X1 U556 ( .A1(A[15]), .A2(n1), .ZN(ab_15__23_) );
  NOR2_X1 U557 ( .A1(n15), .A2(n45), .ZN(ab_15__22_) );
  NOR2_X1 U558 ( .A1(n16), .A2(n45), .ZN(ab_15__21_) );
  NOR2_X1 U559 ( .A1(n17), .A2(n45), .ZN(ab_15__20_) );
  NOR2_X1 U560 ( .A1(n18), .A2(n45), .ZN(ab_15__1_) );
  NOR2_X1 U561 ( .A1(n19), .A2(n45), .ZN(ab_15__19_) );
  NOR2_X1 U562 ( .A1(n20), .A2(n45), .ZN(ab_15__18_) );
  NOR2_X1 U563 ( .A1(n21), .A2(n45), .ZN(ab_15__17_) );
  NOR2_X1 U564 ( .A1(n22), .A2(n45), .ZN(ab_15__16_) );
  NOR2_X1 U565 ( .A1(n23), .A2(n45), .ZN(ab_15__15_) );
  NOR2_X1 U566 ( .A1(n24), .A2(n45), .ZN(ab_15__14_) );
  NOR2_X1 U567 ( .A1(n25), .A2(n45), .ZN(ab_15__13_) );
  NOR2_X1 U568 ( .A1(n26), .A2(n45), .ZN(ab_15__12_) );
  NOR2_X1 U569 ( .A1(n27), .A2(n45), .ZN(ab_15__11_) );
  NOR2_X1 U570 ( .A1(n28), .A2(n45), .ZN(ab_15__10_) );
  NOR2_X1 U571 ( .A1(n29), .A2(n45), .ZN(ab_15__0_) );
  NOR2_X1 U572 ( .A1(n7), .A2(n46), .ZN(ab_14__9_) );
  NOR2_X1 U573 ( .A1(n8), .A2(n46), .ZN(ab_14__8_) );
  NOR2_X1 U574 ( .A1(n9), .A2(n46), .ZN(ab_14__7_) );
  NOR2_X1 U575 ( .A1(n10), .A2(n46), .ZN(ab_14__6_) );
  NOR2_X1 U576 ( .A1(n11), .A2(n46), .ZN(ab_14__5_) );
  NOR2_X1 U577 ( .A1(n12), .A2(n46), .ZN(ab_14__4_) );
  NOR2_X1 U578 ( .A1(n13), .A2(n46), .ZN(ab_14__3_) );
  NOR2_X1 U579 ( .A1(n14), .A2(n46), .ZN(ab_14__2_) );
  NOR2_X1 U580 ( .A1(A[14]), .A2(n2), .ZN(ab_14__23_) );
  NOR2_X1 U581 ( .A1(n15), .A2(n46), .ZN(ab_14__22_) );
  NOR2_X1 U582 ( .A1(n16), .A2(n46), .ZN(ab_14__21_) );
  NOR2_X1 U583 ( .A1(n17), .A2(n46), .ZN(ab_14__20_) );
  NOR2_X1 U584 ( .A1(n18), .A2(n46), .ZN(ab_14__1_) );
  NOR2_X1 U585 ( .A1(n19), .A2(n46), .ZN(ab_14__19_) );
  NOR2_X1 U586 ( .A1(n20), .A2(n46), .ZN(ab_14__18_) );
  NOR2_X1 U587 ( .A1(n21), .A2(n46), .ZN(ab_14__17_) );
  NOR2_X1 U588 ( .A1(n22), .A2(n46), .ZN(ab_14__16_) );
  NOR2_X1 U589 ( .A1(n23), .A2(n46), .ZN(ab_14__15_) );
  NOR2_X1 U590 ( .A1(n24), .A2(n46), .ZN(ab_14__14_) );
  NOR2_X1 U591 ( .A1(n25), .A2(n46), .ZN(ab_14__13_) );
  NOR2_X1 U592 ( .A1(n26), .A2(n46), .ZN(ab_14__12_) );
  NOR2_X1 U593 ( .A1(n27), .A2(n46), .ZN(ab_14__11_) );
  NOR2_X1 U594 ( .A1(n28), .A2(n46), .ZN(ab_14__10_) );
  NOR2_X1 U595 ( .A1(n29), .A2(n46), .ZN(ab_14__0_) );
  NOR2_X1 U596 ( .A1(n7), .A2(n47), .ZN(ab_13__9_) );
  NOR2_X1 U597 ( .A1(n8), .A2(n47), .ZN(ab_13__8_) );
  NOR2_X1 U598 ( .A1(n9), .A2(n47), .ZN(ab_13__7_) );
  NOR2_X1 U599 ( .A1(n10), .A2(n47), .ZN(ab_13__6_) );
  NOR2_X1 U600 ( .A1(n11), .A2(n47), .ZN(ab_13__5_) );
  NOR2_X1 U601 ( .A1(n12), .A2(n47), .ZN(ab_13__4_) );
  NOR2_X1 U602 ( .A1(n13), .A2(n47), .ZN(ab_13__3_) );
  NOR2_X1 U603 ( .A1(n14), .A2(n47), .ZN(ab_13__2_) );
  NOR2_X1 U604 ( .A1(A[13]), .A2(n2), .ZN(ab_13__23_) );
  NOR2_X1 U605 ( .A1(n15), .A2(n47), .ZN(ab_13__22_) );
  NOR2_X1 U606 ( .A1(n16), .A2(n47), .ZN(ab_13__21_) );
  NOR2_X1 U607 ( .A1(n17), .A2(n47), .ZN(ab_13__20_) );
  NOR2_X1 U608 ( .A1(n18), .A2(n47), .ZN(ab_13__1_) );
  NOR2_X1 U609 ( .A1(n19), .A2(n47), .ZN(ab_13__19_) );
  NOR2_X1 U610 ( .A1(n20), .A2(n47), .ZN(ab_13__18_) );
  NOR2_X1 U611 ( .A1(n21), .A2(n47), .ZN(ab_13__17_) );
  NOR2_X1 U612 ( .A1(n22), .A2(n47), .ZN(ab_13__16_) );
  NOR2_X1 U613 ( .A1(n23), .A2(n47), .ZN(ab_13__15_) );
  NOR2_X1 U614 ( .A1(n24), .A2(n47), .ZN(ab_13__14_) );
  NOR2_X1 U615 ( .A1(n25), .A2(n47), .ZN(ab_13__13_) );
  NOR2_X1 U616 ( .A1(n26), .A2(n47), .ZN(ab_13__12_) );
  NOR2_X1 U617 ( .A1(n27), .A2(n47), .ZN(ab_13__11_) );
  NOR2_X1 U618 ( .A1(n28), .A2(n47), .ZN(ab_13__10_) );
  NOR2_X1 U619 ( .A1(n29), .A2(n47), .ZN(ab_13__0_) );
  NOR2_X1 U620 ( .A1(n7), .A2(n48), .ZN(ab_12__9_) );
  NOR2_X1 U621 ( .A1(n8), .A2(n48), .ZN(ab_12__8_) );
  NOR2_X1 U622 ( .A1(n9), .A2(n48), .ZN(ab_12__7_) );
  NOR2_X1 U623 ( .A1(n10), .A2(n48), .ZN(ab_12__6_) );
  NOR2_X1 U624 ( .A1(n11), .A2(n48), .ZN(ab_12__5_) );
  NOR2_X1 U625 ( .A1(n12), .A2(n48), .ZN(ab_12__4_) );
  NOR2_X1 U626 ( .A1(n13), .A2(n48), .ZN(ab_12__3_) );
  NOR2_X1 U627 ( .A1(n14), .A2(n48), .ZN(ab_12__2_) );
  NOR2_X1 U628 ( .A1(A[12]), .A2(n2), .ZN(ab_12__23_) );
  NOR2_X1 U629 ( .A1(n15), .A2(n48), .ZN(ab_12__22_) );
  NOR2_X1 U630 ( .A1(n16), .A2(n48), .ZN(ab_12__21_) );
  NOR2_X1 U631 ( .A1(n17), .A2(n48), .ZN(ab_12__20_) );
  NOR2_X1 U632 ( .A1(n18), .A2(n48), .ZN(ab_12__1_) );
  NOR2_X1 U633 ( .A1(n19), .A2(n48), .ZN(ab_12__19_) );
  NOR2_X1 U634 ( .A1(n20), .A2(n48), .ZN(ab_12__18_) );
  NOR2_X1 U635 ( .A1(n21), .A2(n48), .ZN(ab_12__17_) );
  NOR2_X1 U636 ( .A1(n22), .A2(n48), .ZN(ab_12__16_) );
  NOR2_X1 U637 ( .A1(n23), .A2(n48), .ZN(ab_12__15_) );
  NOR2_X1 U638 ( .A1(n24), .A2(n48), .ZN(ab_12__14_) );
  NOR2_X1 U639 ( .A1(n25), .A2(n48), .ZN(ab_12__13_) );
  NOR2_X1 U640 ( .A1(n26), .A2(n48), .ZN(ab_12__12_) );
  NOR2_X1 U641 ( .A1(n27), .A2(n48), .ZN(ab_12__11_) );
  NOR2_X1 U642 ( .A1(n28), .A2(n48), .ZN(ab_12__10_) );
  NOR2_X1 U643 ( .A1(n29), .A2(n48), .ZN(ab_12__0_) );
  NOR2_X1 U644 ( .A1(n7), .A2(n49), .ZN(ab_11__9_) );
  NOR2_X1 U645 ( .A1(n8), .A2(n49), .ZN(ab_11__8_) );
  NOR2_X1 U646 ( .A1(n9), .A2(n49), .ZN(ab_11__7_) );
  NOR2_X1 U647 ( .A1(n10), .A2(n49), .ZN(ab_11__6_) );
  NOR2_X1 U648 ( .A1(n11), .A2(n49), .ZN(ab_11__5_) );
  NOR2_X1 U649 ( .A1(n12), .A2(n49), .ZN(ab_11__4_) );
  NOR2_X1 U650 ( .A1(n13), .A2(n49), .ZN(ab_11__3_) );
  NOR2_X1 U651 ( .A1(n14), .A2(n49), .ZN(ab_11__2_) );
  NOR2_X1 U652 ( .A1(A[11]), .A2(n2), .ZN(ab_11__23_) );
  NOR2_X1 U653 ( .A1(n15), .A2(n49), .ZN(ab_11__22_) );
  NOR2_X1 U654 ( .A1(n16), .A2(n49), .ZN(ab_11__21_) );
  NOR2_X1 U655 ( .A1(n17), .A2(n49), .ZN(ab_11__20_) );
  NOR2_X1 U656 ( .A1(n18), .A2(n49), .ZN(ab_11__1_) );
  NOR2_X1 U657 ( .A1(n19), .A2(n49), .ZN(ab_11__19_) );
  NOR2_X1 U658 ( .A1(n20), .A2(n49), .ZN(ab_11__18_) );
  NOR2_X1 U659 ( .A1(n21), .A2(n49), .ZN(ab_11__17_) );
  NOR2_X1 U660 ( .A1(n22), .A2(n49), .ZN(ab_11__16_) );
  NOR2_X1 U661 ( .A1(n23), .A2(n49), .ZN(ab_11__15_) );
  NOR2_X1 U662 ( .A1(n24), .A2(n49), .ZN(ab_11__14_) );
  NOR2_X1 U663 ( .A1(n25), .A2(n49), .ZN(ab_11__13_) );
  NOR2_X1 U664 ( .A1(n26), .A2(n49), .ZN(ab_11__12_) );
  NOR2_X1 U665 ( .A1(n27), .A2(n49), .ZN(ab_11__11_) );
  NOR2_X1 U666 ( .A1(n28), .A2(n49), .ZN(ab_11__10_) );
  NOR2_X1 U667 ( .A1(n29), .A2(n49), .ZN(ab_11__0_) );
  NOR2_X1 U668 ( .A1(n7), .A2(n50), .ZN(ab_10__9_) );
  NOR2_X1 U669 ( .A1(n8), .A2(n50), .ZN(ab_10__8_) );
  NOR2_X1 U670 ( .A1(n9), .A2(n50), .ZN(ab_10__7_) );
  NOR2_X1 U671 ( .A1(n10), .A2(n50), .ZN(ab_10__6_) );
  NOR2_X1 U672 ( .A1(n11), .A2(n50), .ZN(ab_10__5_) );
  NOR2_X1 U673 ( .A1(n12), .A2(n50), .ZN(ab_10__4_) );
  NOR2_X1 U674 ( .A1(n13), .A2(n50), .ZN(ab_10__3_) );
  NOR2_X1 U675 ( .A1(n14), .A2(n50), .ZN(ab_10__2_) );
  NOR2_X1 U676 ( .A1(A[10]), .A2(n2), .ZN(ab_10__23_) );
  NOR2_X1 U677 ( .A1(n15), .A2(n50), .ZN(ab_10__22_) );
  NOR2_X1 U678 ( .A1(n16), .A2(n50), .ZN(ab_10__21_) );
  NOR2_X1 U679 ( .A1(n17), .A2(n50), .ZN(ab_10__20_) );
  NOR2_X1 U680 ( .A1(n18), .A2(n50), .ZN(ab_10__1_) );
  NOR2_X1 U681 ( .A1(n19), .A2(n50), .ZN(ab_10__19_) );
  NOR2_X1 U682 ( .A1(n20), .A2(n50), .ZN(ab_10__18_) );
  NOR2_X1 U683 ( .A1(n21), .A2(n50), .ZN(ab_10__17_) );
  NOR2_X1 U684 ( .A1(n22), .A2(n50), .ZN(ab_10__16_) );
  NOR2_X1 U685 ( .A1(n23), .A2(n50), .ZN(ab_10__15_) );
  NOR2_X1 U686 ( .A1(n24), .A2(n50), .ZN(ab_10__14_) );
  NOR2_X1 U687 ( .A1(n25), .A2(n50), .ZN(ab_10__13_) );
  NOR2_X1 U688 ( .A1(n26), .A2(n50), .ZN(ab_10__12_) );
  NOR2_X1 U689 ( .A1(n27), .A2(n50), .ZN(ab_10__11_) );
  NOR2_X1 U690 ( .A1(n28), .A2(n50), .ZN(ab_10__10_) );
  NOR2_X1 U691 ( .A1(n29), .A2(n50), .ZN(ab_10__0_) );
  NOR2_X1 U692 ( .A1(n7), .A2(n51), .ZN(ab_0__9_) );
  NOR2_X1 U693 ( .A1(n8), .A2(n51), .ZN(ab_0__8_) );
  NOR2_X1 U694 ( .A1(n9), .A2(n51), .ZN(ab_0__7_) );
  NOR2_X1 U695 ( .A1(n10), .A2(n51), .ZN(ab_0__6_) );
  NOR2_X1 U696 ( .A1(n11), .A2(n51), .ZN(ab_0__5_) );
  NOR2_X1 U697 ( .A1(n12), .A2(n51), .ZN(ab_0__4_) );
  NOR2_X1 U698 ( .A1(n13), .A2(n51), .ZN(ab_0__3_) );
  NOR2_X1 U699 ( .A1(n14), .A2(n51), .ZN(ab_0__2_) );
  NOR2_X1 U700 ( .A1(A[0]), .A2(n1), .ZN(ab_0__23_) );
  NOR2_X1 U701 ( .A1(n15), .A2(n51), .ZN(ab_0__22_) );
  NOR2_X1 U702 ( .A1(n16), .A2(n51), .ZN(ab_0__21_) );
  NOR2_X1 U703 ( .A1(n17), .A2(n51), .ZN(ab_0__20_) );
  NOR2_X1 U704 ( .A1(n19), .A2(n51), .ZN(ab_0__19_) );
  NOR2_X1 U705 ( .A1(n20), .A2(n51), .ZN(ab_0__18_) );
  NOR2_X1 U706 ( .A1(n21), .A2(n51), .ZN(ab_0__17_) );
  NOR2_X1 U707 ( .A1(n22), .A2(n51), .ZN(ab_0__16_) );
  NOR2_X1 U708 ( .A1(n23), .A2(n51), .ZN(ab_0__15_) );
  NOR2_X1 U709 ( .A1(n24), .A2(n51), .ZN(ab_0__14_) );
  NOR2_X1 U710 ( .A1(n25), .A2(n51), .ZN(ab_0__13_) );
  NOR2_X1 U711 ( .A1(n26), .A2(n51), .ZN(ab_0__12_) );
  NOR2_X1 U712 ( .A1(n27), .A2(n51), .ZN(ab_0__11_) );
  NOR2_X1 U713 ( .A1(n28), .A2(n51), .ZN(ab_0__10_) );
  INV_X1 U714 ( .A(B[23]), .ZN(QB) );
  INV_X1 U715 ( .A(A[23]), .ZN(QA) );
  AND3_X1 U716 ( .A1(ab_1__1_), .A2(B[0]), .A3(A[0]), .ZN(CARRYB_1__0_) );
  NOR2_X1 U717 ( .A1(n40), .A2(n18), .ZN(ab_1__1_) );
  INV_X1 U719 ( .A(CARRYB_23__23_), .ZN(A1_45_) );
endmodule


module iir_filter_DW01_add_6 ( A, B, CI, SUM, CO );
  input [45:0] A;
  input [45:0] B;
  output [45:0] SUM;
  input CI;
  output CO;
  wire   A_21_, A_20_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112;
  assign SUM[21] = A_21_;
  assign A_21_ = A[21];
  assign SUM[20] = A_20_;
  assign A_20_ = A[20];

  XOR2_X1 U2 ( .A(n1), .B(n2), .Z(SUM[45]) );
  XOR2_X1 U3 ( .A(B[45]), .B(A[45]), .Z(n2) );
  OAI21_X1 U4 ( .B1(n3), .B2(n4), .A(n5), .ZN(n1) );
  OAI21_X1 U5 ( .B1(A[44]), .B2(n6), .A(B[44]), .ZN(n5) );
  INV_X1 U6 ( .A(n3), .ZN(n6) );
  INV_X1 U7 ( .A(A[44]), .ZN(n4) );
  AOI21_X1 U8 ( .B1(A[43]), .B2(B[43]), .A(n7), .ZN(n3) );
  INV_X1 U9 ( .A(n8), .ZN(n7) );
  OAI22_X1 U10 ( .A1(n9), .A2(n10), .B1(A[43]), .B2(B[43]), .ZN(n8) );
  AOI21_X1 U11 ( .B1(n11), .B2(n12), .A(n13), .ZN(n9) );
  NAND3_X1 U12 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n12) );
  AOI21_X1 U13 ( .B1(n17), .B2(n16), .A(n18), .ZN(n11) );
  INV_X1 U14 ( .A(n19), .ZN(n18) );
  XOR2_X1 U15 ( .A(n20), .B(n21), .Z(SUM[42]) );
  NOR2_X1 U16 ( .A1(n10), .A2(n13), .ZN(n21) );
  NOR2_X1 U17 ( .A1(B[42]), .A2(A[42]), .ZN(n13) );
  AND2_X1 U18 ( .A1(B[42]), .A2(A[42]), .ZN(n10) );
  OAI21_X1 U19 ( .B1(n22), .B2(n23), .A(n19), .ZN(n20) );
  XOR2_X1 U20 ( .A(n24), .B(n23), .Z(SUM[41]) );
  AOI21_X1 U21 ( .B1(n15), .B2(n14), .A(n17), .ZN(n23) );
  INV_X1 U22 ( .A(n25), .ZN(n15) );
  NAND2_X1 U23 ( .A1(n16), .A2(n19), .ZN(n24) );
  NAND2_X1 U24 ( .A1(B[41]), .A2(A[41]), .ZN(n19) );
  INV_X1 U25 ( .A(n22), .ZN(n16) );
  NOR2_X1 U26 ( .A1(B[41]), .A2(A[41]), .ZN(n22) );
  XOR2_X1 U27 ( .A(n14), .B(n26), .Z(SUM[40]) );
  NOR2_X1 U28 ( .A1(n17), .A2(n25), .ZN(n26) );
  NOR2_X1 U29 ( .A1(B[40]), .A2(A[40]), .ZN(n25) );
  AND2_X1 U30 ( .A1(B[40]), .A2(A[40]), .ZN(n17) );
  OAI21_X1 U31 ( .B1(n27), .B2(n28), .A(n29), .ZN(n14) );
  XOR2_X1 U32 ( .A(n30), .B(n28), .Z(SUM[39]) );
  AOI21_X1 U33 ( .B1(n31), .B2(n32), .A(n33), .ZN(n28) );
  INV_X1 U34 ( .A(n34), .ZN(n31) );
  NAND2_X1 U35 ( .A1(n35), .A2(n29), .ZN(n30) );
  NAND2_X1 U36 ( .A1(B[39]), .A2(A[39]), .ZN(n29) );
  INV_X1 U37 ( .A(n27), .ZN(n35) );
  NOR2_X1 U38 ( .A1(B[39]), .A2(A[39]), .ZN(n27) );
  XOR2_X1 U39 ( .A(n32), .B(n36), .Z(SUM[38]) );
  NOR2_X1 U40 ( .A1(n33), .A2(n34), .ZN(n36) );
  NOR2_X1 U41 ( .A1(B[38]), .A2(A[38]), .ZN(n34) );
  AND2_X1 U42 ( .A1(B[38]), .A2(A[38]), .ZN(n33) );
  OAI21_X1 U43 ( .B1(n37), .B2(n38), .A(n39), .ZN(n32) );
  XOR2_X1 U44 ( .A(n40), .B(n38), .Z(SUM[37]) );
  AOI21_X1 U45 ( .B1(n41), .B2(n42), .A(n43), .ZN(n38) );
  INV_X1 U46 ( .A(n44), .ZN(n41) );
  NAND2_X1 U47 ( .A1(n45), .A2(n39), .ZN(n40) );
  NAND2_X1 U48 ( .A1(B[37]), .A2(A[37]), .ZN(n39) );
  INV_X1 U49 ( .A(n37), .ZN(n45) );
  NOR2_X1 U50 ( .A1(B[37]), .A2(A[37]), .ZN(n37) );
  XOR2_X1 U51 ( .A(n42), .B(n46), .Z(SUM[36]) );
  NOR2_X1 U52 ( .A1(n43), .A2(n44), .ZN(n46) );
  NOR2_X1 U53 ( .A1(B[36]), .A2(A[36]), .ZN(n44) );
  AND2_X1 U54 ( .A1(B[36]), .A2(A[36]), .ZN(n43) );
  OAI21_X1 U55 ( .B1(n47), .B2(n48), .A(n49), .ZN(n42) );
  XOR2_X1 U56 ( .A(n50), .B(n48), .Z(SUM[35]) );
  AOI21_X1 U57 ( .B1(n51), .B2(n52), .A(n53), .ZN(n48) );
  INV_X1 U58 ( .A(n54), .ZN(n51) );
  NAND2_X1 U59 ( .A1(n55), .A2(n49), .ZN(n50) );
  NAND2_X1 U60 ( .A1(B[35]), .A2(A[35]), .ZN(n49) );
  INV_X1 U61 ( .A(n47), .ZN(n55) );
  NOR2_X1 U62 ( .A1(B[35]), .A2(A[35]), .ZN(n47) );
  XOR2_X1 U63 ( .A(n52), .B(n56), .Z(SUM[34]) );
  NOR2_X1 U64 ( .A1(n53), .A2(n54), .ZN(n56) );
  NOR2_X1 U65 ( .A1(B[34]), .A2(A[34]), .ZN(n54) );
  AND2_X1 U66 ( .A1(B[34]), .A2(A[34]), .ZN(n53) );
  OAI21_X1 U67 ( .B1(n57), .B2(n58), .A(n59), .ZN(n52) );
  XOR2_X1 U68 ( .A(n60), .B(n58), .Z(SUM[33]) );
  AOI21_X1 U69 ( .B1(n61), .B2(n62), .A(n63), .ZN(n58) );
  INV_X1 U70 ( .A(n64), .ZN(n61) );
  NAND2_X1 U71 ( .A1(n65), .A2(n59), .ZN(n60) );
  NAND2_X1 U72 ( .A1(B[33]), .A2(A[33]), .ZN(n59) );
  INV_X1 U73 ( .A(n57), .ZN(n65) );
  NOR2_X1 U74 ( .A1(B[33]), .A2(A[33]), .ZN(n57) );
  XOR2_X1 U75 ( .A(n62), .B(n66), .Z(SUM[32]) );
  NOR2_X1 U76 ( .A1(n63), .A2(n64), .ZN(n66) );
  NOR2_X1 U77 ( .A1(B[32]), .A2(A[32]), .ZN(n64) );
  AND2_X1 U78 ( .A1(B[32]), .A2(A[32]), .ZN(n63) );
  OAI21_X1 U79 ( .B1(n67), .B2(n68), .A(n69), .ZN(n62) );
  XOR2_X1 U80 ( .A(n70), .B(n68), .Z(SUM[31]) );
  AOI21_X1 U81 ( .B1(n71), .B2(n72), .A(n73), .ZN(n68) );
  INV_X1 U82 ( .A(n74), .ZN(n71) );
  NAND2_X1 U83 ( .A1(n75), .A2(n69), .ZN(n70) );
  NAND2_X1 U84 ( .A1(B[31]), .A2(A[31]), .ZN(n69) );
  INV_X1 U85 ( .A(n67), .ZN(n75) );
  NOR2_X1 U86 ( .A1(B[31]), .A2(A[31]), .ZN(n67) );
  XOR2_X1 U87 ( .A(n72), .B(n76), .Z(SUM[30]) );
  NOR2_X1 U88 ( .A1(n73), .A2(n74), .ZN(n76) );
  NOR2_X1 U89 ( .A1(B[30]), .A2(A[30]), .ZN(n74) );
  AND2_X1 U90 ( .A1(B[30]), .A2(A[30]), .ZN(n73) );
  OAI21_X1 U91 ( .B1(n77), .B2(n78), .A(n79), .ZN(n72) );
  XOR2_X1 U92 ( .A(n80), .B(n78), .Z(SUM[29]) );
  AOI21_X1 U93 ( .B1(n81), .B2(n82), .A(n83), .ZN(n78) );
  INV_X1 U94 ( .A(n84), .ZN(n81) );
  NAND2_X1 U95 ( .A1(n85), .A2(n79), .ZN(n80) );
  NAND2_X1 U96 ( .A1(B[29]), .A2(A[29]), .ZN(n79) );
  INV_X1 U97 ( .A(n77), .ZN(n85) );
  NOR2_X1 U98 ( .A1(B[29]), .A2(A[29]), .ZN(n77) );
  XOR2_X1 U99 ( .A(n82), .B(n86), .Z(SUM[28]) );
  NOR2_X1 U100 ( .A1(n83), .A2(n84), .ZN(n86) );
  NOR2_X1 U101 ( .A1(B[28]), .A2(A[28]), .ZN(n84) );
  AND2_X1 U102 ( .A1(B[28]), .A2(A[28]), .ZN(n83) );
  OAI21_X1 U103 ( .B1(n87), .B2(n88), .A(n89), .ZN(n82) );
  XOR2_X1 U104 ( .A(n90), .B(n88), .Z(SUM[27]) );
  AOI21_X1 U105 ( .B1(n91), .B2(n92), .A(n93), .ZN(n88) );
  INV_X1 U106 ( .A(n94), .ZN(n92) );
  NAND2_X1 U107 ( .A1(n95), .A2(n89), .ZN(n90) );
  NAND2_X1 U108 ( .A1(B[27]), .A2(A[27]), .ZN(n89) );
  INV_X1 U109 ( .A(n87), .ZN(n95) );
  NOR2_X1 U110 ( .A1(B[27]), .A2(A[27]), .ZN(n87) );
  XOR2_X1 U111 ( .A(n91), .B(n96), .Z(SUM[26]) );
  NOR2_X1 U112 ( .A1(n93), .A2(n94), .ZN(n96) );
  NOR2_X1 U113 ( .A1(B[26]), .A2(A[26]), .ZN(n94) );
  AND2_X1 U114 ( .A1(B[26]), .A2(A[26]), .ZN(n93) );
  OAI21_X1 U115 ( .B1(n97), .B2(n98), .A(n99), .ZN(n91) );
  XOR2_X1 U116 ( .A(n100), .B(n98), .Z(SUM[25]) );
  AOI21_X1 U117 ( .B1(n101), .B2(n102), .A(n103), .ZN(n98) );
  INV_X1 U118 ( .A(n104), .ZN(n101) );
  NAND2_X1 U119 ( .A1(n105), .A2(n99), .ZN(n100) );
  NAND2_X1 U120 ( .A1(B[25]), .A2(A[25]), .ZN(n99) );
  INV_X1 U121 ( .A(n97), .ZN(n105) );
  NOR2_X1 U122 ( .A1(B[25]), .A2(A[25]), .ZN(n97) );
  XOR2_X1 U123 ( .A(n102), .B(n106), .Z(SUM[24]) );
  NOR2_X1 U124 ( .A1(n103), .A2(n104), .ZN(n106) );
  NOR2_X1 U125 ( .A1(B[24]), .A2(A[24]), .ZN(n104) );
  AND2_X1 U126 ( .A1(B[24]), .A2(A[24]), .ZN(n103) );
  OAI21_X1 U127 ( .B1(n107), .B2(n108), .A(n109), .ZN(n102) );
  XOR2_X1 U128 ( .A(n108), .B(n110), .Z(SUM[23]) );
  NAND2_X1 U129 ( .A1(n111), .A2(n109), .ZN(n110) );
  NAND2_X1 U130 ( .A1(B[23]), .A2(A[23]), .ZN(n109) );
  INV_X1 U131 ( .A(n107), .ZN(n111) );
  NOR2_X1 U132 ( .A1(B[23]), .A2(A[23]), .ZN(n107) );
  INV_X1 U133 ( .A(n112), .ZN(SUM[22]) );
  OAI21_X1 U134 ( .B1(B[22]), .B2(A[22]), .A(n108), .ZN(n112) );
  NAND2_X1 U135 ( .A1(B[22]), .A2(A[22]), .ZN(n108) );
endmodule


module iir_filter_DW02_mult_2 ( A, B, TC, PRODUCT );
  input [23:0] A;
  input [23:0] B;
  output [47:0] PRODUCT;
  input TC;
  wire   ab_23__23_, ab_23__22_, ab_23__21_, ab_23__20_, ab_23__19_,
         ab_23__18_, ab_23__17_, ab_23__16_, ab_23__15_, ab_23__14_,
         ab_23__13_, ab_23__12_, ab_23__11_, ab_23__10_, ab_23__9_, ab_23__8_,
         ab_23__7_, ab_23__6_, ab_23__5_, ab_23__4_, ab_23__3_, ab_23__2_,
         ab_23__1_, ab_23__0_, ab_22__23_, ab_22__22_, ab_22__21_, ab_22__20_,
         ab_22__19_, ab_22__18_, ab_22__17_, ab_22__16_, ab_22__15_,
         ab_22__14_, ab_22__13_, ab_22__12_, ab_22__11_, ab_22__10_, ab_22__9_,
         ab_22__8_, ab_22__7_, ab_22__6_, ab_22__5_, ab_22__4_, ab_22__3_,
         ab_22__2_, ab_22__1_, ab_22__0_, ab_21__23_, ab_21__22_, ab_21__21_,
         ab_21__20_, ab_21__19_, ab_21__18_, ab_21__17_, ab_21__16_,
         ab_21__15_, ab_21__14_, ab_21__13_, ab_21__12_, ab_21__11_,
         ab_21__10_, ab_21__9_, ab_21__8_, ab_21__7_, ab_21__6_, ab_21__5_,
         ab_21__4_, ab_21__3_, ab_21__2_, ab_21__1_, ab_21__0_, ab_20__23_,
         ab_20__22_, ab_20__21_, ab_20__20_, ab_20__19_, ab_20__18_,
         ab_20__17_, ab_20__16_, ab_20__15_, ab_20__14_, ab_20__13_,
         ab_20__12_, ab_20__11_, ab_20__10_, ab_20__9_, ab_20__8_, ab_20__7_,
         ab_20__6_, ab_20__5_, ab_20__4_, ab_20__3_, ab_20__2_, ab_20__1_,
         ab_20__0_, ab_19__23_, ab_19__22_, ab_19__21_, ab_19__20_, ab_19__19_,
         ab_19__18_, ab_19__17_, ab_19__16_, ab_19__15_, ab_19__14_,
         ab_19__13_, ab_19__12_, ab_19__11_, ab_19__10_, ab_19__9_, ab_19__8_,
         ab_19__7_, ab_19__6_, ab_19__5_, ab_19__4_, ab_19__3_, ab_19__2_,
         ab_19__1_, ab_19__0_, ab_18__23_, ab_18__22_, ab_18__21_, ab_18__20_,
         ab_18__19_, ab_18__18_, ab_18__17_, ab_18__16_, ab_18__15_,
         ab_18__14_, ab_18__13_, ab_18__12_, ab_18__11_, ab_18__10_, ab_18__9_,
         ab_18__8_, ab_18__7_, ab_18__6_, ab_18__5_, ab_18__4_, ab_18__3_,
         ab_18__2_, ab_18__1_, ab_18__0_, ab_17__23_, ab_17__22_, ab_17__21_,
         ab_17__20_, ab_17__19_, ab_17__18_, ab_17__17_, ab_17__16_,
         ab_17__15_, ab_17__14_, ab_17__13_, ab_17__12_, ab_17__11_,
         ab_17__10_, ab_17__9_, ab_17__8_, ab_17__7_, ab_17__6_, ab_17__5_,
         ab_17__4_, ab_17__3_, ab_17__2_, ab_17__1_, ab_17__0_, ab_16__23_,
         ab_16__22_, ab_16__21_, ab_16__20_, ab_16__19_, ab_16__18_,
         ab_16__17_, ab_16__16_, ab_16__15_, ab_16__14_, ab_16__13_,
         ab_16__12_, ab_16__11_, ab_16__10_, ab_16__9_, ab_16__8_, ab_16__7_,
         ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_, ab_16__1_,
         ab_16__0_, ab_15__23_, ab_15__22_, ab_15__21_, ab_15__20_, ab_15__19_,
         ab_15__18_, ab_15__17_, ab_15__16_, ab_15__15_, ab_15__14_,
         ab_15__13_, ab_15__12_, ab_15__11_, ab_15__10_, ab_15__9_, ab_15__8_,
         ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_, ab_15__3_, ab_15__2_,
         ab_15__1_, ab_15__0_, ab_14__23_, ab_14__22_, ab_14__21_, ab_14__20_,
         ab_14__19_, ab_14__18_, ab_14__17_, ab_14__16_, ab_14__15_,
         ab_14__14_, ab_14__13_, ab_14__12_, ab_14__11_, ab_14__10_, ab_14__9_,
         ab_14__8_, ab_14__7_, ab_14__6_, ab_14__5_, ab_14__4_, ab_14__3_,
         ab_14__2_, ab_14__1_, ab_14__0_, ab_13__23_, ab_13__22_, ab_13__21_,
         ab_13__20_, ab_13__19_, ab_13__18_, ab_13__17_, ab_13__16_,
         ab_13__15_, ab_13__14_, ab_13__13_, ab_13__12_, ab_13__11_,
         ab_13__10_, ab_13__9_, ab_13__8_, ab_13__7_, ab_13__6_, ab_13__5_,
         ab_13__4_, ab_13__3_, ab_13__2_, ab_13__1_, ab_13__0_, ab_12__23_,
         ab_12__22_, ab_12__21_, ab_12__20_, ab_12__19_, ab_12__18_,
         ab_12__17_, ab_12__16_, ab_12__15_, ab_12__14_, ab_12__13_,
         ab_12__12_, ab_12__11_, ab_12__10_, ab_12__9_, ab_12__8_, ab_12__7_,
         ab_12__6_, ab_12__5_, ab_12__4_, ab_12__3_, ab_12__2_, ab_12__1_,
         ab_12__0_, ab_11__23_, ab_11__22_, ab_11__21_, ab_11__20_, ab_11__19_,
         ab_11__18_, ab_11__17_, ab_11__16_, ab_11__15_, ab_11__14_,
         ab_11__13_, ab_11__12_, ab_11__11_, ab_11__10_, ab_11__9_, ab_11__8_,
         ab_11__7_, ab_11__6_, ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_,
         ab_11__1_, ab_11__0_, ab_10__23_, ab_10__22_, ab_10__21_, ab_10__20_,
         ab_10__19_, ab_10__18_, ab_10__17_, ab_10__16_, ab_10__15_,
         ab_10__14_, ab_10__13_, ab_10__12_, ab_10__11_, ab_10__10_, ab_10__9_,
         ab_10__8_, ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_,
         ab_10__2_, ab_10__1_, ab_10__0_, ab_9__23_, ab_9__22_, ab_9__21_,
         ab_9__20_, ab_9__19_, ab_9__18_, ab_9__17_, ab_9__16_, ab_9__15_,
         ab_9__14_, ab_9__13_, ab_9__12_, ab_9__11_, ab_9__10_, ab_9__9_,
         ab_9__8_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_,
         ab_9__1_, ab_9__0_, ab_8__23_, ab_8__22_, ab_8__21_, ab_8__20_,
         ab_8__19_, ab_8__18_, ab_8__17_, ab_8__16_, ab_8__15_, ab_8__14_,
         ab_8__13_, ab_8__12_, ab_8__11_, ab_8__10_, ab_8__9_, ab_8__8_,
         ab_8__7_, ab_8__6_, ab_8__5_, ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_,
         ab_8__0_, ab_7__23_, ab_7__22_, ab_7__21_, ab_7__20_, ab_7__19_,
         ab_7__18_, ab_7__17_, ab_7__16_, ab_7__15_, ab_7__14_, ab_7__13_,
         ab_7__12_, ab_7__11_, ab_7__10_, ab_7__9_, ab_7__8_, ab_7__7_,
         ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_,
         ab_6__23_, ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_, ab_6__18_,
         ab_6__17_, ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_, ab_6__12_,
         ab_6__11_, ab_6__10_, ab_6__9_, ab_6__8_, ab_6__7_, ab_6__6_,
         ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_, ab_5__23_,
         ab_5__22_, ab_5__21_, ab_5__20_, ab_5__19_, ab_5__18_, ab_5__17_,
         ab_5__16_, ab_5__15_, ab_5__14_, ab_5__13_, ab_5__12_, ab_5__11_,
         ab_5__10_, ab_5__9_, ab_5__8_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_,
         ab_5__3_, ab_5__2_, ab_5__1_, ab_5__0_, ab_4__23_, ab_4__22_,
         ab_4__21_, ab_4__20_, ab_4__19_, ab_4__18_, ab_4__17_, ab_4__16_,
         ab_4__15_, ab_4__14_, ab_4__13_, ab_4__12_, ab_4__11_, ab_4__10_,
         ab_4__9_, ab_4__8_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_,
         ab_4__2_, ab_4__1_, ab_4__0_, ab_3__23_, ab_3__22_, ab_3__21_,
         ab_3__20_, ab_3__19_, ab_3__18_, ab_3__17_, ab_3__16_, ab_3__15_,
         ab_3__14_, ab_3__13_, ab_3__12_, ab_3__11_, ab_3__10_, ab_3__9_,
         ab_3__8_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_, ab_3__2_,
         ab_3__1_, ab_3__0_, ab_2__23_, ab_2__22_, ab_2__21_, ab_2__20_,
         ab_2__19_, ab_2__18_, ab_2__17_, ab_2__16_, ab_2__15_, ab_2__14_,
         ab_2__13_, ab_2__12_, ab_2__11_, ab_2__10_, ab_2__9_, ab_2__8_,
         ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_,
         ab_2__0_, ab_1__23_, ab_1__22_, ab_1__21_, ab_1__20_, ab_1__19_,
         ab_1__18_, ab_1__17_, ab_1__16_, ab_1__15_, ab_1__14_, ab_1__13_,
         ab_1__12_, ab_1__11_, ab_1__10_, ab_1__9_, ab_1__8_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_0__23_,
         ab_0__22_, ab_0__21_, ab_0__20_, ab_0__19_, ab_0__18_, ab_0__17_,
         ab_0__16_, ab_0__15_, ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_,
         ab_0__10_, ab_0__9_, ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_23__23_, CARRYB_23__22_, CARRYB_23__21_,
         CARRYB_23__20_, CARRYB_23__19_, CARRYB_23__18_, CARRYB_23__17_,
         CARRYB_23__16_, CARRYB_23__15_, CARRYB_23__14_, CARRYB_23__13_,
         CARRYB_23__12_, CARRYB_23__11_, CARRYB_23__10_, CARRYB_23__9_,
         CARRYB_23__8_, CARRYB_23__7_, CARRYB_23__6_, CARRYB_23__5_,
         CARRYB_23__4_, CARRYB_23__3_, CARRYB_23__2_, CARRYB_23__1_,
         CARRYB_23__0_, CARRYB_22__22_, CARRYB_22__21_, CARRYB_22__20_,
         CARRYB_22__19_, CARRYB_22__18_, CARRYB_22__17_, CARRYB_22__16_,
         CARRYB_22__15_, CARRYB_22__14_, CARRYB_22__13_, CARRYB_22__12_,
         CARRYB_22__11_, CARRYB_22__10_, CARRYB_22__9_, CARRYB_22__8_,
         CARRYB_22__7_, CARRYB_22__6_, CARRYB_22__5_, CARRYB_22__4_,
         CARRYB_22__3_, CARRYB_22__2_, CARRYB_22__1_, CARRYB_22__0_,
         CARRYB_21__22_, CARRYB_21__21_, CARRYB_21__20_, CARRYB_21__19_,
         CARRYB_21__18_, CARRYB_21__17_, CARRYB_21__16_, CARRYB_21__15_,
         CARRYB_21__14_, CARRYB_21__13_, CARRYB_21__12_, CARRYB_21__11_,
         CARRYB_21__10_, CARRYB_21__9_, CARRYB_21__8_, CARRYB_21__7_,
         CARRYB_21__6_, CARRYB_21__5_, CARRYB_21__4_, CARRYB_21__3_,
         CARRYB_21__2_, CARRYB_21__1_, CARRYB_21__0_, CARRYB_20__22_,
         CARRYB_20__21_, CARRYB_20__20_, CARRYB_20__19_, CARRYB_20__18_,
         CARRYB_20__17_, CARRYB_20__16_, CARRYB_20__15_, CARRYB_20__14_,
         CARRYB_20__13_, CARRYB_20__12_, CARRYB_20__11_, CARRYB_20__10_,
         CARRYB_20__9_, CARRYB_20__8_, CARRYB_20__7_, CARRYB_20__6_,
         CARRYB_20__5_, CARRYB_20__4_, CARRYB_20__3_, CARRYB_20__2_,
         CARRYB_20__1_, CARRYB_20__0_, CARRYB_19__22_, CARRYB_19__21_,
         CARRYB_19__20_, CARRYB_19__19_, CARRYB_19__18_, CARRYB_19__17_,
         CARRYB_19__16_, CARRYB_19__15_, CARRYB_19__14_, CARRYB_19__13_,
         CARRYB_19__12_, CARRYB_19__11_, CARRYB_19__10_, CARRYB_19__9_,
         CARRYB_19__8_, CARRYB_19__7_, CARRYB_19__6_, CARRYB_19__5_,
         CARRYB_19__4_, CARRYB_19__3_, CARRYB_19__2_, CARRYB_19__1_,
         CARRYB_19__0_, CARRYB_18__22_, CARRYB_18__21_, CARRYB_18__20_,
         CARRYB_18__19_, CARRYB_18__18_, CARRYB_18__17_, CARRYB_18__16_,
         CARRYB_18__15_, CARRYB_18__14_, CARRYB_18__13_, CARRYB_18__12_,
         CARRYB_18__11_, CARRYB_18__10_, CARRYB_18__9_, CARRYB_18__8_,
         CARRYB_18__7_, CARRYB_18__6_, CARRYB_18__5_, CARRYB_18__4_,
         CARRYB_18__3_, CARRYB_18__2_, CARRYB_18__1_, CARRYB_18__0_,
         CARRYB_17__22_, CARRYB_17__21_, CARRYB_17__20_, CARRYB_17__19_,
         CARRYB_17__18_, CARRYB_17__17_, CARRYB_17__16_, CARRYB_17__15_,
         CARRYB_17__14_, CARRYB_17__13_, CARRYB_17__12_, CARRYB_17__11_,
         CARRYB_17__10_, CARRYB_17__9_, CARRYB_17__8_, CARRYB_17__7_,
         CARRYB_17__6_, CARRYB_17__5_, CARRYB_17__4_, CARRYB_17__3_,
         CARRYB_17__2_, CARRYB_17__1_, CARRYB_17__0_, CARRYB_16__22_,
         CARRYB_16__21_, CARRYB_16__20_, CARRYB_16__19_, CARRYB_16__18_,
         CARRYB_16__17_, CARRYB_16__16_, CARRYB_16__15_, CARRYB_16__14_,
         CARRYB_16__13_, CARRYB_16__12_, CARRYB_16__11_, CARRYB_16__10_,
         CARRYB_16__9_, CARRYB_16__8_, CARRYB_16__7_, CARRYB_16__6_,
         CARRYB_16__5_, CARRYB_16__4_, CARRYB_16__3_, CARRYB_16__2_,
         CARRYB_16__1_, CARRYB_16__0_, CARRYB_15__22_, CARRYB_15__21_,
         CARRYB_15__20_, CARRYB_15__19_, CARRYB_15__18_, CARRYB_15__17_,
         CARRYB_15__16_, CARRYB_15__15_, CARRYB_15__14_, CARRYB_15__13_,
         CARRYB_15__12_, CARRYB_15__11_, CARRYB_15__10_, CARRYB_15__9_,
         CARRYB_15__8_, CARRYB_15__7_, CARRYB_15__6_, CARRYB_15__5_,
         CARRYB_15__4_, CARRYB_15__3_, CARRYB_15__2_, CARRYB_15__1_,
         CARRYB_15__0_, CARRYB_14__22_, CARRYB_14__21_, CARRYB_14__20_,
         CARRYB_14__19_, CARRYB_14__18_, CARRYB_14__17_, CARRYB_14__16_,
         CARRYB_14__15_, CARRYB_14__14_, CARRYB_14__13_, CARRYB_14__12_,
         CARRYB_14__11_, CARRYB_14__10_, CARRYB_14__9_, CARRYB_14__8_,
         CARRYB_14__7_, CARRYB_14__6_, CARRYB_14__5_, CARRYB_14__4_,
         CARRYB_14__3_, CARRYB_14__2_, CARRYB_14__1_, CARRYB_14__0_,
         CARRYB_13__22_, CARRYB_13__21_, CARRYB_13__20_, CARRYB_13__19_,
         CARRYB_13__18_, CARRYB_13__17_, CARRYB_13__16_, CARRYB_13__15_,
         CARRYB_13__14_, CARRYB_13__13_, CARRYB_13__12_, CARRYB_13__11_,
         CARRYB_13__10_, CARRYB_13__9_, CARRYB_13__8_, CARRYB_13__7_,
         CARRYB_13__6_, CARRYB_13__5_, CARRYB_13__4_, CARRYB_13__3_,
         CARRYB_13__2_, CARRYB_13__1_, CARRYB_13__0_, CARRYB_12__22_,
         CARRYB_12__21_, CARRYB_12__20_, CARRYB_12__19_, CARRYB_12__18_,
         CARRYB_12__17_, CARRYB_12__16_, CARRYB_12__15_, CARRYB_12__14_,
         CARRYB_12__13_, CARRYB_12__12_, CARRYB_12__11_, CARRYB_12__10_,
         CARRYB_12__9_, CARRYB_12__8_, CARRYB_12__7_, CARRYB_12__6_,
         CARRYB_12__5_, CARRYB_12__4_, CARRYB_12__3_, CARRYB_12__2_,
         CARRYB_12__1_, CARRYB_12__0_, CARRYB_11__22_, CARRYB_11__21_,
         CARRYB_11__20_, CARRYB_11__19_, CARRYB_11__18_, CARRYB_11__17_,
         CARRYB_11__16_, CARRYB_11__15_, CARRYB_11__14_, CARRYB_11__13_,
         CARRYB_11__12_, CARRYB_11__11_, CARRYB_11__10_, CARRYB_11__9_,
         CARRYB_11__8_, CARRYB_11__7_, CARRYB_11__6_, CARRYB_11__5_,
         CARRYB_11__4_, CARRYB_11__3_, CARRYB_11__2_, CARRYB_11__1_,
         CARRYB_11__0_, CARRYB_10__22_, CARRYB_10__21_, CARRYB_10__20_,
         CARRYB_10__19_, CARRYB_10__18_, CARRYB_10__17_, CARRYB_10__16_,
         CARRYB_10__15_, CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_,
         CARRYB_10__11_, CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_,
         CARRYB_10__7_, CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_,
         CARRYB_10__3_, CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_,
         CARRYB_9__22_, CARRYB_9__21_, CARRYB_9__20_, CARRYB_9__19_,
         CARRYB_9__18_, CARRYB_9__17_, CARRYB_9__16_, CARRYB_9__15_,
         CARRYB_9__14_, CARRYB_9__13_, CARRYB_9__12_, CARRYB_9__11_,
         CARRYB_9__10_, CARRYB_9__9_, CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_,
         CARRYB_9__5_, CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_,
         CARRYB_9__0_, CARRYB_8__22_, CARRYB_8__21_, CARRYB_8__20_,
         CARRYB_8__19_, CARRYB_8__18_, CARRYB_8__17_, CARRYB_8__16_,
         CARRYB_8__15_, CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_,
         CARRYB_8__11_, CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_,
         CARRYB_8__7_, CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_,
         CARRYB_8__2_, CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__22_,
         CARRYB_7__21_, CARRYB_7__20_, CARRYB_7__19_, CARRYB_7__18_,
         CARRYB_7__17_, CARRYB_7__16_, CARRYB_7__15_, CARRYB_7__14_,
         CARRYB_7__13_, CARRYB_7__12_, CARRYB_7__11_, CARRYB_7__10_,
         CARRYB_7__9_, CARRYB_7__8_, CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_,
         CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_,
         CARRYB_6__22_, CARRYB_6__21_, CARRYB_6__20_, CARRYB_6__19_,
         CARRYB_6__18_, CARRYB_6__17_, CARRYB_6__16_, CARRYB_6__15_,
         CARRYB_6__14_, CARRYB_6__13_, CARRYB_6__12_, CARRYB_6__11_,
         CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_, CARRYB_6__7_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__22_, CARRYB_5__21_, CARRYB_5__20_,
         CARRYB_5__19_, CARRYB_5__18_, CARRYB_5__17_, CARRYB_5__16_,
         CARRYB_5__15_, CARRYB_5__14_, CARRYB_5__13_, CARRYB_5__12_,
         CARRYB_5__11_, CARRYB_5__10_, CARRYB_5__9_, CARRYB_5__8_,
         CARRYB_5__7_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__22_,
         CARRYB_4__21_, CARRYB_4__20_, CARRYB_4__19_, CARRYB_4__18_,
         CARRYB_4__17_, CARRYB_4__16_, CARRYB_4__15_, CARRYB_4__14_,
         CARRYB_4__13_, CARRYB_4__12_, CARRYB_4__11_, CARRYB_4__10_,
         CARRYB_4__9_, CARRYB_4__8_, CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__22_, CARRYB_3__21_, CARRYB_3__20_, CARRYB_3__19_,
         CARRYB_3__18_, CARRYB_3__17_, CARRYB_3__16_, CARRYB_3__15_,
         CARRYB_3__14_, CARRYB_3__13_, CARRYB_3__12_, CARRYB_3__11_,
         CARRYB_3__10_, CARRYB_3__9_, CARRYB_3__8_, CARRYB_3__7_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__22_, CARRYB_2__21_, CARRYB_2__20_,
         CARRYB_2__19_, CARRYB_2__18_, CARRYB_2__17_, CARRYB_2__16_,
         CARRYB_2__15_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__22_,
         CARRYB_1__21_, CARRYB_1__20_, CARRYB_1__19_, CARRYB_1__18_,
         CARRYB_1__17_, CARRYB_1__16_, CARRYB_1__15_, CARRYB_1__14_,
         CARRYB_1__13_, CARRYB_1__12_, CARRYB_1__11_, CARRYB_1__10_,
         CARRYB_1__9_, CARRYB_1__8_, CARRYB_1__7_, CARRYB_1__6_, CARRYB_1__5_,
         CARRYB_1__4_, CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_,
         SUMB_23__23_, SUMB_23__22_, SUMB_23__21_, SUMB_23__20_, SUMB_23__19_,
         SUMB_23__18_, SUMB_23__17_, SUMB_23__16_, SUMB_23__15_, SUMB_23__14_,
         SUMB_23__13_, SUMB_23__12_, SUMB_23__11_, SUMB_23__10_, SUMB_23__9_,
         SUMB_23__8_, SUMB_23__7_, SUMB_23__6_, SUMB_23__5_, SUMB_23__4_,
         SUMB_23__3_, SUMB_23__2_, SUMB_23__1_, SUMB_23__0_, SUMB_22__22_,
         SUMB_22__21_, SUMB_22__20_, SUMB_22__19_, SUMB_22__18_, SUMB_22__17_,
         SUMB_22__16_, SUMB_22__15_, SUMB_22__14_, SUMB_22__13_, SUMB_22__12_,
         SUMB_22__11_, SUMB_22__10_, SUMB_22__9_, SUMB_22__8_, SUMB_22__7_,
         SUMB_22__6_, SUMB_22__5_, SUMB_22__4_, SUMB_22__3_, SUMB_22__2_,
         SUMB_22__1_, SUMB_21__22_, SUMB_21__21_, SUMB_21__20_, SUMB_21__19_,
         SUMB_21__18_, SUMB_21__17_, SUMB_21__16_, SUMB_21__15_, SUMB_21__14_,
         SUMB_21__13_, SUMB_21__12_, SUMB_21__11_, SUMB_21__10_, SUMB_21__9_,
         SUMB_21__8_, SUMB_21__7_, SUMB_21__6_, SUMB_21__5_, SUMB_21__4_,
         SUMB_21__3_, SUMB_21__2_, SUMB_21__1_, SUMB_20__22_, SUMB_20__21_,
         SUMB_20__20_, SUMB_20__19_, SUMB_20__18_, SUMB_20__17_, SUMB_20__16_,
         SUMB_20__15_, SUMB_20__14_, SUMB_20__13_, SUMB_20__12_, SUMB_20__11_,
         SUMB_20__10_, SUMB_20__9_, SUMB_20__8_, SUMB_20__7_, SUMB_20__6_,
         SUMB_20__5_, SUMB_20__4_, SUMB_20__3_, SUMB_20__2_, SUMB_20__1_,
         SUMB_19__22_, SUMB_19__21_, SUMB_19__20_, SUMB_19__19_, SUMB_19__18_,
         SUMB_19__17_, SUMB_19__16_, SUMB_19__15_, SUMB_19__14_, SUMB_19__13_,
         SUMB_19__12_, SUMB_19__11_, SUMB_19__10_, SUMB_19__9_, SUMB_19__8_,
         SUMB_19__7_, SUMB_19__6_, SUMB_19__5_, SUMB_19__4_, SUMB_19__3_,
         SUMB_19__2_, SUMB_19__1_, SUMB_18__22_, SUMB_18__21_, SUMB_18__20_,
         SUMB_18__19_, SUMB_18__18_, SUMB_18__17_, SUMB_18__16_, SUMB_18__15_,
         SUMB_18__14_, SUMB_18__13_, SUMB_18__12_, SUMB_18__11_, SUMB_18__10_,
         SUMB_18__9_, SUMB_18__8_, SUMB_18__7_, SUMB_18__6_, SUMB_18__5_,
         SUMB_18__4_, SUMB_18__3_, SUMB_18__2_, SUMB_18__1_, SUMB_17__22_,
         SUMB_17__21_, SUMB_17__20_, SUMB_17__19_, SUMB_17__18_, SUMB_17__17_,
         SUMB_17__16_, SUMB_17__15_, SUMB_17__14_, SUMB_17__13_, SUMB_17__12_,
         SUMB_17__11_, SUMB_17__10_, SUMB_17__9_, SUMB_17__8_, SUMB_17__7_,
         SUMB_17__6_, SUMB_17__5_, SUMB_17__4_, SUMB_17__3_, SUMB_17__2_,
         SUMB_17__1_, SUMB_16__22_, SUMB_16__21_, SUMB_16__20_, SUMB_16__19_,
         SUMB_16__18_, SUMB_16__17_, SUMB_16__16_, SUMB_16__15_, SUMB_16__14_,
         SUMB_16__13_, SUMB_16__12_, SUMB_16__11_, SUMB_16__10_, SUMB_16__9_,
         SUMB_16__8_, SUMB_16__7_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_,
         SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, SUMB_15__22_, SUMB_15__21_,
         SUMB_15__20_, SUMB_15__19_, SUMB_15__18_, SUMB_15__17_, SUMB_15__16_,
         SUMB_15__15_, SUMB_15__14_, SUMB_15__13_, SUMB_15__12_, SUMB_15__11_,
         SUMB_15__10_, SUMB_15__9_, SUMB_15__8_, SUMB_15__7_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_14__22_, SUMB_14__21_, SUMB_14__20_, SUMB_14__19_, SUMB_14__18_,
         SUMB_14__17_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_, SUMB_14__13_,
         SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_, SUMB_14__8_,
         SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_,
         SUMB_14__2_, SUMB_14__1_, SUMB_13__22_, SUMB_13__21_, SUMB_13__20_,
         SUMB_13__19_, SUMB_13__18_, SUMB_13__17_, SUMB_13__16_, SUMB_13__15_,
         SUMB_13__14_, SUMB_13__13_, SUMB_13__12_, SUMB_13__11_, SUMB_13__10_,
         SUMB_13__9_, SUMB_13__8_, SUMB_13__7_, SUMB_13__6_, SUMB_13__5_,
         SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_, SUMB_12__22_,
         SUMB_12__21_, SUMB_12__20_, SUMB_12__19_, SUMB_12__18_, SUMB_12__17_,
         SUMB_12__16_, SUMB_12__15_, SUMB_12__14_, SUMB_12__13_, SUMB_12__12_,
         SUMB_12__11_, SUMB_12__10_, SUMB_12__9_, SUMB_12__8_, SUMB_12__7_,
         SUMB_12__6_, SUMB_12__5_, SUMB_12__4_, SUMB_12__3_, SUMB_12__2_,
         SUMB_12__1_, SUMB_11__22_, SUMB_11__21_, SUMB_11__20_, SUMB_11__19_,
         SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_, SUMB_11__14_,
         SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_, SUMB_11__9_,
         SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_, SUMB_11__4_,
         SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__22_, SUMB_10__21_,
         SUMB_10__20_, SUMB_10__19_, SUMB_10__18_, SUMB_10__17_, SUMB_10__16_,
         SUMB_10__15_, SUMB_10__14_, SUMB_10__13_, SUMB_10__12_, SUMB_10__11_,
         SUMB_10__10_, SUMB_10__9_, SUMB_10__8_, SUMB_10__7_, SUMB_10__6_,
         SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_,
         SUMB_9__22_, SUMB_9__21_, SUMB_9__20_, SUMB_9__19_, SUMB_9__18_,
         SUMB_9__17_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_, SUMB_9__13_,
         SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_, SUMB_9__8_,
         SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_,
         SUMB_9__2_, SUMB_9__1_, SUMB_8__22_, SUMB_8__21_, SUMB_8__20_,
         SUMB_8__19_, SUMB_8__18_, SUMB_8__17_, SUMB_8__16_, SUMB_8__15_,
         SUMB_8__14_, SUMB_8__13_, SUMB_8__12_, SUMB_8__11_, SUMB_8__10_,
         SUMB_8__9_, SUMB_8__8_, SUMB_8__7_, SUMB_8__6_, SUMB_8__5_,
         SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_, SUMB_7__22_,
         SUMB_7__21_, SUMB_7__20_, SUMB_7__19_, SUMB_7__18_, SUMB_7__17_,
         SUMB_7__16_, SUMB_7__15_, SUMB_7__14_, SUMB_7__13_, SUMB_7__12_,
         SUMB_7__11_, SUMB_7__10_, SUMB_7__9_, SUMB_7__8_, SUMB_7__7_,
         SUMB_7__6_, SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_,
         SUMB_7__1_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_, SUMB_6__19_,
         SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_, SUMB_6__14_,
         SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_, SUMB_6__9_,
         SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_,
         SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__22_, SUMB_5__21_,
         SUMB_5__20_, SUMB_5__19_, SUMB_5__18_, SUMB_5__17_, SUMB_5__16_,
         SUMB_5__15_, SUMB_5__14_, SUMB_5__13_, SUMB_5__12_, SUMB_5__11_,
         SUMB_5__10_, SUMB_5__9_, SUMB_5__8_, SUMB_5__7_, SUMB_5__6_,
         SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_,
         SUMB_4__22_, SUMB_4__21_, SUMB_4__20_, SUMB_4__19_, SUMB_4__18_,
         SUMB_4__17_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_, SUMB_4__13_,
         SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_, SUMB_4__8_,
         SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_,
         SUMB_4__2_, SUMB_4__1_, SUMB_3__22_, SUMB_3__21_, SUMB_3__20_,
         SUMB_3__19_, SUMB_3__18_, SUMB_3__17_, SUMB_3__16_, SUMB_3__15_,
         SUMB_3__14_, SUMB_3__13_, SUMB_3__12_, SUMB_3__11_, SUMB_3__10_,
         SUMB_3__9_, SUMB_3__8_, SUMB_3__7_, SUMB_3__6_, SUMB_3__5_,
         SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_, SUMB_2__22_,
         SUMB_2__21_, SUMB_2__20_, SUMB_2__19_, SUMB_2__18_, SUMB_2__17_,
         SUMB_2__16_, SUMB_2__15_, SUMB_2__14_, SUMB_2__13_, SUMB_2__12_,
         SUMB_2__11_, SUMB_2__10_, SUMB_2__9_, SUMB_2__8_, SUMB_2__7_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__22_, SUMB_1__21_, SUMB_1__20_, SUMB_1__19_,
         SUMB_1__18_, SUMB_1__17_, SUMB_1__16_, SUMB_1__15_, SUMB_1__14_,
         SUMB_1__13_, SUMB_1__12_, SUMB_1__11_, SUMB_1__10_, SUMB_1__9_,
         SUMB_1__8_, SUMB_1__7_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_,
         SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, QA, QB, A1_45_, A1_44_, A1_43_,
         A1_42_, A1_41_, A1_40_, A1_39_, A1_38_, A1_37_, A1_36_, A1_35_,
         A1_34_, A1_33_, A1_32_, A1_31_, A1_30_, A1_29_, A1_28_, A1_27_,
         A1_26_, A1_25_, A1_24_, A1_23_, A1_22_, A1_21_, A1_20_, A1_19_,
         A1_18_, A1_17_, A1_16_, A1_15_, A1_14_, A1_13_, A1_12_, A1_11_,
         A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_,
         A1_0_, A2_45_, A2_44_, A2_43_, A2_42_, A2_41_, A2_40_, A2_39_, A2_38_,
         A2_37_, A2_36_, A2_35_, A2_34_, A2_33_, A2_32_, A2_31_, A2_30_,
         A2_29_, A2_28_, A2_27_, A2_26_, A2_25_, A2_24_, A2_23_, A2_22_, n1,
         n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21;

  FA_X1 S14_23_0 ( .A(A[23]), .B(B[23]), .CI(SUMB_23__0_), .CO(A2_22_), .S(
        A1_21_) );
  FA_X1 S4_0 ( .A(ab_23__0_), .B(CARRYB_22__0_), .CI(SUMB_22__1_), .CO(
        CARRYB_23__0_), .S(SUMB_23__0_) );
  FA_X1 S4_1 ( .A(ab_23__1_), .B(CARRYB_22__1_), .CI(SUMB_22__2_), .CO(
        CARRYB_23__1_), .S(SUMB_23__1_) );
  FA_X1 S4_2 ( .A(ab_23__2_), .B(CARRYB_22__2_), .CI(SUMB_22__3_), .CO(
        CARRYB_23__2_), .S(SUMB_23__2_) );
  FA_X1 S4_3 ( .A(ab_23__3_), .B(CARRYB_22__3_), .CI(SUMB_22__4_), .CO(
        CARRYB_23__3_), .S(SUMB_23__3_) );
  FA_X1 S4_4 ( .A(ab_23__4_), .B(CARRYB_22__4_), .CI(SUMB_22__5_), .CO(
        CARRYB_23__4_), .S(SUMB_23__4_) );
  FA_X1 S4_5 ( .A(ab_23__5_), .B(CARRYB_22__5_), .CI(SUMB_22__6_), .CO(
        CARRYB_23__5_), .S(SUMB_23__5_) );
  FA_X1 S4_6 ( .A(ab_23__6_), .B(CARRYB_22__6_), .CI(SUMB_22__7_), .CO(
        CARRYB_23__6_), .S(SUMB_23__6_) );
  FA_X1 S4_7 ( .A(ab_23__7_), .B(CARRYB_22__7_), .CI(SUMB_22__8_), .CO(
        CARRYB_23__7_), .S(SUMB_23__7_) );
  FA_X1 S4_8 ( .A(ab_23__8_), .B(CARRYB_22__8_), .CI(SUMB_22__9_), .CO(
        CARRYB_23__8_), .S(SUMB_23__8_) );
  FA_X1 S4_9 ( .A(ab_23__9_), .B(CARRYB_22__9_), .CI(SUMB_22__10_), .CO(
        CARRYB_23__9_), .S(SUMB_23__9_) );
  FA_X1 S4_10 ( .A(ab_23__10_), .B(CARRYB_22__10_), .CI(SUMB_22__11_), .CO(
        CARRYB_23__10_), .S(SUMB_23__10_) );
  FA_X1 S4_11 ( .A(ab_23__11_), .B(CARRYB_22__11_), .CI(SUMB_22__12_), .CO(
        CARRYB_23__11_), .S(SUMB_23__11_) );
  FA_X1 S4_12 ( .A(ab_23__12_), .B(CARRYB_22__12_), .CI(SUMB_22__13_), .CO(
        CARRYB_23__12_), .S(SUMB_23__12_) );
  FA_X1 S4_13 ( .A(ab_23__13_), .B(CARRYB_22__13_), .CI(SUMB_22__14_), .CO(
        CARRYB_23__13_), .S(SUMB_23__13_) );
  FA_X1 S4_14 ( .A(ab_23__14_), .B(CARRYB_22__14_), .CI(SUMB_22__15_), .CO(
        CARRYB_23__14_), .S(SUMB_23__14_) );
  FA_X1 S4_15 ( .A(ab_23__15_), .B(CARRYB_22__15_), .CI(SUMB_22__16_), .CO(
        CARRYB_23__15_), .S(SUMB_23__15_) );
  FA_X1 S4_16 ( .A(ab_23__16_), .B(CARRYB_22__16_), .CI(SUMB_22__17_), .CO(
        CARRYB_23__16_), .S(SUMB_23__16_) );
  FA_X1 S4_17 ( .A(ab_23__17_), .B(CARRYB_22__17_), .CI(SUMB_22__18_), .CO(
        CARRYB_23__17_), .S(SUMB_23__17_) );
  FA_X1 S4_18 ( .A(ab_23__18_), .B(CARRYB_22__18_), .CI(SUMB_22__19_), .CO(
        CARRYB_23__18_), .S(SUMB_23__18_) );
  FA_X1 S4_19 ( .A(ab_23__19_), .B(CARRYB_22__19_), .CI(SUMB_22__20_), .CO(
        CARRYB_23__19_), .S(SUMB_23__19_) );
  FA_X1 S4_20 ( .A(ab_23__20_), .B(CARRYB_22__20_), .CI(SUMB_22__21_), .CO(
        CARRYB_23__20_), .S(SUMB_23__20_) );
  FA_X1 S4_21 ( .A(ab_23__21_), .B(CARRYB_22__21_), .CI(SUMB_22__22_), .CO(
        CARRYB_23__21_), .S(SUMB_23__21_) );
  FA_X1 S5_22 ( .A(ab_23__22_), .B(CARRYB_22__22_), .CI(ab_22__23_), .CO(
        CARRYB_23__22_), .S(SUMB_23__22_) );
  FA_X1 S14_23 ( .A(n3), .B(n1), .CI(ab_23__23_), .CO(CARRYB_23__23_), .S(
        SUMB_23__23_) );
  FA_X1 S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), .CO(
        CARRYB_22__0_), .S(A1_20_) );
  FA_X1 S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), .CO(
        CARRYB_22__1_), .S(SUMB_22__1_) );
  FA_X1 S2_22_2 ( .A(ab_22__2_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), .CO(
        CARRYB_22__2_), .S(SUMB_22__2_) );
  FA_X1 S2_22_3 ( .A(ab_22__3_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), .CO(
        CARRYB_22__3_), .S(SUMB_22__3_) );
  FA_X1 S2_22_4 ( .A(ab_22__4_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), .CO(
        CARRYB_22__4_), .S(SUMB_22__4_) );
  FA_X1 S2_22_5 ( .A(ab_22__5_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), .CO(
        CARRYB_22__5_), .S(SUMB_22__5_) );
  FA_X1 S2_22_6 ( .A(ab_22__6_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), .CO(
        CARRYB_22__6_), .S(SUMB_22__6_) );
  FA_X1 S2_22_7 ( .A(ab_22__7_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), .CO(
        CARRYB_22__7_), .S(SUMB_22__7_) );
  FA_X1 S2_22_8 ( .A(ab_22__8_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), .CO(
        CARRYB_22__8_), .S(SUMB_22__8_) );
  FA_X1 S2_22_9 ( .A(ab_22__9_), .B(CARRYB_21__9_), .CI(SUMB_21__10_), .CO(
        CARRYB_22__9_), .S(SUMB_22__9_) );
  FA_X1 S2_22_10 ( .A(ab_22__10_), .B(CARRYB_21__10_), .CI(SUMB_21__11_), .CO(
        CARRYB_22__10_), .S(SUMB_22__10_) );
  FA_X1 S2_22_11 ( .A(ab_22__11_), .B(CARRYB_21__11_), .CI(SUMB_21__12_), .CO(
        CARRYB_22__11_), .S(SUMB_22__11_) );
  FA_X1 S2_22_12 ( .A(ab_22__12_), .B(CARRYB_21__12_), .CI(SUMB_21__13_), .CO(
        CARRYB_22__12_), .S(SUMB_22__12_) );
  FA_X1 S2_22_13 ( .A(ab_22__13_), .B(CARRYB_21__13_), .CI(SUMB_21__14_), .CO(
        CARRYB_22__13_), .S(SUMB_22__13_) );
  FA_X1 S2_22_14 ( .A(ab_22__14_), .B(CARRYB_21__14_), .CI(SUMB_21__15_), .CO(
        CARRYB_22__14_), .S(SUMB_22__14_) );
  FA_X1 S2_22_15 ( .A(ab_22__15_), .B(CARRYB_21__15_), .CI(SUMB_21__16_), .CO(
        CARRYB_22__15_), .S(SUMB_22__15_) );
  FA_X1 S2_22_16 ( .A(ab_22__16_), .B(CARRYB_21__16_), .CI(SUMB_21__17_), .CO(
        CARRYB_22__16_), .S(SUMB_22__16_) );
  FA_X1 S2_22_17 ( .A(ab_22__17_), .B(CARRYB_21__17_), .CI(SUMB_21__18_), .CO(
        CARRYB_22__17_), .S(SUMB_22__17_) );
  FA_X1 S2_22_18 ( .A(ab_22__18_), .B(CARRYB_21__18_), .CI(SUMB_21__19_), .CO(
        CARRYB_22__18_), .S(SUMB_22__18_) );
  FA_X1 S2_22_19 ( .A(ab_22__19_), .B(CARRYB_21__19_), .CI(SUMB_21__20_), .CO(
        CARRYB_22__19_), .S(SUMB_22__19_) );
  FA_X1 S2_22_20 ( .A(ab_22__20_), .B(CARRYB_21__20_), .CI(SUMB_21__21_), .CO(
        CARRYB_22__20_), .S(SUMB_22__20_) );
  FA_X1 S2_22_21 ( .A(ab_22__21_), .B(CARRYB_21__21_), .CI(SUMB_21__22_), .CO(
        CARRYB_22__21_), .S(SUMB_22__21_) );
  FA_X1 S3_22_22 ( .A(ab_22__22_), .B(CARRYB_21__22_), .CI(ab_21__23_), .CO(
        CARRYB_22__22_), .S(SUMB_22__22_) );
  FA_X1 S1_21_0 ( .A(ab_21__0_), .B(CARRYB_20__0_), .CI(SUMB_20__1_), .CO(
        CARRYB_21__0_), .S(A1_19_) );
  FA_X1 S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), .CO(
        CARRYB_21__1_), .S(SUMB_21__1_) );
  FA_X1 S2_21_2 ( .A(ab_21__2_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), .CO(
        CARRYB_21__2_), .S(SUMB_21__2_) );
  FA_X1 S2_21_3 ( .A(ab_21__3_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), .CO(
        CARRYB_21__3_), .S(SUMB_21__3_) );
  FA_X1 S2_21_4 ( .A(ab_21__4_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), .CO(
        CARRYB_21__4_), .S(SUMB_21__4_) );
  FA_X1 S2_21_5 ( .A(ab_21__5_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), .CO(
        CARRYB_21__5_), .S(SUMB_21__5_) );
  FA_X1 S2_21_6 ( .A(ab_21__6_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), .CO(
        CARRYB_21__6_), .S(SUMB_21__6_) );
  FA_X1 S2_21_7 ( .A(ab_21__7_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), .CO(
        CARRYB_21__7_), .S(SUMB_21__7_) );
  FA_X1 S2_21_8 ( .A(ab_21__8_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), .CO(
        CARRYB_21__8_), .S(SUMB_21__8_) );
  FA_X1 S2_21_9 ( .A(ab_21__9_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), .CO(
        CARRYB_21__9_), .S(SUMB_21__9_) );
  FA_X1 S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .CI(SUMB_20__11_), .CO(
        CARRYB_21__10_), .S(SUMB_21__10_) );
  FA_X1 S2_21_11 ( .A(ab_21__11_), .B(CARRYB_20__11_), .CI(SUMB_20__12_), .CO(
        CARRYB_21__11_), .S(SUMB_21__11_) );
  FA_X1 S2_21_12 ( .A(ab_21__12_), .B(CARRYB_20__12_), .CI(SUMB_20__13_), .CO(
        CARRYB_21__12_), .S(SUMB_21__12_) );
  FA_X1 S2_21_13 ( .A(ab_21__13_), .B(CARRYB_20__13_), .CI(SUMB_20__14_), .CO(
        CARRYB_21__13_), .S(SUMB_21__13_) );
  FA_X1 S2_21_14 ( .A(ab_21__14_), .B(CARRYB_20__14_), .CI(SUMB_20__15_), .CO(
        CARRYB_21__14_), .S(SUMB_21__14_) );
  FA_X1 S2_21_15 ( .A(ab_21__15_), .B(CARRYB_20__15_), .CI(SUMB_20__16_), .CO(
        CARRYB_21__15_), .S(SUMB_21__15_) );
  FA_X1 S2_21_16 ( .A(ab_21__16_), .B(CARRYB_20__16_), .CI(SUMB_20__17_), .CO(
        CARRYB_21__16_), .S(SUMB_21__16_) );
  FA_X1 S2_21_17 ( .A(ab_21__17_), .B(CARRYB_20__17_), .CI(SUMB_20__18_), .CO(
        CARRYB_21__17_), .S(SUMB_21__17_) );
  FA_X1 S2_21_18 ( .A(ab_21__18_), .B(CARRYB_20__18_), .CI(SUMB_20__19_), .CO(
        CARRYB_21__18_), .S(SUMB_21__18_) );
  FA_X1 S2_21_19 ( .A(ab_21__19_), .B(CARRYB_20__19_), .CI(SUMB_20__20_), .CO(
        CARRYB_21__19_), .S(SUMB_21__19_) );
  FA_X1 S2_21_20 ( .A(ab_21__20_), .B(CARRYB_20__20_), .CI(SUMB_20__21_), .CO(
        CARRYB_21__20_), .S(SUMB_21__20_) );
  FA_X1 S2_21_21 ( .A(ab_21__21_), .B(CARRYB_20__21_), .CI(SUMB_20__22_), .CO(
        CARRYB_21__21_), .S(SUMB_21__21_) );
  FA_X1 S3_21_22 ( .A(ab_21__22_), .B(CARRYB_20__22_), .CI(ab_20__23_), .CO(
        CARRYB_21__22_), .S(SUMB_21__22_) );
  FA_X1 S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), .CO(
        CARRYB_20__0_), .S(A1_18_) );
  FA_X1 S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), .CO(
        CARRYB_20__1_), .S(SUMB_20__1_) );
  FA_X1 S2_20_2 ( .A(ab_20__2_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), .CO(
        CARRYB_20__2_), .S(SUMB_20__2_) );
  FA_X1 S2_20_3 ( .A(ab_20__3_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), .CO(
        CARRYB_20__3_), .S(SUMB_20__3_) );
  FA_X1 S2_20_4 ( .A(ab_20__4_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), .CO(
        CARRYB_20__4_), .S(SUMB_20__4_) );
  FA_X1 S2_20_5 ( .A(ab_20__5_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), .CO(
        CARRYB_20__5_), .S(SUMB_20__5_) );
  FA_X1 S2_20_6 ( .A(ab_20__6_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), .CO(
        CARRYB_20__6_), .S(SUMB_20__6_) );
  FA_X1 S2_20_7 ( .A(ab_20__7_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), .CO(
        CARRYB_20__7_), .S(SUMB_20__7_) );
  FA_X1 S2_20_8 ( .A(ab_20__8_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), .CO(
        CARRYB_20__8_), .S(SUMB_20__8_) );
  FA_X1 S2_20_9 ( .A(ab_20__9_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), .CO(
        CARRYB_20__9_), .S(SUMB_20__9_) );
  FA_X1 S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), .CO(
        CARRYB_20__10_), .S(SUMB_20__10_) );
  FA_X1 S2_20_11 ( .A(ab_20__11_), .B(CARRYB_19__11_), .CI(SUMB_19__12_), .CO(
        CARRYB_20__11_), .S(SUMB_20__11_) );
  FA_X1 S2_20_12 ( .A(ab_20__12_), .B(CARRYB_19__12_), .CI(SUMB_19__13_), .CO(
        CARRYB_20__12_), .S(SUMB_20__12_) );
  FA_X1 S2_20_13 ( .A(ab_20__13_), .B(CARRYB_19__13_), .CI(SUMB_19__14_), .CO(
        CARRYB_20__13_), .S(SUMB_20__13_) );
  FA_X1 S2_20_14 ( .A(ab_20__14_), .B(CARRYB_19__14_), .CI(SUMB_19__15_), .CO(
        CARRYB_20__14_), .S(SUMB_20__14_) );
  FA_X1 S2_20_15 ( .A(ab_20__15_), .B(CARRYB_19__15_), .CI(SUMB_19__16_), .CO(
        CARRYB_20__15_), .S(SUMB_20__15_) );
  FA_X1 S2_20_16 ( .A(ab_20__16_), .B(CARRYB_19__16_), .CI(SUMB_19__17_), .CO(
        CARRYB_20__16_), .S(SUMB_20__16_) );
  FA_X1 S2_20_17 ( .A(ab_20__17_), .B(CARRYB_19__17_), .CI(SUMB_19__18_), .CO(
        CARRYB_20__17_), .S(SUMB_20__17_) );
  FA_X1 S2_20_18 ( .A(ab_20__18_), .B(CARRYB_19__18_), .CI(SUMB_19__19_), .CO(
        CARRYB_20__18_), .S(SUMB_20__18_) );
  FA_X1 S2_20_19 ( .A(ab_20__19_), .B(CARRYB_19__19_), .CI(SUMB_19__20_), .CO(
        CARRYB_20__19_), .S(SUMB_20__19_) );
  FA_X1 S2_20_20 ( .A(ab_20__20_), .B(CARRYB_19__20_), .CI(SUMB_19__21_), .CO(
        CARRYB_20__20_), .S(SUMB_20__20_) );
  FA_X1 S2_20_21 ( .A(ab_20__21_), .B(CARRYB_19__21_), .CI(SUMB_19__22_), .CO(
        CARRYB_20__21_), .S(SUMB_20__21_) );
  FA_X1 S3_20_22 ( .A(ab_20__22_), .B(CARRYB_19__22_), .CI(ab_19__23_), .CO(
        CARRYB_20__22_), .S(SUMB_20__22_) );
  FA_X1 S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), .CO(
        CARRYB_19__0_), .S(A1_17_) );
  FA_X1 S2_19_1 ( .A(ab_19__1_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), .CO(
        CARRYB_19__1_), .S(SUMB_19__1_) );
  FA_X1 S2_19_2 ( .A(ab_19__2_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), .CO(
        CARRYB_19__2_), .S(SUMB_19__2_) );
  FA_X1 S2_19_3 ( .A(ab_19__3_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), .CO(
        CARRYB_19__3_), .S(SUMB_19__3_) );
  FA_X1 S2_19_4 ( .A(ab_19__4_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), .CO(
        CARRYB_19__4_), .S(SUMB_19__4_) );
  FA_X1 S2_19_5 ( .A(ab_19__5_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), .CO(
        CARRYB_19__5_), .S(SUMB_19__5_) );
  FA_X1 S2_19_6 ( .A(ab_19__6_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), .CO(
        CARRYB_19__6_), .S(SUMB_19__6_) );
  FA_X1 S2_19_7 ( .A(ab_19__7_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), .CO(
        CARRYB_19__7_), .S(SUMB_19__7_) );
  FA_X1 S2_19_8 ( .A(ab_19__8_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), .CO(
        CARRYB_19__8_), .S(SUMB_19__8_) );
  FA_X1 S2_19_9 ( .A(ab_19__9_), .B(CARRYB_18__9_), .CI(SUMB_18__10_), .CO(
        CARRYB_19__9_), .S(SUMB_19__9_) );
  FA_X1 S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), .CO(
        CARRYB_19__10_), .S(SUMB_19__10_) );
  FA_X1 S2_19_11 ( .A(ab_19__11_), .B(CARRYB_18__11_), .CI(SUMB_18__12_), .CO(
        CARRYB_19__11_), .S(SUMB_19__11_) );
  FA_X1 S2_19_12 ( .A(ab_19__12_), .B(CARRYB_18__12_), .CI(SUMB_18__13_), .CO(
        CARRYB_19__12_), .S(SUMB_19__12_) );
  FA_X1 S2_19_13 ( .A(ab_19__13_), .B(CARRYB_18__13_), .CI(SUMB_18__14_), .CO(
        CARRYB_19__13_), .S(SUMB_19__13_) );
  FA_X1 S2_19_14 ( .A(ab_19__14_), .B(CARRYB_18__14_), .CI(SUMB_18__15_), .CO(
        CARRYB_19__14_), .S(SUMB_19__14_) );
  FA_X1 S2_19_15 ( .A(ab_19__15_), .B(CARRYB_18__15_), .CI(SUMB_18__16_), .CO(
        CARRYB_19__15_), .S(SUMB_19__15_) );
  FA_X1 S2_19_16 ( .A(ab_19__16_), .B(CARRYB_18__16_), .CI(SUMB_18__17_), .CO(
        CARRYB_19__16_), .S(SUMB_19__16_) );
  FA_X1 S2_19_17 ( .A(ab_19__17_), .B(CARRYB_18__17_), .CI(SUMB_18__18_), .CO(
        CARRYB_19__17_), .S(SUMB_19__17_) );
  FA_X1 S2_19_18 ( .A(ab_19__18_), .B(CARRYB_18__18_), .CI(SUMB_18__19_), .CO(
        CARRYB_19__18_), .S(SUMB_19__18_) );
  FA_X1 S2_19_19 ( .A(ab_19__19_), .B(CARRYB_18__19_), .CI(SUMB_18__20_), .CO(
        CARRYB_19__19_), .S(SUMB_19__19_) );
  FA_X1 S2_19_20 ( .A(ab_19__20_), .B(CARRYB_18__20_), .CI(SUMB_18__21_), .CO(
        CARRYB_19__20_), .S(SUMB_19__20_) );
  FA_X1 S2_19_21 ( .A(ab_19__21_), .B(CARRYB_18__21_), .CI(SUMB_18__22_), .CO(
        CARRYB_19__21_), .S(SUMB_19__21_) );
  FA_X1 S3_19_22 ( .A(ab_19__22_), .B(CARRYB_18__22_), .CI(ab_18__23_), .CO(
        CARRYB_19__22_), .S(SUMB_19__22_) );
  FA_X1 S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), .CO(
        CARRYB_18__0_), .S(A1_16_) );
  FA_X1 S2_18_1 ( .A(ab_18__1_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), .CO(
        CARRYB_18__1_), .S(SUMB_18__1_) );
  FA_X1 S2_18_2 ( .A(ab_18__2_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), .CO(
        CARRYB_18__2_), .S(SUMB_18__2_) );
  FA_X1 S2_18_3 ( .A(ab_18__3_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), .CO(
        CARRYB_18__3_), .S(SUMB_18__3_) );
  FA_X1 S2_18_4 ( .A(ab_18__4_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), .CO(
        CARRYB_18__4_), .S(SUMB_18__4_) );
  FA_X1 S2_18_5 ( .A(ab_18__5_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), .CO(
        CARRYB_18__5_), .S(SUMB_18__5_) );
  FA_X1 S2_18_6 ( .A(ab_18__6_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), .CO(
        CARRYB_18__6_), .S(SUMB_18__6_) );
  FA_X1 S2_18_7 ( .A(ab_18__7_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), .CO(
        CARRYB_18__7_), .S(SUMB_18__7_) );
  FA_X1 S2_18_8 ( .A(ab_18__8_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), .CO(
        CARRYB_18__8_), .S(SUMB_18__8_) );
  FA_X1 S2_18_9 ( .A(ab_18__9_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), .CO(
        CARRYB_18__9_), .S(SUMB_18__9_) );
  FA_X1 S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), .CO(
        CARRYB_18__10_), .S(SUMB_18__10_) );
  FA_X1 S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), .CO(
        CARRYB_18__11_), .S(SUMB_18__11_) );
  FA_X1 S2_18_12 ( .A(ab_18__12_), .B(CARRYB_17__12_), .CI(SUMB_17__13_), .CO(
        CARRYB_18__12_), .S(SUMB_18__12_) );
  FA_X1 S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .CI(SUMB_17__14_), .CO(
        CARRYB_18__13_), .S(SUMB_18__13_) );
  FA_X1 S2_18_14 ( .A(ab_18__14_), .B(CARRYB_17__14_), .CI(SUMB_17__15_), .CO(
        CARRYB_18__14_), .S(SUMB_18__14_) );
  FA_X1 S2_18_15 ( .A(ab_18__15_), .B(CARRYB_17__15_), .CI(SUMB_17__16_), .CO(
        CARRYB_18__15_), .S(SUMB_18__15_) );
  FA_X1 S2_18_16 ( .A(ab_18__16_), .B(CARRYB_17__16_), .CI(SUMB_17__17_), .CO(
        CARRYB_18__16_), .S(SUMB_18__16_) );
  FA_X1 S2_18_17 ( .A(ab_18__17_), .B(CARRYB_17__17_), .CI(SUMB_17__18_), .CO(
        CARRYB_18__17_), .S(SUMB_18__17_) );
  FA_X1 S2_18_18 ( .A(ab_18__18_), .B(CARRYB_17__18_), .CI(SUMB_17__19_), .CO(
        CARRYB_18__18_), .S(SUMB_18__18_) );
  FA_X1 S2_18_19 ( .A(ab_18__19_), .B(CARRYB_17__19_), .CI(SUMB_17__20_), .CO(
        CARRYB_18__19_), .S(SUMB_18__19_) );
  FA_X1 S2_18_20 ( .A(ab_18__20_), .B(CARRYB_17__20_), .CI(SUMB_17__21_), .CO(
        CARRYB_18__20_), .S(SUMB_18__20_) );
  FA_X1 S2_18_21 ( .A(ab_18__21_), .B(CARRYB_17__21_), .CI(SUMB_17__22_), .CO(
        CARRYB_18__21_), .S(SUMB_18__21_) );
  FA_X1 S3_18_22 ( .A(ab_18__22_), .B(CARRYB_17__22_), .CI(ab_17__23_), .CO(
        CARRYB_18__22_), .S(SUMB_18__22_) );
  FA_X1 S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), .CO(
        CARRYB_17__0_), .S(A1_15_) );
  FA_X1 S2_17_1 ( .A(ab_17__1_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), .CO(
        CARRYB_17__1_), .S(SUMB_17__1_) );
  FA_X1 S2_17_2 ( .A(ab_17__2_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), .CO(
        CARRYB_17__2_), .S(SUMB_17__2_) );
  FA_X1 S2_17_3 ( .A(ab_17__3_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), .CO(
        CARRYB_17__3_), .S(SUMB_17__3_) );
  FA_X1 S2_17_4 ( .A(ab_17__4_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), .CO(
        CARRYB_17__4_), .S(SUMB_17__4_) );
  FA_X1 S2_17_5 ( .A(ab_17__5_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), .CO(
        CARRYB_17__5_), .S(SUMB_17__5_) );
  FA_X1 S2_17_6 ( .A(ab_17__6_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), .CO(
        CARRYB_17__6_), .S(SUMB_17__6_) );
  FA_X1 S2_17_7 ( .A(ab_17__7_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), .CO(
        CARRYB_17__7_), .S(SUMB_17__7_) );
  FA_X1 S2_17_8 ( .A(ab_17__8_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), .CO(
        CARRYB_17__8_), .S(SUMB_17__8_) );
  FA_X1 S2_17_9 ( .A(ab_17__9_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), .CO(
        CARRYB_17__9_), .S(SUMB_17__9_) );
  FA_X1 S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), .CO(
        CARRYB_17__10_), .S(SUMB_17__10_) );
  FA_X1 S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), .CO(
        CARRYB_17__11_), .S(SUMB_17__11_) );
  FA_X1 S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), .CO(
        CARRYB_17__12_), .S(SUMB_17__12_) );
  FA_X1 S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), .CO(
        CARRYB_17__13_), .S(SUMB_17__13_) );
  FA_X1 S2_17_14 ( .A(ab_17__14_), .B(CARRYB_16__14_), .CI(SUMB_16__15_), .CO(
        CARRYB_17__14_), .S(SUMB_17__14_) );
  FA_X1 S2_17_15 ( .A(ab_17__15_), .B(CARRYB_16__15_), .CI(SUMB_16__16_), .CO(
        CARRYB_17__15_), .S(SUMB_17__15_) );
  FA_X1 S2_17_16 ( .A(ab_17__16_), .B(CARRYB_16__16_), .CI(SUMB_16__17_), .CO(
        CARRYB_17__16_), .S(SUMB_17__16_) );
  FA_X1 S2_17_17 ( .A(ab_17__17_), .B(CARRYB_16__17_), .CI(SUMB_16__18_), .CO(
        CARRYB_17__17_), .S(SUMB_17__17_) );
  FA_X1 S2_17_18 ( .A(ab_17__18_), .B(CARRYB_16__18_), .CI(SUMB_16__19_), .CO(
        CARRYB_17__18_), .S(SUMB_17__18_) );
  FA_X1 S2_17_19 ( .A(ab_17__19_), .B(CARRYB_16__19_), .CI(SUMB_16__20_), .CO(
        CARRYB_17__19_), .S(SUMB_17__19_) );
  FA_X1 S2_17_20 ( .A(ab_17__20_), .B(CARRYB_16__20_), .CI(SUMB_16__21_), .CO(
        CARRYB_17__20_), .S(SUMB_17__20_) );
  FA_X1 S2_17_21 ( .A(ab_17__21_), .B(CARRYB_16__21_), .CI(SUMB_16__22_), .CO(
        CARRYB_17__21_), .S(SUMB_17__21_) );
  FA_X1 S3_17_22 ( .A(ab_17__22_), .B(CARRYB_16__22_), .CI(ab_16__23_), .CO(
        CARRYB_17__22_), .S(SUMB_17__22_) );
  FA_X1 S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(A1_14_) );
  FA_X1 S2_16_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  FA_X1 S2_16_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  FA_X1 S2_16_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  FA_X1 S2_16_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  FA_X1 S2_16_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  FA_X1 S2_16_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  FA_X1 S2_16_7 ( .A(ab_16__7_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), .CO(
        CARRYB_16__7_), .S(SUMB_16__7_) );
  FA_X1 S2_16_8 ( .A(ab_16__8_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), .CO(
        CARRYB_16__8_), .S(SUMB_16__8_) );
  FA_X1 S2_16_9 ( .A(ab_16__9_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), .CO(
        CARRYB_16__9_), .S(SUMB_16__9_) );
  FA_X1 S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), .CO(
        CARRYB_16__10_), .S(SUMB_16__10_) );
  FA_X1 S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), .CO(
        CARRYB_16__11_), .S(SUMB_16__11_) );
  FA_X1 S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), .CO(
        CARRYB_16__12_), .S(SUMB_16__12_) );
  FA_X1 S2_16_13 ( .A(ab_16__13_), .B(CARRYB_15__13_), .CI(SUMB_15__14_), .CO(
        CARRYB_16__13_), .S(SUMB_16__13_) );
  FA_X1 S2_16_14 ( .A(ab_16__14_), .B(CARRYB_15__14_), .CI(SUMB_15__15_), .CO(
        CARRYB_16__14_), .S(SUMB_16__14_) );
  FA_X1 S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .CI(SUMB_15__16_), .CO(
        CARRYB_16__15_), .S(SUMB_16__15_) );
  FA_X1 S2_16_16 ( .A(ab_16__16_), .B(CARRYB_15__16_), .CI(SUMB_15__17_), .CO(
        CARRYB_16__16_), .S(SUMB_16__16_) );
  FA_X1 S2_16_17 ( .A(ab_16__17_), .B(CARRYB_15__17_), .CI(SUMB_15__18_), .CO(
        CARRYB_16__17_), .S(SUMB_16__17_) );
  FA_X1 S2_16_18 ( .A(ab_16__18_), .B(CARRYB_15__18_), .CI(SUMB_15__19_), .CO(
        CARRYB_16__18_), .S(SUMB_16__18_) );
  FA_X1 S2_16_19 ( .A(ab_16__19_), .B(CARRYB_15__19_), .CI(SUMB_15__20_), .CO(
        CARRYB_16__19_), .S(SUMB_16__19_) );
  FA_X1 S2_16_20 ( .A(ab_16__20_), .B(CARRYB_15__20_), .CI(SUMB_15__21_), .CO(
        CARRYB_16__20_), .S(SUMB_16__20_) );
  FA_X1 S2_16_21 ( .A(ab_16__21_), .B(CARRYB_15__21_), .CI(SUMB_15__22_), .CO(
        CARRYB_16__21_), .S(SUMB_16__21_) );
  FA_X1 S3_16_22 ( .A(ab_16__22_), .B(CARRYB_15__22_), .CI(ab_15__23_), .CO(
        CARRYB_16__22_), .S(SUMB_16__22_) );
  FA_X1 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  FA_X1 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  FA_X1 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  FA_X1 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  FA_X1 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  FA_X1 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  FA_X1 S2_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  FA_X1 S2_15_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), .CO(
        CARRYB_15__7_), .S(SUMB_15__7_) );
  FA_X1 S2_15_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), .CO(
        CARRYB_15__8_), .S(SUMB_15__8_) );
  FA_X1 S2_15_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), .CO(
        CARRYB_15__9_), .S(SUMB_15__9_) );
  FA_X1 S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), .CO(
        CARRYB_15__10_), .S(SUMB_15__10_) );
  FA_X1 S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), .CO(
        CARRYB_15__11_), .S(SUMB_15__11_) );
  FA_X1 S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), .CO(
        CARRYB_15__12_), .S(SUMB_15__12_) );
  FA_X1 S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), .CO(
        CARRYB_15__13_), .S(SUMB_15__13_) );
  FA_X1 S2_15_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), .CO(
        CARRYB_15__14_), .S(SUMB_15__14_) );
  FA_X1 S2_15_15 ( .A(ab_15__15_), .B(CARRYB_14__15_), .CI(SUMB_14__16_), .CO(
        CARRYB_15__15_), .S(SUMB_15__15_) );
  FA_X1 S2_15_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .CI(SUMB_14__17_), .CO(
        CARRYB_15__16_), .S(SUMB_15__16_) );
  FA_X1 S2_15_17 ( .A(ab_15__17_), .B(CARRYB_14__17_), .CI(SUMB_14__18_), .CO(
        CARRYB_15__17_), .S(SUMB_15__17_) );
  FA_X1 S2_15_18 ( .A(ab_15__18_), .B(CARRYB_14__18_), .CI(SUMB_14__19_), .CO(
        CARRYB_15__18_), .S(SUMB_15__18_) );
  FA_X1 S2_15_19 ( .A(ab_15__19_), .B(CARRYB_14__19_), .CI(SUMB_14__20_), .CO(
        CARRYB_15__19_), .S(SUMB_15__19_) );
  FA_X1 S2_15_20 ( .A(ab_15__20_), .B(CARRYB_14__20_), .CI(SUMB_14__21_), .CO(
        CARRYB_15__20_), .S(SUMB_15__20_) );
  FA_X1 S2_15_21 ( .A(ab_15__21_), .B(CARRYB_14__21_), .CI(SUMB_14__22_), .CO(
        CARRYB_15__21_), .S(SUMB_15__21_) );
  FA_X1 S3_15_22 ( .A(ab_15__22_), .B(CARRYB_14__22_), .CI(ab_14__23_), .CO(
        CARRYB_15__22_), .S(SUMB_15__22_) );
  FA_X1 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  FA_X1 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  FA_X1 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  FA_X1 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  FA_X1 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  FA_X1 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  FA_X1 S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  FA_X1 S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), .CO(
        CARRYB_14__7_), .S(SUMB_14__7_) );
  FA_X1 S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), .CO(
        CARRYB_14__8_), .S(SUMB_14__8_) );
  FA_X1 S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), .CO(
        CARRYB_14__9_), .S(SUMB_14__9_) );
  FA_X1 S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), .CO(
        CARRYB_14__10_), .S(SUMB_14__10_) );
  FA_X1 S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), .CO(
        CARRYB_14__11_), .S(SUMB_14__11_) );
  FA_X1 S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), .CO(
        CARRYB_14__12_), .S(SUMB_14__12_) );
  FA_X1 S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), .CO(
        CARRYB_14__13_), .S(SUMB_14__13_) );
  FA_X1 S2_14_14 ( .A(ab_14__14_), .B(CARRYB_13__14_), .CI(SUMB_13__15_), .CO(
        CARRYB_14__14_), .S(SUMB_14__14_) );
  FA_X1 S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), .CO(
        CARRYB_14__15_), .S(SUMB_14__15_) );
  FA_X1 S2_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), .CO(
        CARRYB_14__16_), .S(SUMB_14__16_) );
  FA_X1 S2_14_17 ( .A(ab_14__17_), .B(CARRYB_13__17_), .CI(SUMB_13__18_), .CO(
        CARRYB_14__17_), .S(SUMB_14__17_) );
  FA_X1 S2_14_18 ( .A(ab_14__18_), .B(CARRYB_13__18_), .CI(SUMB_13__19_), .CO(
        CARRYB_14__18_), .S(SUMB_14__18_) );
  FA_X1 S2_14_19 ( .A(ab_14__19_), .B(CARRYB_13__19_), .CI(SUMB_13__20_), .CO(
        CARRYB_14__19_), .S(SUMB_14__19_) );
  FA_X1 S2_14_20 ( .A(ab_14__20_), .B(CARRYB_13__20_), .CI(SUMB_13__21_), .CO(
        CARRYB_14__20_), .S(SUMB_14__20_) );
  FA_X1 S2_14_21 ( .A(ab_14__21_), .B(CARRYB_13__21_), .CI(SUMB_13__22_), .CO(
        CARRYB_14__21_), .S(SUMB_14__21_) );
  FA_X1 S3_14_22 ( .A(ab_14__22_), .B(CARRYB_13__22_), .CI(ab_13__23_), .CO(
        CARRYB_14__22_), .S(SUMB_14__22_) );
  FA_X1 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  FA_X1 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  FA_X1 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  FA_X1 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  FA_X1 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  FA_X1 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  FA_X1 S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  FA_X1 S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), .CO(
        CARRYB_13__7_), .S(SUMB_13__7_) );
  FA_X1 S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), .CO(
        CARRYB_13__8_), .S(SUMB_13__8_) );
  FA_X1 S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), .CO(
        CARRYB_13__9_), .S(SUMB_13__9_) );
  FA_X1 S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), .CO(
        CARRYB_13__10_), .S(SUMB_13__10_) );
  FA_X1 S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), .CO(
        CARRYB_13__11_), .S(SUMB_13__11_) );
  FA_X1 S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), .CO(
        CARRYB_13__12_), .S(SUMB_13__12_) );
  FA_X1 S2_13_13 ( .A(ab_13__13_), .B(CARRYB_12__13_), .CI(SUMB_12__14_), .CO(
        CARRYB_13__13_), .S(SUMB_13__13_) );
  FA_X1 S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), .CO(
        CARRYB_13__14_), .S(SUMB_13__14_) );
  FA_X1 S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), .CO(
        CARRYB_13__15_), .S(SUMB_13__15_) );
  FA_X1 S2_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), .CO(
        CARRYB_13__16_), .S(SUMB_13__16_) );
  FA_X1 S2_13_17 ( .A(ab_13__17_), .B(CARRYB_12__17_), .CI(SUMB_12__18_), .CO(
        CARRYB_13__17_), .S(SUMB_13__17_) );
  FA_X1 S2_13_18 ( .A(ab_13__18_), .B(CARRYB_12__18_), .CI(SUMB_12__19_), .CO(
        CARRYB_13__18_), .S(SUMB_13__18_) );
  FA_X1 S2_13_19 ( .A(ab_13__19_), .B(CARRYB_12__19_), .CI(SUMB_12__20_), .CO(
        CARRYB_13__19_), .S(SUMB_13__19_) );
  FA_X1 S2_13_20 ( .A(ab_13__20_), .B(CARRYB_12__20_), .CI(SUMB_12__21_), .CO(
        CARRYB_13__20_), .S(SUMB_13__20_) );
  FA_X1 S2_13_21 ( .A(ab_13__21_), .B(CARRYB_12__21_), .CI(SUMB_12__22_), .CO(
        CARRYB_13__21_), .S(SUMB_13__21_) );
  FA_X1 S3_13_22 ( .A(ab_13__22_), .B(CARRYB_12__22_), .CI(ab_12__23_), .CO(
        CARRYB_13__22_), .S(SUMB_13__22_) );
  FA_X1 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  FA_X1 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  FA_X1 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  FA_X1 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  FA_X1 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  FA_X1 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  FA_X1 S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  FA_X1 S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), .CO(
        CARRYB_12__7_), .S(SUMB_12__7_) );
  FA_X1 S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), .CO(
        CARRYB_12__8_), .S(SUMB_12__8_) );
  FA_X1 S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), .CO(
        CARRYB_12__9_), .S(SUMB_12__9_) );
  FA_X1 S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), .CO(
        CARRYB_12__10_), .S(SUMB_12__10_) );
  FA_X1 S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), .CO(
        CARRYB_12__11_), .S(SUMB_12__11_) );
  FA_X1 S2_12_12 ( .A(ab_12__12_), .B(CARRYB_11__12_), .CI(SUMB_11__13_), .CO(
        CARRYB_12__12_), .S(SUMB_12__12_) );
  FA_X1 S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), .CO(
        CARRYB_12__13_), .S(SUMB_12__13_) );
  FA_X1 S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), .CO(
        CARRYB_12__14_), .S(SUMB_12__14_) );
  FA_X1 S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), .CO(
        CARRYB_12__15_), .S(SUMB_12__15_) );
  FA_X1 S2_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), .CO(
        CARRYB_12__16_), .S(SUMB_12__16_) );
  FA_X1 S2_12_17 ( .A(ab_12__17_), .B(CARRYB_11__17_), .CI(SUMB_11__18_), .CO(
        CARRYB_12__17_), .S(SUMB_12__17_) );
  FA_X1 S2_12_18 ( .A(ab_12__18_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), .CO(
        CARRYB_12__18_), .S(SUMB_12__18_) );
  FA_X1 S2_12_19 ( .A(ab_12__19_), .B(CARRYB_11__19_), .CI(SUMB_11__20_), .CO(
        CARRYB_12__19_), .S(SUMB_12__19_) );
  FA_X1 S2_12_20 ( .A(ab_12__20_), .B(CARRYB_11__20_), .CI(SUMB_11__21_), .CO(
        CARRYB_12__20_), .S(SUMB_12__20_) );
  FA_X1 S2_12_21 ( .A(ab_12__21_), .B(CARRYB_11__21_), .CI(SUMB_11__22_), .CO(
        CARRYB_12__21_), .S(SUMB_12__21_) );
  FA_X1 S3_12_22 ( .A(ab_12__22_), .B(CARRYB_11__22_), .CI(ab_11__23_), .CO(
        CARRYB_12__22_), .S(SUMB_12__22_) );
  FA_X1 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  FA_X1 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  FA_X1 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  FA_X1 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  FA_X1 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  FA_X1 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  FA_X1 S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  FA_X1 S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), .CO(
        CARRYB_11__7_), .S(SUMB_11__7_) );
  FA_X1 S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), .CO(
        CARRYB_11__8_), .S(SUMB_11__8_) );
  FA_X1 S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), .CO(
        CARRYB_11__9_), .S(SUMB_11__9_) );
  FA_X1 S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), .CO(
        CARRYB_11__10_), .S(SUMB_11__10_) );
  FA_X1 S2_11_11 ( .A(ab_11__11_), .B(CARRYB_10__11_), .CI(SUMB_10__12_), .CO(
        CARRYB_11__11_), .S(SUMB_11__11_) );
  FA_X1 S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), .CO(
        CARRYB_11__12_), .S(SUMB_11__12_) );
  FA_X1 S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), .CO(
        CARRYB_11__13_), .S(SUMB_11__13_) );
  FA_X1 S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), .CO(
        CARRYB_11__14_), .S(SUMB_11__14_) );
  FA_X1 S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), .CO(
        CARRYB_11__15_), .S(SUMB_11__15_) );
  FA_X1 S2_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(SUMB_10__17_), .CO(
        CARRYB_11__16_), .S(SUMB_11__16_) );
  FA_X1 S2_11_17 ( .A(ab_11__17_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), .CO(
        CARRYB_11__17_), .S(SUMB_11__17_) );
  FA_X1 S2_11_18 ( .A(ab_11__18_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), .CO(
        CARRYB_11__18_), .S(SUMB_11__18_) );
  FA_X1 S2_11_19 ( .A(ab_11__19_), .B(CARRYB_10__19_), .CI(SUMB_10__20_), .CO(
        CARRYB_11__19_), .S(SUMB_11__19_) );
  FA_X1 S2_11_20 ( .A(ab_11__20_), .B(CARRYB_10__20_), .CI(SUMB_10__21_), .CO(
        CARRYB_11__20_), .S(SUMB_11__20_) );
  FA_X1 S2_11_21 ( .A(ab_11__21_), .B(CARRYB_10__21_), .CI(SUMB_10__22_), .CO(
        CARRYB_11__21_), .S(SUMB_11__21_) );
  FA_X1 S3_11_22 ( .A(ab_11__22_), .B(CARRYB_10__22_), .CI(ab_10__23_), .CO(
        CARRYB_11__22_), .S(SUMB_11__22_) );
  FA_X1 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  FA_X1 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  FA_X1 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  FA_X1 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  FA_X1 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  FA_X1 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  FA_X1 S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  FA_X1 S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  FA_X1 S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  FA_X1 S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  FA_X1 S2_10_10 ( .A(ab_10__10_), .B(CARRYB_9__10_), .CI(SUMB_9__11_), .CO(
        CARRYB_10__10_), .S(SUMB_10__10_) );
  FA_X1 S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), .CO(
        CARRYB_10__11_), .S(SUMB_10__11_) );
  FA_X1 S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), .CO(
        CARRYB_10__12_), .S(SUMB_10__12_) );
  FA_X1 S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), .CO(
        CARRYB_10__13_), .S(SUMB_10__13_) );
  FA_X1 S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), .CO(
        CARRYB_10__14_), .S(SUMB_10__14_) );
  FA_X1 S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), .CO(
        CARRYB_10__15_), .S(SUMB_10__15_) );
  FA_X1 S2_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), .CO(
        CARRYB_10__16_), .S(SUMB_10__16_) );
  FA_X1 S2_10_17 ( .A(ab_10__17_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), .CO(
        CARRYB_10__17_), .S(SUMB_10__17_) );
  FA_X1 S2_10_18 ( .A(ab_10__18_), .B(CARRYB_9__18_), .CI(SUMB_9__19_), .CO(
        CARRYB_10__18_), .S(SUMB_10__18_) );
  FA_X1 S2_10_19 ( .A(ab_10__19_), .B(CARRYB_9__19_), .CI(SUMB_9__20_), .CO(
        CARRYB_10__19_), .S(SUMB_10__19_) );
  FA_X1 S2_10_20 ( .A(ab_10__20_), .B(CARRYB_9__20_), .CI(SUMB_9__21_), .CO(
        CARRYB_10__20_), .S(SUMB_10__20_) );
  FA_X1 S2_10_21 ( .A(ab_10__21_), .B(CARRYB_9__21_), .CI(SUMB_9__22_), .CO(
        CARRYB_10__21_), .S(SUMB_10__21_) );
  FA_X1 S3_10_22 ( .A(ab_10__22_), .B(CARRYB_9__22_), .CI(ab_9__23_), .CO(
        CARRYB_10__22_), .S(SUMB_10__22_) );
  FA_X1 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  FA_X1 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  FA_X1 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  FA_X1 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  FA_X1 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  FA_X1 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  FA_X1 S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  FA_X1 S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  FA_X1 S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  FA_X1 S2_9_9 ( .A(ab_9__9_), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  FA_X1 S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), .CO(
        CARRYB_9__10_), .S(SUMB_9__10_) );
  FA_X1 S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), .CO(
        CARRYB_9__11_), .S(SUMB_9__11_) );
  FA_X1 S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), .CO(
        CARRYB_9__12_), .S(SUMB_9__12_) );
  FA_X1 S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), .CO(
        CARRYB_9__13_), .S(SUMB_9__13_) );
  FA_X1 S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), .CO(
        CARRYB_9__14_), .S(SUMB_9__14_) );
  FA_X1 S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), .CO(
        CARRYB_9__15_), .S(SUMB_9__15_) );
  FA_X1 S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), .CO(
        CARRYB_9__16_), .S(SUMB_9__16_) );
  FA_X1 S2_9_17 ( .A(ab_9__17_), .B(CARRYB_8__17_), .CI(SUMB_8__18_), .CO(
        CARRYB_9__17_), .S(SUMB_9__17_) );
  FA_X1 S2_9_18 ( .A(ab_9__18_), .B(CARRYB_8__18_), .CI(SUMB_8__19_), .CO(
        CARRYB_9__18_), .S(SUMB_9__18_) );
  FA_X1 S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), .CO(
        CARRYB_9__19_), .S(SUMB_9__19_) );
  FA_X1 S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(SUMB_8__21_), .CO(
        CARRYB_9__20_), .S(SUMB_9__20_) );
  FA_X1 S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), .CO(
        CARRYB_9__21_), .S(SUMB_9__21_) );
  FA_X1 S3_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .CI(ab_8__23_), .CO(
        CARRYB_9__22_), .S(SUMB_9__22_) );
  FA_X1 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  FA_X1 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  FA_X1 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  FA_X1 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  FA_X1 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  FA_X1 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  FA_X1 S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  FA_X1 S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  FA_X1 S2_8_8 ( .A(ab_8__8_), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  FA_X1 S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  FA_X1 S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), .CO(
        CARRYB_8__10_), .S(SUMB_8__10_) );
  FA_X1 S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), .CO(
        CARRYB_8__11_), .S(SUMB_8__11_) );
  FA_X1 S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), .CO(
        CARRYB_8__12_), .S(SUMB_8__12_) );
  FA_X1 S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), .CO(
        CARRYB_8__13_), .S(SUMB_8__13_) );
  FA_X1 S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), .CO(
        CARRYB_8__14_), .S(SUMB_8__14_) );
  FA_X1 S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), .CO(
        CARRYB_8__15_), .S(SUMB_8__15_) );
  FA_X1 S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), .CO(
        CARRYB_8__16_), .S(SUMB_8__16_) );
  FA_X1 S2_8_17 ( .A(ab_8__17_), .B(CARRYB_7__17_), .CI(SUMB_7__18_), .CO(
        CARRYB_8__17_), .S(SUMB_8__17_) );
  FA_X1 S2_8_18 ( .A(ab_8__18_), .B(CARRYB_7__18_), .CI(SUMB_7__19_), .CO(
        CARRYB_8__18_), .S(SUMB_8__18_) );
  FA_X1 S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), .CO(
        CARRYB_8__19_), .S(SUMB_8__19_) );
  FA_X1 S2_8_20 ( .A(ab_8__20_), .B(CARRYB_7__20_), .CI(SUMB_7__21_), .CO(
        CARRYB_8__20_), .S(SUMB_8__20_) );
  FA_X1 S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), .CO(
        CARRYB_8__21_), .S(SUMB_8__21_) );
  FA_X1 S3_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(ab_7__23_), .CO(
        CARRYB_8__22_), .S(SUMB_8__22_) );
  FA_X1 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(A1_5_) );
  FA_X1 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S2_7_7 ( .A(ab_7__7_), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  FA_X1 S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  FA_X1 S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  FA_X1 S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), .CO(
        CARRYB_7__10_), .S(SUMB_7__10_) );
  FA_X1 S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), .CO(
        CARRYB_7__11_), .S(SUMB_7__11_) );
  FA_X1 S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), .CO(
        CARRYB_7__12_), .S(SUMB_7__12_) );
  FA_X1 S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), .CO(
        CARRYB_7__13_), .S(SUMB_7__13_) );
  FA_X1 S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), .CO(
        CARRYB_7__14_), .S(SUMB_7__14_) );
  FA_X1 S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), .CO(
        CARRYB_7__15_), .S(SUMB_7__15_) );
  FA_X1 S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), .CO(
        CARRYB_7__16_), .S(SUMB_7__16_) );
  FA_X1 S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), .CO(
        CARRYB_7__17_), .S(SUMB_7__17_) );
  FA_X1 S2_7_18 ( .A(ab_7__18_), .B(CARRYB_6__18_), .CI(SUMB_6__19_), .CO(
        CARRYB_7__18_), .S(SUMB_7__18_) );
  FA_X1 S2_7_19 ( .A(ab_7__19_), .B(CARRYB_6__19_), .CI(SUMB_6__20_), .CO(
        CARRYB_7__19_), .S(SUMB_7__19_) );
  FA_X1 S2_7_20 ( .A(ab_7__20_), .B(CARRYB_6__20_), .CI(SUMB_6__21_), .CO(
        CARRYB_7__20_), .S(SUMB_7__20_) );
  FA_X1 S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), .CO(
        CARRYB_7__21_), .S(SUMB_7__21_) );
  FA_X1 S3_7_22 ( .A(ab_7__22_), .B(CARRYB_6__22_), .CI(ab_6__23_), .CO(
        CARRYB_7__22_), .S(SUMB_7__22_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S2_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  FA_X1 S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  FA_X1 S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  FA_X1 S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), .CO(
        CARRYB_6__10_), .S(SUMB_6__10_) );
  FA_X1 S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), .CO(
        CARRYB_6__11_), .S(SUMB_6__11_) );
  FA_X1 S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), .CO(
        CARRYB_6__12_), .S(SUMB_6__12_) );
  FA_X1 S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), .CO(
        CARRYB_6__13_), .S(SUMB_6__13_) );
  FA_X1 S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), .CO(
        CARRYB_6__14_), .S(SUMB_6__14_) );
  FA_X1 S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), .CO(
        CARRYB_6__15_), .S(SUMB_6__15_) );
  FA_X1 S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), .CO(
        CARRYB_6__16_), .S(SUMB_6__16_) );
  FA_X1 S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), .CO(
        CARRYB_6__17_), .S(SUMB_6__17_) );
  FA_X1 S2_6_18 ( .A(ab_6__18_), .B(CARRYB_5__18_), .CI(SUMB_5__19_), .CO(
        CARRYB_6__18_), .S(SUMB_6__18_) );
  FA_X1 S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), .CO(
        CARRYB_6__19_), .S(SUMB_6__19_) );
  FA_X1 S2_6_20 ( .A(ab_6__20_), .B(CARRYB_5__20_), .CI(SUMB_5__21_), .CO(
        CARRYB_6__20_), .S(SUMB_6__20_) );
  FA_X1 S2_6_21 ( .A(ab_6__21_), .B(CARRYB_5__21_), .CI(SUMB_5__22_), .CO(
        CARRYB_6__21_), .S(SUMB_6__21_) );
  FA_X1 S3_6_22 ( .A(ab_6__22_), .B(CARRYB_5__22_), .CI(ab_5__23_), .CO(
        CARRYB_6__22_), .S(SUMB_6__22_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  FA_X1 S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  FA_X1 S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  FA_X1 S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), .CO(
        CARRYB_5__10_), .S(SUMB_5__10_) );
  FA_X1 S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), .CO(
        CARRYB_5__11_), .S(SUMB_5__11_) );
  FA_X1 S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), .CO(
        CARRYB_5__12_), .S(SUMB_5__12_) );
  FA_X1 S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), .CO(
        CARRYB_5__13_), .S(SUMB_5__13_) );
  FA_X1 S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), .CO(
        CARRYB_5__14_), .S(SUMB_5__14_) );
  FA_X1 S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), .CO(
        CARRYB_5__15_), .S(SUMB_5__15_) );
  FA_X1 S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), .CO(
        CARRYB_5__16_), .S(SUMB_5__16_) );
  FA_X1 S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), .CO(
        CARRYB_5__17_), .S(SUMB_5__17_) );
  FA_X1 S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), .CO(
        CARRYB_5__18_), .S(SUMB_5__18_) );
  FA_X1 S2_5_19 ( .A(ab_5__19_), .B(CARRYB_4__19_), .CI(SUMB_4__20_), .CO(
        CARRYB_5__19_), .S(SUMB_5__19_) );
  FA_X1 S2_5_20 ( .A(ab_5__20_), .B(CARRYB_4__20_), .CI(SUMB_4__21_), .CO(
        CARRYB_5__20_), .S(SUMB_5__20_) );
  FA_X1 S2_5_21 ( .A(ab_5__21_), .B(CARRYB_4__21_), .CI(SUMB_4__22_), .CO(
        CARRYB_5__21_), .S(SUMB_5__21_) );
  FA_X1 S3_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(ab_4__23_), .CO(
        CARRYB_5__22_), .S(SUMB_5__22_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  FA_X1 S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  FA_X1 S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  FA_X1 S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), .CO(
        CARRYB_4__10_), .S(SUMB_4__10_) );
  FA_X1 S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), .CO(
        CARRYB_4__11_), .S(SUMB_4__11_) );
  FA_X1 S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), .CO(
        CARRYB_4__12_), .S(SUMB_4__12_) );
  FA_X1 S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), .CO(
        CARRYB_4__13_), .S(SUMB_4__13_) );
  FA_X1 S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), .CO(
        CARRYB_4__14_), .S(SUMB_4__14_) );
  FA_X1 S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), .CO(
        CARRYB_4__15_), .S(SUMB_4__15_) );
  FA_X1 S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), .CO(
        CARRYB_4__16_), .S(SUMB_4__16_) );
  FA_X1 S2_4_17 ( .A(ab_4__17_), .B(CARRYB_3__17_), .CI(SUMB_3__18_), .CO(
        CARRYB_4__17_), .S(SUMB_4__17_) );
  FA_X1 S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), .CO(
        CARRYB_4__18_), .S(SUMB_4__18_) );
  FA_X1 S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), .CO(
        CARRYB_4__19_), .S(SUMB_4__19_) );
  FA_X1 S2_4_20 ( .A(ab_4__20_), .B(CARRYB_3__20_), .CI(SUMB_3__21_), .CO(
        CARRYB_4__20_), .S(SUMB_4__20_) );
  FA_X1 S2_4_21 ( .A(ab_4__21_), .B(CARRYB_3__21_), .CI(SUMB_3__22_), .CO(
        CARRYB_4__21_), .S(SUMB_4__21_) );
  FA_X1 S3_4_22 ( .A(ab_4__22_), .B(CARRYB_3__22_), .CI(ab_3__23_), .CO(
        CARRYB_4__22_), .S(SUMB_4__22_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  FA_X1 S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  FA_X1 S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  FA_X1 S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), .CO(
        CARRYB_3__10_), .S(SUMB_3__10_) );
  FA_X1 S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), .CO(
        CARRYB_3__11_), .S(SUMB_3__11_) );
  FA_X1 S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), .CO(
        CARRYB_3__12_), .S(SUMB_3__12_) );
  FA_X1 S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), .CO(
        CARRYB_3__13_), .S(SUMB_3__13_) );
  FA_X1 S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), .CO(
        CARRYB_3__14_), .S(SUMB_3__14_) );
  FA_X1 S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), .CO(
        CARRYB_3__15_), .S(SUMB_3__15_) );
  FA_X1 S2_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(SUMB_2__17_), .CO(
        CARRYB_3__16_), .S(SUMB_3__16_) );
  FA_X1 S2_3_17 ( .A(ab_3__17_), .B(CARRYB_2__17_), .CI(SUMB_2__18_), .CO(
        CARRYB_3__17_), .S(SUMB_3__17_) );
  FA_X1 S2_3_18 ( .A(ab_3__18_), .B(CARRYB_2__18_), .CI(SUMB_2__19_), .CO(
        CARRYB_3__18_), .S(SUMB_3__18_) );
  FA_X1 S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), .CO(
        CARRYB_3__19_), .S(SUMB_3__19_) );
  FA_X1 S2_3_20 ( .A(ab_3__20_), .B(CARRYB_2__20_), .CI(SUMB_2__21_), .CO(
        CARRYB_3__20_), .S(SUMB_3__20_) );
  FA_X1 S2_3_21 ( .A(ab_3__21_), .B(CARRYB_2__21_), .CI(SUMB_2__22_), .CO(
        CARRYB_3__21_), .S(SUMB_3__21_) );
  FA_X1 S3_3_22 ( .A(ab_3__22_), .B(CARRYB_2__22_), .CI(ab_2__23_), .CO(
        CARRYB_3__22_), .S(SUMB_3__22_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S2_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(SUMB_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  FA_X1 S2_2_7 ( .A(ab_2__7_), .B(CARRYB_1__7_), .CI(SUMB_1__8_), .CO(
        CARRYB_2__7_), .S(SUMB_2__7_) );
  FA_X1 S2_2_8 ( .A(ab_2__8_), .B(CARRYB_1__8_), .CI(SUMB_1__9_), .CO(
        CARRYB_2__8_), .S(SUMB_2__8_) );
  FA_X1 S2_2_9 ( .A(ab_2__9_), .B(CARRYB_1__9_), .CI(SUMB_1__10_), .CO(
        CARRYB_2__9_), .S(SUMB_2__9_) );
  FA_X1 S2_2_10 ( .A(ab_2__10_), .B(CARRYB_1__10_), .CI(SUMB_1__11_), .CO(
        CARRYB_2__10_), .S(SUMB_2__10_) );
  FA_X1 S2_2_11 ( .A(ab_2__11_), .B(CARRYB_1__11_), .CI(SUMB_1__12_), .CO(
        CARRYB_2__11_), .S(SUMB_2__11_) );
  FA_X1 S2_2_12 ( .A(ab_2__12_), .B(CARRYB_1__12_), .CI(SUMB_1__13_), .CO(
        CARRYB_2__12_), .S(SUMB_2__12_) );
  FA_X1 S2_2_13 ( .A(ab_2__13_), .B(CARRYB_1__13_), .CI(SUMB_1__14_), .CO(
        CARRYB_2__13_), .S(SUMB_2__13_) );
  FA_X1 S2_2_14 ( .A(ab_2__14_), .B(CARRYB_1__14_), .CI(SUMB_1__15_), .CO(
        CARRYB_2__14_), .S(SUMB_2__14_) );
  FA_X1 S2_2_15 ( .A(ab_2__15_), .B(CARRYB_1__15_), .CI(SUMB_1__16_), .CO(
        CARRYB_2__15_), .S(SUMB_2__15_) );
  FA_X1 S2_2_16 ( .A(ab_2__16_), .B(CARRYB_1__16_), .CI(SUMB_1__17_), .CO(
        CARRYB_2__16_), .S(SUMB_2__16_) );
  FA_X1 S2_2_17 ( .A(ab_2__17_), .B(CARRYB_1__17_), .CI(SUMB_1__18_), .CO(
        CARRYB_2__17_), .S(SUMB_2__17_) );
  FA_X1 S2_2_18 ( .A(ab_2__18_), .B(CARRYB_1__18_), .CI(SUMB_1__19_), .CO(
        CARRYB_2__18_), .S(SUMB_2__18_) );
  FA_X1 S2_2_19 ( .A(ab_2__19_), .B(CARRYB_1__19_), .CI(SUMB_1__20_), .CO(
        CARRYB_2__19_), .S(SUMB_2__19_) );
  FA_X1 S2_2_20 ( .A(ab_2__20_), .B(CARRYB_1__20_), .CI(SUMB_1__21_), .CO(
        CARRYB_2__20_), .S(SUMB_2__20_) );
  FA_X1 S2_2_21 ( .A(ab_2__21_), .B(CARRYB_1__21_), .CI(SUMB_1__22_), .CO(
        CARRYB_2__21_), .S(SUMB_2__21_) );
  FA_X1 S3_2_22 ( .A(ab_2__22_), .B(CARRYB_1__22_), .CI(ab_1__23_), .CO(
        CARRYB_2__22_), .S(SUMB_2__22_) );
  iir_filter_DW01_add_6 FS_1 ( .A({A1_45_, A1_44_, A1_43_, A1_42_, A1_41_, 
        A1_40_, A1_39_, A1_38_, A1_37_, A1_36_, A1_35_, A1_34_, A1_33_, A1_32_, 
        A1_31_, A1_30_, A1_29_, A1_28_, A1_27_, A1_26_, A1_25_, A1_24_, A1_23_, 
        A1_22_, A1_21_, A1_20_, A1_19_, A1_18_, A1_17_, A1_16_, A1_15_, A1_14_, 
        A1_13_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, A1_5_, 
        A1_4_, A1_3_, A1_2_, A1_1_, A1_0_}), .B({A2_45_, A2_44_, A2_43_, 
        A2_42_, A2_41_, A2_40_, A2_39_, A2_38_, A2_37_, A2_36_, A2_35_, A2_34_, 
        A2_33_, A2_32_, A2_31_, A2_30_, A2_29_, A2_28_, A2_27_, A2_26_, A2_25_, 
        A2_24_, A2_23_, A2_22_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({PRODUCT[47], SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, PRODUCT[44:22], SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21}) );
  BUF_X1 U2 ( .A(QB), .Z(n1) );
  BUF_X1 U3 ( .A(QB), .Z(n2) );
  BUF_X1 U4 ( .A(QA), .Z(n3) );
  BUF_X1 U5 ( .A(QA), .Z(n4) );
  INV_X1 U6 ( .A(A[2]), .ZN(n36) );
  INV_X1 U7 ( .A(A[3]), .ZN(n35) );
  INV_X1 U8 ( .A(A[4]), .ZN(n34) );
  INV_X1 U9 ( .A(A[5]), .ZN(n33) );
  INV_X1 U10 ( .A(A[6]), .ZN(n32) );
  INV_X1 U11 ( .A(B[1]), .ZN(n18) );
  INV_X1 U12 ( .A(A[1]), .ZN(n40) );
  INV_X1 U13 ( .A(B[0]), .ZN(n29) );
  INV_X1 U14 ( .A(A[0]), .ZN(n51) );
  INV_X1 U15 ( .A(B[22]), .ZN(n15) );
  INV_X1 U16 ( .A(B[21]), .ZN(n16) );
  INV_X1 U17 ( .A(B[20]), .ZN(n17) );
  INV_X1 U18 ( .A(B[19]), .ZN(n19) );
  INV_X1 U19 ( .A(B[18]), .ZN(n20) );
  INV_X1 U20 ( .A(B[17]), .ZN(n21) );
  INV_X1 U21 ( .A(B[16]), .ZN(n22) );
  INV_X1 U22 ( .A(B[15]), .ZN(n23) );
  INV_X1 U23 ( .A(B[14]), .ZN(n24) );
  INV_X1 U24 ( .A(B[13]), .ZN(n25) );
  INV_X1 U25 ( .A(B[12]), .ZN(n26) );
  INV_X1 U26 ( .A(B[11]), .ZN(n27) );
  INV_X1 U27 ( .A(B[10]), .ZN(n28) );
  INV_X1 U28 ( .A(B[9]), .ZN(n7) );
  INV_X1 U29 ( .A(B[8]), .ZN(n8) );
  INV_X1 U30 ( .A(B[7]), .ZN(n9) );
  INV_X1 U31 ( .A(B[6]), .ZN(n10) );
  INV_X1 U32 ( .A(B[5]), .ZN(n11) );
  INV_X1 U33 ( .A(B[4]), .ZN(n12) );
  INV_X1 U34 ( .A(B[3]), .ZN(n13) );
  INV_X1 U35 ( .A(B[2]), .ZN(n14) );
  INV_X1 U36 ( .A(A[7]), .ZN(n31) );
  INV_X1 U37 ( .A(A[8]), .ZN(n30) );
  INV_X1 U38 ( .A(A[10]), .ZN(n50) );
  INV_X1 U39 ( .A(A[11]), .ZN(n49) );
  INV_X1 U40 ( .A(A[12]), .ZN(n48) );
  INV_X1 U41 ( .A(A[13]), .ZN(n47) );
  INV_X1 U42 ( .A(A[14]), .ZN(n46) );
  INV_X1 U43 ( .A(A[9]), .ZN(n6) );
  INV_X1 U44 ( .A(A[22]), .ZN(n37) );
  INV_X1 U45 ( .A(A[15]), .ZN(n45) );
  INV_X1 U46 ( .A(A[16]), .ZN(n44) );
  INV_X1 U47 ( .A(A[17]), .ZN(n43) );
  INV_X1 U48 ( .A(A[18]), .ZN(n42) );
  INV_X1 U49 ( .A(A[19]), .ZN(n41) );
  INV_X1 U50 ( .A(A[20]), .ZN(n39) );
  INV_X1 U51 ( .A(A[21]), .ZN(n38) );
  AND2_X1 U52 ( .A1(SUMB_23__23_), .A2(CARRYB_23__22_), .ZN(A2_45_) );
  XOR2_X1 U53 ( .A(CARRYB_23__22_), .B(SUMB_23__23_), .Z(A1_44_) );
  AND2_X1 U54 ( .A1(SUMB_23__22_), .A2(CARRYB_23__21_), .ZN(A2_44_) );
  XOR2_X1 U55 ( .A(CARRYB_23__21_), .B(SUMB_23__22_), .Z(A1_43_) );
  AND2_X1 U56 ( .A1(SUMB_23__21_), .A2(CARRYB_23__20_), .ZN(A2_43_) );
  XOR2_X1 U57 ( .A(CARRYB_23__20_), .B(SUMB_23__21_), .Z(A1_42_) );
  AND2_X1 U58 ( .A1(SUMB_23__20_), .A2(CARRYB_23__19_), .ZN(A2_42_) );
  XOR2_X1 U59 ( .A(CARRYB_23__19_), .B(SUMB_23__20_), .Z(A1_41_) );
  AND2_X1 U60 ( .A1(SUMB_23__19_), .A2(CARRYB_23__18_), .ZN(A2_41_) );
  XOR2_X1 U61 ( .A(CARRYB_23__18_), .B(SUMB_23__19_), .Z(A1_40_) );
  AND2_X1 U62 ( .A1(SUMB_23__18_), .A2(CARRYB_23__17_), .ZN(A2_40_) );
  XOR2_X1 U63 ( .A(CARRYB_23__17_), .B(SUMB_23__18_), .Z(A1_39_) );
  AND2_X1 U64 ( .A1(SUMB_23__17_), .A2(CARRYB_23__16_), .ZN(A2_39_) );
  XOR2_X1 U65 ( .A(CARRYB_23__16_), .B(SUMB_23__17_), .Z(A1_38_) );
  AND2_X1 U66 ( .A1(SUMB_23__16_), .A2(CARRYB_23__15_), .ZN(A2_38_) );
  XOR2_X1 U67 ( .A(CARRYB_23__15_), .B(SUMB_23__16_), .Z(A1_37_) );
  AND2_X1 U68 ( .A1(SUMB_23__15_), .A2(CARRYB_23__14_), .ZN(A2_37_) );
  XOR2_X1 U69 ( .A(CARRYB_23__14_), .B(SUMB_23__15_), .Z(A1_36_) );
  AND2_X1 U70 ( .A1(SUMB_23__14_), .A2(CARRYB_23__13_), .ZN(A2_36_) );
  XOR2_X1 U71 ( .A(CARRYB_23__13_), .B(SUMB_23__14_), .Z(A1_35_) );
  AND2_X1 U72 ( .A1(SUMB_23__13_), .A2(CARRYB_23__12_), .ZN(A2_35_) );
  XOR2_X1 U73 ( .A(CARRYB_23__12_), .B(SUMB_23__13_), .Z(A1_34_) );
  AND2_X1 U74 ( .A1(SUMB_23__12_), .A2(CARRYB_23__11_), .ZN(A2_34_) );
  XOR2_X1 U75 ( .A(CARRYB_23__11_), .B(SUMB_23__12_), .Z(A1_33_) );
  AND2_X1 U76 ( .A1(SUMB_23__11_), .A2(CARRYB_23__10_), .ZN(A2_33_) );
  XOR2_X1 U77 ( .A(CARRYB_23__10_), .B(SUMB_23__11_), .Z(A1_32_) );
  AND2_X1 U78 ( .A1(SUMB_23__10_), .A2(CARRYB_23__9_), .ZN(A2_32_) );
  XOR2_X1 U79 ( .A(CARRYB_23__9_), .B(SUMB_23__10_), .Z(A1_31_) );
  AND2_X1 U80 ( .A1(SUMB_23__9_), .A2(CARRYB_23__8_), .ZN(A2_31_) );
  XOR2_X1 U81 ( .A(CARRYB_23__8_), .B(SUMB_23__9_), .Z(A1_30_) );
  AND2_X1 U82 ( .A1(SUMB_23__8_), .A2(CARRYB_23__7_), .ZN(A2_30_) );
  XOR2_X1 U83 ( .A(CARRYB_23__7_), .B(SUMB_23__8_), .Z(A1_29_) );
  AND2_X1 U84 ( .A1(SUMB_23__7_), .A2(CARRYB_23__6_), .ZN(A2_29_) );
  XOR2_X1 U85 ( .A(CARRYB_23__6_), .B(SUMB_23__7_), .Z(A1_28_) );
  AND2_X1 U86 ( .A1(SUMB_23__6_), .A2(CARRYB_23__5_), .ZN(A2_28_) );
  XOR2_X1 U87 ( .A(CARRYB_23__5_), .B(SUMB_23__6_), .Z(A1_27_) );
  AND2_X1 U88 ( .A1(SUMB_23__5_), .A2(CARRYB_23__4_), .ZN(A2_27_) );
  XOR2_X1 U89 ( .A(CARRYB_23__4_), .B(SUMB_23__5_), .Z(A1_26_) );
  AND2_X1 U90 ( .A1(SUMB_23__4_), .A2(CARRYB_23__3_), .ZN(A2_26_) );
  XOR2_X1 U91 ( .A(CARRYB_23__3_), .B(SUMB_23__4_), .Z(A1_25_) );
  AND2_X1 U92 ( .A1(SUMB_23__3_), .A2(CARRYB_23__2_), .ZN(A2_25_) );
  XOR2_X1 U93 ( .A(CARRYB_23__2_), .B(SUMB_23__3_), .Z(A1_24_) );
  AND2_X1 U94 ( .A1(SUMB_23__2_), .A2(CARRYB_23__1_), .ZN(A2_24_) );
  XOR2_X1 U95 ( .A(CARRYB_23__1_), .B(SUMB_23__2_), .Z(A1_23_) );
  AND2_X1 U96 ( .A1(SUMB_23__1_), .A2(CARRYB_23__0_), .ZN(A2_23_) );
  XOR2_X1 U97 ( .A(CARRYB_23__0_), .B(SUMB_23__1_), .Z(A1_22_) );
  AND2_X1 U98 ( .A1(ab_1__22_), .A2(ab_0__23_), .ZN(CARRYB_1__22_) );
  XOR2_X1 U99 ( .A(ab_1__22_), .B(ab_0__23_), .Z(SUMB_1__22_) );
  AND2_X1 U100 ( .A1(ab_1__21_), .A2(ab_0__22_), .ZN(CARRYB_1__21_) );
  XOR2_X1 U101 ( .A(ab_1__21_), .B(ab_0__22_), .Z(SUMB_1__21_) );
  AND2_X1 U102 ( .A1(ab_1__20_), .A2(ab_0__21_), .ZN(CARRYB_1__20_) );
  XOR2_X1 U103 ( .A(ab_1__20_), .B(ab_0__21_), .Z(SUMB_1__20_) );
  AND2_X1 U104 ( .A1(ab_1__19_), .A2(ab_0__20_), .ZN(CARRYB_1__19_) );
  XOR2_X1 U105 ( .A(ab_1__19_), .B(ab_0__20_), .Z(SUMB_1__19_) );
  AND2_X1 U106 ( .A1(ab_1__18_), .A2(ab_0__19_), .ZN(CARRYB_1__18_) );
  XOR2_X1 U107 ( .A(ab_1__18_), .B(ab_0__19_), .Z(SUMB_1__18_) );
  AND2_X1 U108 ( .A1(ab_1__17_), .A2(ab_0__18_), .ZN(CARRYB_1__17_) );
  XOR2_X1 U109 ( .A(ab_1__17_), .B(ab_0__18_), .Z(SUMB_1__17_) );
  AND2_X1 U110 ( .A1(ab_1__16_), .A2(ab_0__17_), .ZN(CARRYB_1__16_) );
  XOR2_X1 U111 ( .A(ab_1__16_), .B(ab_0__17_), .Z(SUMB_1__16_) );
  AND2_X1 U112 ( .A1(ab_1__15_), .A2(ab_0__16_), .ZN(CARRYB_1__15_) );
  XOR2_X1 U113 ( .A(ab_1__15_), .B(ab_0__16_), .Z(SUMB_1__15_) );
  AND2_X1 U114 ( .A1(ab_1__14_), .A2(ab_0__15_), .ZN(CARRYB_1__14_) );
  XOR2_X1 U115 ( .A(ab_1__14_), .B(ab_0__15_), .Z(SUMB_1__14_) );
  AND2_X1 U116 ( .A1(ab_1__13_), .A2(ab_0__14_), .ZN(CARRYB_1__13_) );
  XOR2_X1 U117 ( .A(ab_1__13_), .B(ab_0__14_), .Z(SUMB_1__13_) );
  AND2_X1 U118 ( .A1(ab_1__12_), .A2(ab_0__13_), .ZN(CARRYB_1__12_) );
  XOR2_X1 U119 ( .A(ab_1__12_), .B(ab_0__13_), .Z(SUMB_1__12_) );
  AND2_X1 U120 ( .A1(ab_1__11_), .A2(ab_0__12_), .ZN(CARRYB_1__11_) );
  XOR2_X1 U121 ( .A(ab_1__11_), .B(ab_0__12_), .Z(SUMB_1__11_) );
  AND2_X1 U122 ( .A1(ab_1__10_), .A2(ab_0__11_), .ZN(CARRYB_1__10_) );
  XOR2_X1 U123 ( .A(ab_1__10_), .B(ab_0__11_), .Z(SUMB_1__10_) );
  AND2_X1 U124 ( .A1(ab_1__9_), .A2(ab_0__10_), .ZN(CARRYB_1__9_) );
  XOR2_X1 U125 ( .A(ab_1__9_), .B(ab_0__10_), .Z(SUMB_1__9_) );
  AND2_X1 U126 ( .A1(ab_1__8_), .A2(ab_0__9_), .ZN(CARRYB_1__8_) );
  XOR2_X1 U127 ( .A(ab_1__8_), .B(ab_0__9_), .Z(SUMB_1__8_) );
  AND2_X1 U128 ( .A1(ab_1__7_), .A2(ab_0__8_), .ZN(CARRYB_1__7_) );
  XOR2_X1 U129 ( .A(ab_1__7_), .B(ab_0__8_), .Z(SUMB_1__7_) );
  AND2_X1 U130 ( .A1(ab_1__6_), .A2(ab_0__7_), .ZN(CARRYB_1__6_) );
  XOR2_X1 U131 ( .A(ab_1__6_), .B(ab_0__7_), .Z(SUMB_1__6_) );
  AND2_X1 U132 ( .A1(ab_1__5_), .A2(ab_0__6_), .ZN(CARRYB_1__5_) );
  XOR2_X1 U133 ( .A(ab_1__5_), .B(ab_0__6_), .Z(SUMB_1__5_) );
  AND2_X1 U134 ( .A1(ab_1__4_), .A2(ab_0__5_), .ZN(CARRYB_1__4_) );
  XOR2_X1 U135 ( .A(ab_1__4_), .B(ab_0__5_), .Z(SUMB_1__4_) );
  AND2_X1 U136 ( .A1(ab_1__3_), .A2(ab_0__4_), .ZN(CARRYB_1__3_) );
  XOR2_X1 U137 ( .A(ab_1__3_), .B(ab_0__4_), .Z(SUMB_1__3_) );
  AND2_X1 U138 ( .A1(ab_1__2_), .A2(ab_0__3_), .ZN(CARRYB_1__2_) );
  XOR2_X1 U139 ( .A(ab_1__2_), .B(ab_0__3_), .Z(SUMB_1__2_) );
  AND2_X1 U140 ( .A1(ab_1__1_), .A2(ab_0__2_), .ZN(CARRYB_1__1_) );
  XOR2_X1 U141 ( .A(ab_1__1_), .B(ab_0__2_), .Z(SUMB_1__1_) );
  NOR2_X1 U142 ( .A1(n6), .A2(n7), .ZN(ab_9__9_) );
  NOR2_X1 U143 ( .A1(n6), .A2(n8), .ZN(ab_9__8_) );
  NOR2_X1 U144 ( .A1(n6), .A2(n9), .ZN(ab_9__7_) );
  NOR2_X1 U145 ( .A1(n6), .A2(n10), .ZN(ab_9__6_) );
  NOR2_X1 U146 ( .A1(n6), .A2(n11), .ZN(ab_9__5_) );
  NOR2_X1 U147 ( .A1(n6), .A2(n12), .ZN(ab_9__4_) );
  NOR2_X1 U148 ( .A1(n6), .A2(n13), .ZN(ab_9__3_) );
  NOR2_X1 U149 ( .A1(n6), .A2(n14), .ZN(ab_9__2_) );
  NOR2_X1 U150 ( .A1(A[9]), .A2(n1), .ZN(ab_9__23_) );
  NOR2_X1 U151 ( .A1(n6), .A2(n15), .ZN(ab_9__22_) );
  NOR2_X1 U152 ( .A1(n6), .A2(n16), .ZN(ab_9__21_) );
  NOR2_X1 U153 ( .A1(n6), .A2(n17), .ZN(ab_9__20_) );
  NOR2_X1 U154 ( .A1(n6), .A2(n18), .ZN(ab_9__1_) );
  NOR2_X1 U155 ( .A1(n6), .A2(n19), .ZN(ab_9__19_) );
  NOR2_X1 U156 ( .A1(n6), .A2(n20), .ZN(ab_9__18_) );
  NOR2_X1 U157 ( .A1(n6), .A2(n21), .ZN(ab_9__17_) );
  NOR2_X1 U158 ( .A1(n6), .A2(n22), .ZN(ab_9__16_) );
  NOR2_X1 U159 ( .A1(n6), .A2(n23), .ZN(ab_9__15_) );
  NOR2_X1 U160 ( .A1(n6), .A2(n24), .ZN(ab_9__14_) );
  NOR2_X1 U161 ( .A1(n6), .A2(n25), .ZN(ab_9__13_) );
  NOR2_X1 U162 ( .A1(n6), .A2(n26), .ZN(ab_9__12_) );
  NOR2_X1 U163 ( .A1(n6), .A2(n27), .ZN(ab_9__11_) );
  NOR2_X1 U164 ( .A1(n6), .A2(n28), .ZN(ab_9__10_) );
  NOR2_X1 U165 ( .A1(n6), .A2(n29), .ZN(ab_9__0_) );
  NOR2_X1 U166 ( .A1(n7), .A2(n30), .ZN(ab_8__9_) );
  NOR2_X1 U167 ( .A1(n8), .A2(n30), .ZN(ab_8__8_) );
  NOR2_X1 U168 ( .A1(n9), .A2(n30), .ZN(ab_8__7_) );
  NOR2_X1 U169 ( .A1(n10), .A2(n30), .ZN(ab_8__6_) );
  NOR2_X1 U170 ( .A1(n11), .A2(n30), .ZN(ab_8__5_) );
  NOR2_X1 U171 ( .A1(n12), .A2(n30), .ZN(ab_8__4_) );
  NOR2_X1 U172 ( .A1(n13), .A2(n30), .ZN(ab_8__3_) );
  NOR2_X1 U173 ( .A1(n14), .A2(n30), .ZN(ab_8__2_) );
  NOR2_X1 U174 ( .A1(A[8]), .A2(n1), .ZN(ab_8__23_) );
  NOR2_X1 U175 ( .A1(n15), .A2(n30), .ZN(ab_8__22_) );
  NOR2_X1 U176 ( .A1(n16), .A2(n30), .ZN(ab_8__21_) );
  NOR2_X1 U177 ( .A1(n17), .A2(n30), .ZN(ab_8__20_) );
  NOR2_X1 U178 ( .A1(n18), .A2(n30), .ZN(ab_8__1_) );
  NOR2_X1 U179 ( .A1(n19), .A2(n30), .ZN(ab_8__19_) );
  NOR2_X1 U180 ( .A1(n20), .A2(n30), .ZN(ab_8__18_) );
  NOR2_X1 U181 ( .A1(n21), .A2(n30), .ZN(ab_8__17_) );
  NOR2_X1 U182 ( .A1(n22), .A2(n30), .ZN(ab_8__16_) );
  NOR2_X1 U183 ( .A1(n23), .A2(n30), .ZN(ab_8__15_) );
  NOR2_X1 U184 ( .A1(n24), .A2(n30), .ZN(ab_8__14_) );
  NOR2_X1 U185 ( .A1(n25), .A2(n30), .ZN(ab_8__13_) );
  NOR2_X1 U186 ( .A1(n26), .A2(n30), .ZN(ab_8__12_) );
  NOR2_X1 U187 ( .A1(n27), .A2(n30), .ZN(ab_8__11_) );
  NOR2_X1 U188 ( .A1(n28), .A2(n30), .ZN(ab_8__10_) );
  NOR2_X1 U189 ( .A1(n29), .A2(n30), .ZN(ab_8__0_) );
  NOR2_X1 U190 ( .A1(n7), .A2(n31), .ZN(ab_7__9_) );
  NOR2_X1 U191 ( .A1(n8), .A2(n31), .ZN(ab_7__8_) );
  NOR2_X1 U192 ( .A1(n9), .A2(n31), .ZN(ab_7__7_) );
  NOR2_X1 U193 ( .A1(n10), .A2(n31), .ZN(ab_7__6_) );
  NOR2_X1 U194 ( .A1(n11), .A2(n31), .ZN(ab_7__5_) );
  NOR2_X1 U195 ( .A1(n12), .A2(n31), .ZN(ab_7__4_) );
  NOR2_X1 U196 ( .A1(n13), .A2(n31), .ZN(ab_7__3_) );
  NOR2_X1 U197 ( .A1(n14), .A2(n31), .ZN(ab_7__2_) );
  NOR2_X1 U198 ( .A1(A[7]), .A2(n1), .ZN(ab_7__23_) );
  NOR2_X1 U199 ( .A1(n15), .A2(n31), .ZN(ab_7__22_) );
  NOR2_X1 U200 ( .A1(n16), .A2(n31), .ZN(ab_7__21_) );
  NOR2_X1 U201 ( .A1(n17), .A2(n31), .ZN(ab_7__20_) );
  NOR2_X1 U202 ( .A1(n18), .A2(n31), .ZN(ab_7__1_) );
  NOR2_X1 U203 ( .A1(n19), .A2(n31), .ZN(ab_7__19_) );
  NOR2_X1 U204 ( .A1(n20), .A2(n31), .ZN(ab_7__18_) );
  NOR2_X1 U205 ( .A1(n21), .A2(n31), .ZN(ab_7__17_) );
  NOR2_X1 U206 ( .A1(n22), .A2(n31), .ZN(ab_7__16_) );
  NOR2_X1 U207 ( .A1(n23), .A2(n31), .ZN(ab_7__15_) );
  NOR2_X1 U208 ( .A1(n24), .A2(n31), .ZN(ab_7__14_) );
  NOR2_X1 U209 ( .A1(n25), .A2(n31), .ZN(ab_7__13_) );
  NOR2_X1 U210 ( .A1(n26), .A2(n31), .ZN(ab_7__12_) );
  NOR2_X1 U211 ( .A1(n27), .A2(n31), .ZN(ab_7__11_) );
  NOR2_X1 U212 ( .A1(n28), .A2(n31), .ZN(ab_7__10_) );
  NOR2_X1 U213 ( .A1(n29), .A2(n31), .ZN(ab_7__0_) );
  NOR2_X1 U214 ( .A1(n7), .A2(n32), .ZN(ab_6__9_) );
  NOR2_X1 U215 ( .A1(n8), .A2(n32), .ZN(ab_6__8_) );
  NOR2_X1 U216 ( .A1(n9), .A2(n32), .ZN(ab_6__7_) );
  NOR2_X1 U217 ( .A1(n10), .A2(n32), .ZN(ab_6__6_) );
  NOR2_X1 U218 ( .A1(n11), .A2(n32), .ZN(ab_6__5_) );
  NOR2_X1 U219 ( .A1(n12), .A2(n32), .ZN(ab_6__4_) );
  NOR2_X1 U220 ( .A1(n13), .A2(n32), .ZN(ab_6__3_) );
  NOR2_X1 U221 ( .A1(n14), .A2(n32), .ZN(ab_6__2_) );
  NOR2_X1 U222 ( .A1(A[6]), .A2(n1), .ZN(ab_6__23_) );
  NOR2_X1 U223 ( .A1(n15), .A2(n32), .ZN(ab_6__22_) );
  NOR2_X1 U224 ( .A1(n16), .A2(n32), .ZN(ab_6__21_) );
  NOR2_X1 U225 ( .A1(n17), .A2(n32), .ZN(ab_6__20_) );
  NOR2_X1 U226 ( .A1(n18), .A2(n32), .ZN(ab_6__1_) );
  NOR2_X1 U227 ( .A1(n19), .A2(n32), .ZN(ab_6__19_) );
  NOR2_X1 U228 ( .A1(n20), .A2(n32), .ZN(ab_6__18_) );
  NOR2_X1 U229 ( .A1(n21), .A2(n32), .ZN(ab_6__17_) );
  NOR2_X1 U230 ( .A1(n22), .A2(n32), .ZN(ab_6__16_) );
  NOR2_X1 U231 ( .A1(n23), .A2(n32), .ZN(ab_6__15_) );
  NOR2_X1 U232 ( .A1(n24), .A2(n32), .ZN(ab_6__14_) );
  NOR2_X1 U233 ( .A1(n25), .A2(n32), .ZN(ab_6__13_) );
  NOR2_X1 U234 ( .A1(n26), .A2(n32), .ZN(ab_6__12_) );
  NOR2_X1 U235 ( .A1(n27), .A2(n32), .ZN(ab_6__11_) );
  NOR2_X1 U236 ( .A1(n28), .A2(n32), .ZN(ab_6__10_) );
  NOR2_X1 U237 ( .A1(n29), .A2(n32), .ZN(ab_6__0_) );
  NOR2_X1 U238 ( .A1(n7), .A2(n33), .ZN(ab_5__9_) );
  NOR2_X1 U239 ( .A1(n8), .A2(n33), .ZN(ab_5__8_) );
  NOR2_X1 U240 ( .A1(n9), .A2(n33), .ZN(ab_5__7_) );
  NOR2_X1 U241 ( .A1(n10), .A2(n33), .ZN(ab_5__6_) );
  NOR2_X1 U242 ( .A1(n11), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U243 ( .A1(n12), .A2(n33), .ZN(ab_5__4_) );
  NOR2_X1 U244 ( .A1(n13), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U245 ( .A1(n14), .A2(n33), .ZN(ab_5__2_) );
  NOR2_X1 U246 ( .A1(A[5]), .A2(n1), .ZN(ab_5__23_) );
  NOR2_X1 U247 ( .A1(n15), .A2(n33), .ZN(ab_5__22_) );
  NOR2_X1 U248 ( .A1(n16), .A2(n33), .ZN(ab_5__21_) );
  NOR2_X1 U249 ( .A1(n17), .A2(n33), .ZN(ab_5__20_) );
  NOR2_X1 U250 ( .A1(n18), .A2(n33), .ZN(ab_5__1_) );
  NOR2_X1 U251 ( .A1(n19), .A2(n33), .ZN(ab_5__19_) );
  NOR2_X1 U252 ( .A1(n20), .A2(n33), .ZN(ab_5__18_) );
  NOR2_X1 U253 ( .A1(n21), .A2(n33), .ZN(ab_5__17_) );
  NOR2_X1 U254 ( .A1(n22), .A2(n33), .ZN(ab_5__16_) );
  NOR2_X1 U255 ( .A1(n23), .A2(n33), .ZN(ab_5__15_) );
  NOR2_X1 U256 ( .A1(n24), .A2(n33), .ZN(ab_5__14_) );
  NOR2_X1 U257 ( .A1(n25), .A2(n33), .ZN(ab_5__13_) );
  NOR2_X1 U258 ( .A1(n26), .A2(n33), .ZN(ab_5__12_) );
  NOR2_X1 U259 ( .A1(n27), .A2(n33), .ZN(ab_5__11_) );
  NOR2_X1 U260 ( .A1(n28), .A2(n33), .ZN(ab_5__10_) );
  NOR2_X1 U261 ( .A1(n29), .A2(n33), .ZN(ab_5__0_) );
  NOR2_X1 U262 ( .A1(n7), .A2(n34), .ZN(ab_4__9_) );
  NOR2_X1 U263 ( .A1(n8), .A2(n34), .ZN(ab_4__8_) );
  NOR2_X1 U264 ( .A1(n9), .A2(n34), .ZN(ab_4__7_) );
  NOR2_X1 U265 ( .A1(n10), .A2(n34), .ZN(ab_4__6_) );
  NOR2_X1 U266 ( .A1(n11), .A2(n34), .ZN(ab_4__5_) );
  NOR2_X1 U267 ( .A1(n12), .A2(n34), .ZN(ab_4__4_) );
  NOR2_X1 U268 ( .A1(n13), .A2(n34), .ZN(ab_4__3_) );
  NOR2_X1 U269 ( .A1(n14), .A2(n34), .ZN(ab_4__2_) );
  NOR2_X1 U270 ( .A1(A[4]), .A2(n1), .ZN(ab_4__23_) );
  NOR2_X1 U271 ( .A1(n15), .A2(n34), .ZN(ab_4__22_) );
  NOR2_X1 U272 ( .A1(n16), .A2(n34), .ZN(ab_4__21_) );
  NOR2_X1 U273 ( .A1(n17), .A2(n34), .ZN(ab_4__20_) );
  NOR2_X1 U274 ( .A1(n18), .A2(n34), .ZN(ab_4__1_) );
  NOR2_X1 U275 ( .A1(n19), .A2(n34), .ZN(ab_4__19_) );
  NOR2_X1 U276 ( .A1(n20), .A2(n34), .ZN(ab_4__18_) );
  NOR2_X1 U277 ( .A1(n21), .A2(n34), .ZN(ab_4__17_) );
  NOR2_X1 U278 ( .A1(n22), .A2(n34), .ZN(ab_4__16_) );
  NOR2_X1 U279 ( .A1(n23), .A2(n34), .ZN(ab_4__15_) );
  NOR2_X1 U280 ( .A1(n24), .A2(n34), .ZN(ab_4__14_) );
  NOR2_X1 U281 ( .A1(n25), .A2(n34), .ZN(ab_4__13_) );
  NOR2_X1 U282 ( .A1(n26), .A2(n34), .ZN(ab_4__12_) );
  NOR2_X1 U283 ( .A1(n27), .A2(n34), .ZN(ab_4__11_) );
  NOR2_X1 U284 ( .A1(n28), .A2(n34), .ZN(ab_4__10_) );
  NOR2_X1 U285 ( .A1(n29), .A2(n34), .ZN(ab_4__0_) );
  NOR2_X1 U286 ( .A1(n7), .A2(n35), .ZN(ab_3__9_) );
  NOR2_X1 U287 ( .A1(n8), .A2(n35), .ZN(ab_3__8_) );
  NOR2_X1 U288 ( .A1(n9), .A2(n35), .ZN(ab_3__7_) );
  NOR2_X1 U289 ( .A1(n10), .A2(n35), .ZN(ab_3__6_) );
  NOR2_X1 U290 ( .A1(n11), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U291 ( .A1(n12), .A2(n35), .ZN(ab_3__4_) );
  NOR2_X1 U292 ( .A1(n13), .A2(n35), .ZN(ab_3__3_) );
  NOR2_X1 U293 ( .A1(n14), .A2(n35), .ZN(ab_3__2_) );
  NOR2_X1 U294 ( .A1(A[3]), .A2(n1), .ZN(ab_3__23_) );
  NOR2_X1 U295 ( .A1(n15), .A2(n35), .ZN(ab_3__22_) );
  NOR2_X1 U296 ( .A1(n16), .A2(n35), .ZN(ab_3__21_) );
  NOR2_X1 U297 ( .A1(n17), .A2(n35), .ZN(ab_3__20_) );
  NOR2_X1 U298 ( .A1(n18), .A2(n35), .ZN(ab_3__1_) );
  NOR2_X1 U299 ( .A1(n19), .A2(n35), .ZN(ab_3__19_) );
  NOR2_X1 U300 ( .A1(n20), .A2(n35), .ZN(ab_3__18_) );
  NOR2_X1 U301 ( .A1(n21), .A2(n35), .ZN(ab_3__17_) );
  NOR2_X1 U302 ( .A1(n22), .A2(n35), .ZN(ab_3__16_) );
  NOR2_X1 U303 ( .A1(n23), .A2(n35), .ZN(ab_3__15_) );
  NOR2_X1 U304 ( .A1(n24), .A2(n35), .ZN(ab_3__14_) );
  NOR2_X1 U305 ( .A1(n25), .A2(n35), .ZN(ab_3__13_) );
  NOR2_X1 U306 ( .A1(n26), .A2(n35), .ZN(ab_3__12_) );
  NOR2_X1 U307 ( .A1(n27), .A2(n35), .ZN(ab_3__11_) );
  NOR2_X1 U308 ( .A1(n28), .A2(n35), .ZN(ab_3__10_) );
  NOR2_X1 U309 ( .A1(n29), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U310 ( .A1(n7), .A2(n36), .ZN(ab_2__9_) );
  NOR2_X1 U311 ( .A1(n8), .A2(n36), .ZN(ab_2__8_) );
  NOR2_X1 U312 ( .A1(n9), .A2(n36), .ZN(ab_2__7_) );
  NOR2_X1 U313 ( .A1(n10), .A2(n36), .ZN(ab_2__6_) );
  NOR2_X1 U314 ( .A1(n11), .A2(n36), .ZN(ab_2__5_) );
  NOR2_X1 U315 ( .A1(n12), .A2(n36), .ZN(ab_2__4_) );
  NOR2_X1 U316 ( .A1(n13), .A2(n36), .ZN(ab_2__3_) );
  NOR2_X1 U317 ( .A1(n14), .A2(n36), .ZN(ab_2__2_) );
  NOR2_X1 U318 ( .A1(A[2]), .A2(n1), .ZN(ab_2__23_) );
  NOR2_X1 U319 ( .A1(n15), .A2(n36), .ZN(ab_2__22_) );
  NOR2_X1 U320 ( .A1(n16), .A2(n36), .ZN(ab_2__21_) );
  NOR2_X1 U321 ( .A1(n17), .A2(n36), .ZN(ab_2__20_) );
  NOR2_X1 U322 ( .A1(n18), .A2(n36), .ZN(ab_2__1_) );
  NOR2_X1 U323 ( .A1(n19), .A2(n36), .ZN(ab_2__19_) );
  NOR2_X1 U324 ( .A1(n20), .A2(n36), .ZN(ab_2__18_) );
  NOR2_X1 U325 ( .A1(n21), .A2(n36), .ZN(ab_2__17_) );
  NOR2_X1 U326 ( .A1(n22), .A2(n36), .ZN(ab_2__16_) );
  NOR2_X1 U327 ( .A1(n23), .A2(n36), .ZN(ab_2__15_) );
  NOR2_X1 U328 ( .A1(n24), .A2(n36), .ZN(ab_2__14_) );
  NOR2_X1 U329 ( .A1(n25), .A2(n36), .ZN(ab_2__13_) );
  NOR2_X1 U330 ( .A1(n26), .A2(n36), .ZN(ab_2__12_) );
  NOR2_X1 U331 ( .A1(n27), .A2(n36), .ZN(ab_2__11_) );
  NOR2_X1 U332 ( .A1(n28), .A2(n36), .ZN(ab_2__10_) );
  NOR2_X1 U333 ( .A1(n29), .A2(n36), .ZN(ab_2__0_) );
  NOR2_X1 U334 ( .A1(B[9]), .A2(n4), .ZN(ab_23__9_) );
  NOR2_X1 U335 ( .A1(B[8]), .A2(n4), .ZN(ab_23__8_) );
  NOR2_X1 U336 ( .A1(B[7]), .A2(n4), .ZN(ab_23__7_) );
  NOR2_X1 U337 ( .A1(B[6]), .A2(n4), .ZN(ab_23__6_) );
  NOR2_X1 U338 ( .A1(B[5]), .A2(n3), .ZN(ab_23__5_) );
  NOR2_X1 U339 ( .A1(B[4]), .A2(n3), .ZN(ab_23__4_) );
  NOR2_X1 U340 ( .A1(B[3]), .A2(n3), .ZN(ab_23__3_) );
  NOR2_X1 U341 ( .A1(B[2]), .A2(n3), .ZN(ab_23__2_) );
  NOR2_X1 U342 ( .A1(n1), .A2(n3), .ZN(ab_23__23_) );
  NOR2_X1 U343 ( .A1(B[22]), .A2(n3), .ZN(ab_23__22_) );
  NOR2_X1 U344 ( .A1(B[21]), .A2(n3), .ZN(ab_23__21_) );
  NOR2_X1 U345 ( .A1(B[20]), .A2(n3), .ZN(ab_23__20_) );
  NOR2_X1 U346 ( .A1(B[1]), .A2(n3), .ZN(ab_23__1_) );
  NOR2_X1 U347 ( .A1(B[19]), .A2(n3), .ZN(ab_23__19_) );
  NOR2_X1 U348 ( .A1(B[18]), .A2(n3), .ZN(ab_23__18_) );
  NOR2_X1 U349 ( .A1(B[17]), .A2(n3), .ZN(ab_23__17_) );
  NOR2_X1 U350 ( .A1(B[16]), .A2(n3), .ZN(ab_23__16_) );
  NOR2_X1 U351 ( .A1(B[15]), .A2(n3), .ZN(ab_23__15_) );
  NOR2_X1 U352 ( .A1(B[14]), .A2(n3), .ZN(ab_23__14_) );
  NOR2_X1 U353 ( .A1(B[13]), .A2(n3), .ZN(ab_23__13_) );
  NOR2_X1 U354 ( .A1(B[12]), .A2(n3), .ZN(ab_23__12_) );
  NOR2_X1 U355 ( .A1(B[11]), .A2(n3), .ZN(ab_23__11_) );
  NOR2_X1 U356 ( .A1(B[10]), .A2(n3), .ZN(ab_23__10_) );
  NOR2_X1 U357 ( .A1(B[0]), .A2(n3), .ZN(ab_23__0_) );
  NOR2_X1 U358 ( .A1(n7), .A2(n37), .ZN(ab_22__9_) );
  NOR2_X1 U359 ( .A1(n8), .A2(n37), .ZN(ab_22__8_) );
  NOR2_X1 U360 ( .A1(n9), .A2(n37), .ZN(ab_22__7_) );
  NOR2_X1 U361 ( .A1(n10), .A2(n37), .ZN(ab_22__6_) );
  NOR2_X1 U362 ( .A1(n11), .A2(n37), .ZN(ab_22__5_) );
  NOR2_X1 U363 ( .A1(n12), .A2(n37), .ZN(ab_22__4_) );
  NOR2_X1 U364 ( .A1(n13), .A2(n37), .ZN(ab_22__3_) );
  NOR2_X1 U365 ( .A1(n14), .A2(n37), .ZN(ab_22__2_) );
  NOR2_X1 U366 ( .A1(A[22]), .A2(n1), .ZN(ab_22__23_) );
  NOR2_X1 U367 ( .A1(n15), .A2(n37), .ZN(ab_22__22_) );
  NOR2_X1 U368 ( .A1(n16), .A2(n37), .ZN(ab_22__21_) );
  NOR2_X1 U369 ( .A1(n17), .A2(n37), .ZN(ab_22__20_) );
  NOR2_X1 U370 ( .A1(n18), .A2(n37), .ZN(ab_22__1_) );
  NOR2_X1 U371 ( .A1(n19), .A2(n37), .ZN(ab_22__19_) );
  NOR2_X1 U372 ( .A1(n20), .A2(n37), .ZN(ab_22__18_) );
  NOR2_X1 U373 ( .A1(n21), .A2(n37), .ZN(ab_22__17_) );
  NOR2_X1 U374 ( .A1(n22), .A2(n37), .ZN(ab_22__16_) );
  NOR2_X1 U375 ( .A1(n23), .A2(n37), .ZN(ab_22__15_) );
  NOR2_X1 U376 ( .A1(n24), .A2(n37), .ZN(ab_22__14_) );
  NOR2_X1 U377 ( .A1(n25), .A2(n37), .ZN(ab_22__13_) );
  NOR2_X1 U378 ( .A1(n26), .A2(n37), .ZN(ab_22__12_) );
  NOR2_X1 U379 ( .A1(n27), .A2(n37), .ZN(ab_22__11_) );
  NOR2_X1 U380 ( .A1(n28), .A2(n37), .ZN(ab_22__10_) );
  NOR2_X1 U381 ( .A1(n29), .A2(n37), .ZN(ab_22__0_) );
  NOR2_X1 U382 ( .A1(n7), .A2(n38), .ZN(ab_21__9_) );
  NOR2_X1 U383 ( .A1(n8), .A2(n38), .ZN(ab_21__8_) );
  NOR2_X1 U384 ( .A1(n9), .A2(n38), .ZN(ab_21__7_) );
  NOR2_X1 U385 ( .A1(n10), .A2(n38), .ZN(ab_21__6_) );
  NOR2_X1 U386 ( .A1(n11), .A2(n38), .ZN(ab_21__5_) );
  NOR2_X1 U387 ( .A1(n12), .A2(n38), .ZN(ab_21__4_) );
  NOR2_X1 U388 ( .A1(n13), .A2(n38), .ZN(ab_21__3_) );
  NOR2_X1 U389 ( .A1(n14), .A2(n38), .ZN(ab_21__2_) );
  NOR2_X1 U390 ( .A1(A[21]), .A2(n1), .ZN(ab_21__23_) );
  NOR2_X1 U391 ( .A1(n15), .A2(n38), .ZN(ab_21__22_) );
  NOR2_X1 U392 ( .A1(n16), .A2(n38), .ZN(ab_21__21_) );
  NOR2_X1 U393 ( .A1(n17), .A2(n38), .ZN(ab_21__20_) );
  NOR2_X1 U394 ( .A1(n18), .A2(n38), .ZN(ab_21__1_) );
  NOR2_X1 U395 ( .A1(n19), .A2(n38), .ZN(ab_21__19_) );
  NOR2_X1 U396 ( .A1(n20), .A2(n38), .ZN(ab_21__18_) );
  NOR2_X1 U397 ( .A1(n21), .A2(n38), .ZN(ab_21__17_) );
  NOR2_X1 U398 ( .A1(n22), .A2(n38), .ZN(ab_21__16_) );
  NOR2_X1 U399 ( .A1(n23), .A2(n38), .ZN(ab_21__15_) );
  NOR2_X1 U400 ( .A1(n24), .A2(n38), .ZN(ab_21__14_) );
  NOR2_X1 U401 ( .A1(n25), .A2(n38), .ZN(ab_21__13_) );
  NOR2_X1 U402 ( .A1(n26), .A2(n38), .ZN(ab_21__12_) );
  NOR2_X1 U403 ( .A1(n27), .A2(n38), .ZN(ab_21__11_) );
  NOR2_X1 U404 ( .A1(n28), .A2(n38), .ZN(ab_21__10_) );
  NOR2_X1 U405 ( .A1(n29), .A2(n38), .ZN(ab_21__0_) );
  NOR2_X1 U406 ( .A1(n7), .A2(n39), .ZN(ab_20__9_) );
  NOR2_X1 U407 ( .A1(n8), .A2(n39), .ZN(ab_20__8_) );
  NOR2_X1 U408 ( .A1(n9), .A2(n39), .ZN(ab_20__7_) );
  NOR2_X1 U409 ( .A1(n10), .A2(n39), .ZN(ab_20__6_) );
  NOR2_X1 U410 ( .A1(n11), .A2(n39), .ZN(ab_20__5_) );
  NOR2_X1 U411 ( .A1(n12), .A2(n39), .ZN(ab_20__4_) );
  NOR2_X1 U412 ( .A1(n13), .A2(n39), .ZN(ab_20__3_) );
  NOR2_X1 U413 ( .A1(n14), .A2(n39), .ZN(ab_20__2_) );
  NOR2_X1 U414 ( .A1(A[20]), .A2(n1), .ZN(ab_20__23_) );
  NOR2_X1 U415 ( .A1(n15), .A2(n39), .ZN(ab_20__22_) );
  NOR2_X1 U416 ( .A1(n16), .A2(n39), .ZN(ab_20__21_) );
  NOR2_X1 U417 ( .A1(n17), .A2(n39), .ZN(ab_20__20_) );
  NOR2_X1 U418 ( .A1(n18), .A2(n39), .ZN(ab_20__1_) );
  NOR2_X1 U419 ( .A1(n19), .A2(n39), .ZN(ab_20__19_) );
  NOR2_X1 U420 ( .A1(n20), .A2(n39), .ZN(ab_20__18_) );
  NOR2_X1 U421 ( .A1(n21), .A2(n39), .ZN(ab_20__17_) );
  NOR2_X1 U422 ( .A1(n22), .A2(n39), .ZN(ab_20__16_) );
  NOR2_X1 U423 ( .A1(n23), .A2(n39), .ZN(ab_20__15_) );
  NOR2_X1 U424 ( .A1(n24), .A2(n39), .ZN(ab_20__14_) );
  NOR2_X1 U425 ( .A1(n25), .A2(n39), .ZN(ab_20__13_) );
  NOR2_X1 U426 ( .A1(n26), .A2(n39), .ZN(ab_20__12_) );
  NOR2_X1 U427 ( .A1(n27), .A2(n39), .ZN(ab_20__11_) );
  NOR2_X1 U428 ( .A1(n28), .A2(n39), .ZN(ab_20__10_) );
  NOR2_X1 U429 ( .A1(n29), .A2(n39), .ZN(ab_20__0_) );
  NOR2_X1 U430 ( .A1(n7), .A2(n40), .ZN(ab_1__9_) );
  NOR2_X1 U431 ( .A1(n8), .A2(n40), .ZN(ab_1__8_) );
  NOR2_X1 U432 ( .A1(n9), .A2(n40), .ZN(ab_1__7_) );
  NOR2_X1 U433 ( .A1(n10), .A2(n40), .ZN(ab_1__6_) );
  NOR2_X1 U434 ( .A1(n11), .A2(n40), .ZN(ab_1__5_) );
  NOR2_X1 U435 ( .A1(n12), .A2(n40), .ZN(ab_1__4_) );
  NOR2_X1 U436 ( .A1(n13), .A2(n40), .ZN(ab_1__3_) );
  NOR2_X1 U437 ( .A1(n14), .A2(n40), .ZN(ab_1__2_) );
  NOR2_X1 U438 ( .A1(A[1]), .A2(n1), .ZN(ab_1__23_) );
  NOR2_X1 U439 ( .A1(n15), .A2(n40), .ZN(ab_1__22_) );
  NOR2_X1 U440 ( .A1(n16), .A2(n40), .ZN(ab_1__21_) );
  NOR2_X1 U441 ( .A1(n17), .A2(n40), .ZN(ab_1__20_) );
  NOR2_X1 U442 ( .A1(n19), .A2(n40), .ZN(ab_1__19_) );
  NOR2_X1 U443 ( .A1(n20), .A2(n40), .ZN(ab_1__18_) );
  NOR2_X1 U444 ( .A1(n21), .A2(n40), .ZN(ab_1__17_) );
  NOR2_X1 U445 ( .A1(n22), .A2(n40), .ZN(ab_1__16_) );
  NOR2_X1 U446 ( .A1(n23), .A2(n40), .ZN(ab_1__15_) );
  NOR2_X1 U447 ( .A1(n24), .A2(n40), .ZN(ab_1__14_) );
  NOR2_X1 U448 ( .A1(n25), .A2(n40), .ZN(ab_1__13_) );
  NOR2_X1 U449 ( .A1(n26), .A2(n40), .ZN(ab_1__12_) );
  NOR2_X1 U450 ( .A1(n27), .A2(n40), .ZN(ab_1__11_) );
  NOR2_X1 U451 ( .A1(n28), .A2(n40), .ZN(ab_1__10_) );
  NOR2_X1 U452 ( .A1(n7), .A2(n41), .ZN(ab_19__9_) );
  NOR2_X1 U453 ( .A1(n8), .A2(n41), .ZN(ab_19__8_) );
  NOR2_X1 U454 ( .A1(n9), .A2(n41), .ZN(ab_19__7_) );
  NOR2_X1 U455 ( .A1(n10), .A2(n41), .ZN(ab_19__6_) );
  NOR2_X1 U456 ( .A1(n11), .A2(n41), .ZN(ab_19__5_) );
  NOR2_X1 U457 ( .A1(n12), .A2(n41), .ZN(ab_19__4_) );
  NOR2_X1 U458 ( .A1(n13), .A2(n41), .ZN(ab_19__3_) );
  NOR2_X1 U459 ( .A1(n14), .A2(n41), .ZN(ab_19__2_) );
  NOR2_X1 U460 ( .A1(A[19]), .A2(n1), .ZN(ab_19__23_) );
  NOR2_X1 U461 ( .A1(n15), .A2(n41), .ZN(ab_19__22_) );
  NOR2_X1 U462 ( .A1(n16), .A2(n41), .ZN(ab_19__21_) );
  NOR2_X1 U463 ( .A1(n17), .A2(n41), .ZN(ab_19__20_) );
  NOR2_X1 U464 ( .A1(n18), .A2(n41), .ZN(ab_19__1_) );
  NOR2_X1 U465 ( .A1(n19), .A2(n41), .ZN(ab_19__19_) );
  NOR2_X1 U466 ( .A1(n20), .A2(n41), .ZN(ab_19__18_) );
  NOR2_X1 U467 ( .A1(n21), .A2(n41), .ZN(ab_19__17_) );
  NOR2_X1 U468 ( .A1(n22), .A2(n41), .ZN(ab_19__16_) );
  NOR2_X1 U469 ( .A1(n23), .A2(n41), .ZN(ab_19__15_) );
  NOR2_X1 U470 ( .A1(n24), .A2(n41), .ZN(ab_19__14_) );
  NOR2_X1 U471 ( .A1(n25), .A2(n41), .ZN(ab_19__13_) );
  NOR2_X1 U472 ( .A1(n26), .A2(n41), .ZN(ab_19__12_) );
  NOR2_X1 U473 ( .A1(n27), .A2(n41), .ZN(ab_19__11_) );
  NOR2_X1 U474 ( .A1(n28), .A2(n41), .ZN(ab_19__10_) );
  NOR2_X1 U475 ( .A1(n29), .A2(n41), .ZN(ab_19__0_) );
  NOR2_X1 U476 ( .A1(n7), .A2(n42), .ZN(ab_18__9_) );
  NOR2_X1 U477 ( .A1(n8), .A2(n42), .ZN(ab_18__8_) );
  NOR2_X1 U478 ( .A1(n9), .A2(n42), .ZN(ab_18__7_) );
  NOR2_X1 U479 ( .A1(n10), .A2(n42), .ZN(ab_18__6_) );
  NOR2_X1 U480 ( .A1(n11), .A2(n42), .ZN(ab_18__5_) );
  NOR2_X1 U481 ( .A1(n12), .A2(n42), .ZN(ab_18__4_) );
  NOR2_X1 U482 ( .A1(n13), .A2(n42), .ZN(ab_18__3_) );
  NOR2_X1 U483 ( .A1(n14), .A2(n42), .ZN(ab_18__2_) );
  NOR2_X1 U484 ( .A1(A[18]), .A2(n1), .ZN(ab_18__23_) );
  NOR2_X1 U485 ( .A1(n15), .A2(n42), .ZN(ab_18__22_) );
  NOR2_X1 U486 ( .A1(n16), .A2(n42), .ZN(ab_18__21_) );
  NOR2_X1 U487 ( .A1(n17), .A2(n42), .ZN(ab_18__20_) );
  NOR2_X1 U488 ( .A1(n18), .A2(n42), .ZN(ab_18__1_) );
  NOR2_X1 U489 ( .A1(n19), .A2(n42), .ZN(ab_18__19_) );
  NOR2_X1 U490 ( .A1(n20), .A2(n42), .ZN(ab_18__18_) );
  NOR2_X1 U491 ( .A1(n21), .A2(n42), .ZN(ab_18__17_) );
  NOR2_X1 U492 ( .A1(n22), .A2(n42), .ZN(ab_18__16_) );
  NOR2_X1 U493 ( .A1(n23), .A2(n42), .ZN(ab_18__15_) );
  NOR2_X1 U494 ( .A1(n24), .A2(n42), .ZN(ab_18__14_) );
  NOR2_X1 U495 ( .A1(n25), .A2(n42), .ZN(ab_18__13_) );
  NOR2_X1 U496 ( .A1(n26), .A2(n42), .ZN(ab_18__12_) );
  NOR2_X1 U497 ( .A1(n27), .A2(n42), .ZN(ab_18__11_) );
  NOR2_X1 U498 ( .A1(n28), .A2(n42), .ZN(ab_18__10_) );
  NOR2_X1 U499 ( .A1(n29), .A2(n42), .ZN(ab_18__0_) );
  NOR2_X1 U500 ( .A1(n7), .A2(n43), .ZN(ab_17__9_) );
  NOR2_X1 U501 ( .A1(n8), .A2(n43), .ZN(ab_17__8_) );
  NOR2_X1 U502 ( .A1(n9), .A2(n43), .ZN(ab_17__7_) );
  NOR2_X1 U503 ( .A1(n10), .A2(n43), .ZN(ab_17__6_) );
  NOR2_X1 U504 ( .A1(n11), .A2(n43), .ZN(ab_17__5_) );
  NOR2_X1 U505 ( .A1(n12), .A2(n43), .ZN(ab_17__4_) );
  NOR2_X1 U506 ( .A1(n13), .A2(n43), .ZN(ab_17__3_) );
  NOR2_X1 U507 ( .A1(n14), .A2(n43), .ZN(ab_17__2_) );
  NOR2_X1 U508 ( .A1(A[17]), .A2(n1), .ZN(ab_17__23_) );
  NOR2_X1 U509 ( .A1(n15), .A2(n43), .ZN(ab_17__22_) );
  NOR2_X1 U510 ( .A1(n16), .A2(n43), .ZN(ab_17__21_) );
  NOR2_X1 U511 ( .A1(n17), .A2(n43), .ZN(ab_17__20_) );
  NOR2_X1 U512 ( .A1(n18), .A2(n43), .ZN(ab_17__1_) );
  NOR2_X1 U513 ( .A1(n19), .A2(n43), .ZN(ab_17__19_) );
  NOR2_X1 U514 ( .A1(n20), .A2(n43), .ZN(ab_17__18_) );
  NOR2_X1 U515 ( .A1(n21), .A2(n43), .ZN(ab_17__17_) );
  NOR2_X1 U516 ( .A1(n22), .A2(n43), .ZN(ab_17__16_) );
  NOR2_X1 U517 ( .A1(n23), .A2(n43), .ZN(ab_17__15_) );
  NOR2_X1 U518 ( .A1(n24), .A2(n43), .ZN(ab_17__14_) );
  NOR2_X1 U519 ( .A1(n25), .A2(n43), .ZN(ab_17__13_) );
  NOR2_X1 U520 ( .A1(n26), .A2(n43), .ZN(ab_17__12_) );
  NOR2_X1 U521 ( .A1(n27), .A2(n43), .ZN(ab_17__11_) );
  NOR2_X1 U522 ( .A1(n28), .A2(n43), .ZN(ab_17__10_) );
  NOR2_X1 U523 ( .A1(n29), .A2(n43), .ZN(ab_17__0_) );
  NOR2_X1 U524 ( .A1(n7), .A2(n44), .ZN(ab_16__9_) );
  NOR2_X1 U525 ( .A1(n8), .A2(n44), .ZN(ab_16__8_) );
  NOR2_X1 U526 ( .A1(n9), .A2(n44), .ZN(ab_16__7_) );
  NOR2_X1 U527 ( .A1(n10), .A2(n44), .ZN(ab_16__6_) );
  NOR2_X1 U528 ( .A1(n11), .A2(n44), .ZN(ab_16__5_) );
  NOR2_X1 U529 ( .A1(n12), .A2(n44), .ZN(ab_16__4_) );
  NOR2_X1 U530 ( .A1(n13), .A2(n44), .ZN(ab_16__3_) );
  NOR2_X1 U531 ( .A1(n14), .A2(n44), .ZN(ab_16__2_) );
  NOR2_X1 U532 ( .A1(A[16]), .A2(n1), .ZN(ab_16__23_) );
  NOR2_X1 U533 ( .A1(n15), .A2(n44), .ZN(ab_16__22_) );
  NOR2_X1 U534 ( .A1(n16), .A2(n44), .ZN(ab_16__21_) );
  NOR2_X1 U535 ( .A1(n17), .A2(n44), .ZN(ab_16__20_) );
  NOR2_X1 U536 ( .A1(n18), .A2(n44), .ZN(ab_16__1_) );
  NOR2_X1 U537 ( .A1(n19), .A2(n44), .ZN(ab_16__19_) );
  NOR2_X1 U538 ( .A1(n20), .A2(n44), .ZN(ab_16__18_) );
  NOR2_X1 U539 ( .A1(n21), .A2(n44), .ZN(ab_16__17_) );
  NOR2_X1 U540 ( .A1(n22), .A2(n44), .ZN(ab_16__16_) );
  NOR2_X1 U541 ( .A1(n23), .A2(n44), .ZN(ab_16__15_) );
  NOR2_X1 U542 ( .A1(n24), .A2(n44), .ZN(ab_16__14_) );
  NOR2_X1 U543 ( .A1(n25), .A2(n44), .ZN(ab_16__13_) );
  NOR2_X1 U544 ( .A1(n26), .A2(n44), .ZN(ab_16__12_) );
  NOR2_X1 U545 ( .A1(n27), .A2(n44), .ZN(ab_16__11_) );
  NOR2_X1 U546 ( .A1(n28), .A2(n44), .ZN(ab_16__10_) );
  NOR2_X1 U547 ( .A1(n29), .A2(n44), .ZN(ab_16__0_) );
  NOR2_X1 U548 ( .A1(n7), .A2(n45), .ZN(ab_15__9_) );
  NOR2_X1 U549 ( .A1(n8), .A2(n45), .ZN(ab_15__8_) );
  NOR2_X1 U550 ( .A1(n9), .A2(n45), .ZN(ab_15__7_) );
  NOR2_X1 U551 ( .A1(n10), .A2(n45), .ZN(ab_15__6_) );
  NOR2_X1 U552 ( .A1(n11), .A2(n45), .ZN(ab_15__5_) );
  NOR2_X1 U553 ( .A1(n12), .A2(n45), .ZN(ab_15__4_) );
  NOR2_X1 U554 ( .A1(n13), .A2(n45), .ZN(ab_15__3_) );
  NOR2_X1 U555 ( .A1(n14), .A2(n45), .ZN(ab_15__2_) );
  NOR2_X1 U556 ( .A1(A[15]), .A2(n1), .ZN(ab_15__23_) );
  NOR2_X1 U557 ( .A1(n15), .A2(n45), .ZN(ab_15__22_) );
  NOR2_X1 U558 ( .A1(n16), .A2(n45), .ZN(ab_15__21_) );
  NOR2_X1 U559 ( .A1(n17), .A2(n45), .ZN(ab_15__20_) );
  NOR2_X1 U560 ( .A1(n18), .A2(n45), .ZN(ab_15__1_) );
  NOR2_X1 U561 ( .A1(n19), .A2(n45), .ZN(ab_15__19_) );
  NOR2_X1 U562 ( .A1(n20), .A2(n45), .ZN(ab_15__18_) );
  NOR2_X1 U563 ( .A1(n21), .A2(n45), .ZN(ab_15__17_) );
  NOR2_X1 U564 ( .A1(n22), .A2(n45), .ZN(ab_15__16_) );
  NOR2_X1 U565 ( .A1(n23), .A2(n45), .ZN(ab_15__15_) );
  NOR2_X1 U566 ( .A1(n24), .A2(n45), .ZN(ab_15__14_) );
  NOR2_X1 U567 ( .A1(n25), .A2(n45), .ZN(ab_15__13_) );
  NOR2_X1 U568 ( .A1(n26), .A2(n45), .ZN(ab_15__12_) );
  NOR2_X1 U569 ( .A1(n27), .A2(n45), .ZN(ab_15__11_) );
  NOR2_X1 U570 ( .A1(n28), .A2(n45), .ZN(ab_15__10_) );
  NOR2_X1 U571 ( .A1(n29), .A2(n45), .ZN(ab_15__0_) );
  NOR2_X1 U572 ( .A1(n7), .A2(n46), .ZN(ab_14__9_) );
  NOR2_X1 U573 ( .A1(n8), .A2(n46), .ZN(ab_14__8_) );
  NOR2_X1 U574 ( .A1(n9), .A2(n46), .ZN(ab_14__7_) );
  NOR2_X1 U575 ( .A1(n10), .A2(n46), .ZN(ab_14__6_) );
  NOR2_X1 U576 ( .A1(n11), .A2(n46), .ZN(ab_14__5_) );
  NOR2_X1 U577 ( .A1(n12), .A2(n46), .ZN(ab_14__4_) );
  NOR2_X1 U578 ( .A1(n13), .A2(n46), .ZN(ab_14__3_) );
  NOR2_X1 U579 ( .A1(n14), .A2(n46), .ZN(ab_14__2_) );
  NOR2_X1 U580 ( .A1(A[14]), .A2(n2), .ZN(ab_14__23_) );
  NOR2_X1 U581 ( .A1(n15), .A2(n46), .ZN(ab_14__22_) );
  NOR2_X1 U582 ( .A1(n16), .A2(n46), .ZN(ab_14__21_) );
  NOR2_X1 U583 ( .A1(n17), .A2(n46), .ZN(ab_14__20_) );
  NOR2_X1 U584 ( .A1(n18), .A2(n46), .ZN(ab_14__1_) );
  NOR2_X1 U585 ( .A1(n19), .A2(n46), .ZN(ab_14__19_) );
  NOR2_X1 U586 ( .A1(n20), .A2(n46), .ZN(ab_14__18_) );
  NOR2_X1 U587 ( .A1(n21), .A2(n46), .ZN(ab_14__17_) );
  NOR2_X1 U588 ( .A1(n22), .A2(n46), .ZN(ab_14__16_) );
  NOR2_X1 U589 ( .A1(n23), .A2(n46), .ZN(ab_14__15_) );
  NOR2_X1 U590 ( .A1(n24), .A2(n46), .ZN(ab_14__14_) );
  NOR2_X1 U591 ( .A1(n25), .A2(n46), .ZN(ab_14__13_) );
  NOR2_X1 U592 ( .A1(n26), .A2(n46), .ZN(ab_14__12_) );
  NOR2_X1 U593 ( .A1(n27), .A2(n46), .ZN(ab_14__11_) );
  NOR2_X1 U594 ( .A1(n28), .A2(n46), .ZN(ab_14__10_) );
  NOR2_X1 U595 ( .A1(n29), .A2(n46), .ZN(ab_14__0_) );
  NOR2_X1 U596 ( .A1(n7), .A2(n47), .ZN(ab_13__9_) );
  NOR2_X1 U597 ( .A1(n8), .A2(n47), .ZN(ab_13__8_) );
  NOR2_X1 U598 ( .A1(n9), .A2(n47), .ZN(ab_13__7_) );
  NOR2_X1 U599 ( .A1(n10), .A2(n47), .ZN(ab_13__6_) );
  NOR2_X1 U600 ( .A1(n11), .A2(n47), .ZN(ab_13__5_) );
  NOR2_X1 U601 ( .A1(n12), .A2(n47), .ZN(ab_13__4_) );
  NOR2_X1 U602 ( .A1(n13), .A2(n47), .ZN(ab_13__3_) );
  NOR2_X1 U603 ( .A1(n14), .A2(n47), .ZN(ab_13__2_) );
  NOR2_X1 U604 ( .A1(A[13]), .A2(n2), .ZN(ab_13__23_) );
  NOR2_X1 U605 ( .A1(n15), .A2(n47), .ZN(ab_13__22_) );
  NOR2_X1 U606 ( .A1(n16), .A2(n47), .ZN(ab_13__21_) );
  NOR2_X1 U607 ( .A1(n17), .A2(n47), .ZN(ab_13__20_) );
  NOR2_X1 U608 ( .A1(n18), .A2(n47), .ZN(ab_13__1_) );
  NOR2_X1 U609 ( .A1(n19), .A2(n47), .ZN(ab_13__19_) );
  NOR2_X1 U610 ( .A1(n20), .A2(n47), .ZN(ab_13__18_) );
  NOR2_X1 U611 ( .A1(n21), .A2(n47), .ZN(ab_13__17_) );
  NOR2_X1 U612 ( .A1(n22), .A2(n47), .ZN(ab_13__16_) );
  NOR2_X1 U613 ( .A1(n23), .A2(n47), .ZN(ab_13__15_) );
  NOR2_X1 U614 ( .A1(n24), .A2(n47), .ZN(ab_13__14_) );
  NOR2_X1 U615 ( .A1(n25), .A2(n47), .ZN(ab_13__13_) );
  NOR2_X1 U616 ( .A1(n26), .A2(n47), .ZN(ab_13__12_) );
  NOR2_X1 U617 ( .A1(n27), .A2(n47), .ZN(ab_13__11_) );
  NOR2_X1 U618 ( .A1(n28), .A2(n47), .ZN(ab_13__10_) );
  NOR2_X1 U619 ( .A1(n29), .A2(n47), .ZN(ab_13__0_) );
  NOR2_X1 U620 ( .A1(n7), .A2(n48), .ZN(ab_12__9_) );
  NOR2_X1 U621 ( .A1(n8), .A2(n48), .ZN(ab_12__8_) );
  NOR2_X1 U622 ( .A1(n9), .A2(n48), .ZN(ab_12__7_) );
  NOR2_X1 U623 ( .A1(n10), .A2(n48), .ZN(ab_12__6_) );
  NOR2_X1 U624 ( .A1(n11), .A2(n48), .ZN(ab_12__5_) );
  NOR2_X1 U625 ( .A1(n12), .A2(n48), .ZN(ab_12__4_) );
  NOR2_X1 U626 ( .A1(n13), .A2(n48), .ZN(ab_12__3_) );
  NOR2_X1 U627 ( .A1(n14), .A2(n48), .ZN(ab_12__2_) );
  NOR2_X1 U628 ( .A1(A[12]), .A2(n2), .ZN(ab_12__23_) );
  NOR2_X1 U629 ( .A1(n15), .A2(n48), .ZN(ab_12__22_) );
  NOR2_X1 U630 ( .A1(n16), .A2(n48), .ZN(ab_12__21_) );
  NOR2_X1 U631 ( .A1(n17), .A2(n48), .ZN(ab_12__20_) );
  NOR2_X1 U632 ( .A1(n18), .A2(n48), .ZN(ab_12__1_) );
  NOR2_X1 U633 ( .A1(n19), .A2(n48), .ZN(ab_12__19_) );
  NOR2_X1 U634 ( .A1(n20), .A2(n48), .ZN(ab_12__18_) );
  NOR2_X1 U635 ( .A1(n21), .A2(n48), .ZN(ab_12__17_) );
  NOR2_X1 U636 ( .A1(n22), .A2(n48), .ZN(ab_12__16_) );
  NOR2_X1 U637 ( .A1(n23), .A2(n48), .ZN(ab_12__15_) );
  NOR2_X1 U638 ( .A1(n24), .A2(n48), .ZN(ab_12__14_) );
  NOR2_X1 U639 ( .A1(n25), .A2(n48), .ZN(ab_12__13_) );
  NOR2_X1 U640 ( .A1(n26), .A2(n48), .ZN(ab_12__12_) );
  NOR2_X1 U641 ( .A1(n27), .A2(n48), .ZN(ab_12__11_) );
  NOR2_X1 U642 ( .A1(n28), .A2(n48), .ZN(ab_12__10_) );
  NOR2_X1 U643 ( .A1(n29), .A2(n48), .ZN(ab_12__0_) );
  NOR2_X1 U644 ( .A1(n7), .A2(n49), .ZN(ab_11__9_) );
  NOR2_X1 U645 ( .A1(n8), .A2(n49), .ZN(ab_11__8_) );
  NOR2_X1 U646 ( .A1(n9), .A2(n49), .ZN(ab_11__7_) );
  NOR2_X1 U647 ( .A1(n10), .A2(n49), .ZN(ab_11__6_) );
  NOR2_X1 U648 ( .A1(n11), .A2(n49), .ZN(ab_11__5_) );
  NOR2_X1 U649 ( .A1(n12), .A2(n49), .ZN(ab_11__4_) );
  NOR2_X1 U650 ( .A1(n13), .A2(n49), .ZN(ab_11__3_) );
  NOR2_X1 U651 ( .A1(n14), .A2(n49), .ZN(ab_11__2_) );
  NOR2_X1 U652 ( .A1(A[11]), .A2(n2), .ZN(ab_11__23_) );
  NOR2_X1 U653 ( .A1(n15), .A2(n49), .ZN(ab_11__22_) );
  NOR2_X1 U654 ( .A1(n16), .A2(n49), .ZN(ab_11__21_) );
  NOR2_X1 U655 ( .A1(n17), .A2(n49), .ZN(ab_11__20_) );
  NOR2_X1 U656 ( .A1(n18), .A2(n49), .ZN(ab_11__1_) );
  NOR2_X1 U657 ( .A1(n19), .A2(n49), .ZN(ab_11__19_) );
  NOR2_X1 U658 ( .A1(n20), .A2(n49), .ZN(ab_11__18_) );
  NOR2_X1 U659 ( .A1(n21), .A2(n49), .ZN(ab_11__17_) );
  NOR2_X1 U660 ( .A1(n22), .A2(n49), .ZN(ab_11__16_) );
  NOR2_X1 U661 ( .A1(n23), .A2(n49), .ZN(ab_11__15_) );
  NOR2_X1 U662 ( .A1(n24), .A2(n49), .ZN(ab_11__14_) );
  NOR2_X1 U663 ( .A1(n25), .A2(n49), .ZN(ab_11__13_) );
  NOR2_X1 U664 ( .A1(n26), .A2(n49), .ZN(ab_11__12_) );
  NOR2_X1 U665 ( .A1(n27), .A2(n49), .ZN(ab_11__11_) );
  NOR2_X1 U666 ( .A1(n28), .A2(n49), .ZN(ab_11__10_) );
  NOR2_X1 U667 ( .A1(n29), .A2(n49), .ZN(ab_11__0_) );
  NOR2_X1 U668 ( .A1(n7), .A2(n50), .ZN(ab_10__9_) );
  NOR2_X1 U669 ( .A1(n8), .A2(n50), .ZN(ab_10__8_) );
  NOR2_X1 U670 ( .A1(n9), .A2(n50), .ZN(ab_10__7_) );
  NOR2_X1 U671 ( .A1(n10), .A2(n50), .ZN(ab_10__6_) );
  NOR2_X1 U672 ( .A1(n11), .A2(n50), .ZN(ab_10__5_) );
  NOR2_X1 U673 ( .A1(n12), .A2(n50), .ZN(ab_10__4_) );
  NOR2_X1 U674 ( .A1(n13), .A2(n50), .ZN(ab_10__3_) );
  NOR2_X1 U675 ( .A1(n14), .A2(n50), .ZN(ab_10__2_) );
  NOR2_X1 U676 ( .A1(A[10]), .A2(n2), .ZN(ab_10__23_) );
  NOR2_X1 U677 ( .A1(n15), .A2(n50), .ZN(ab_10__22_) );
  NOR2_X1 U678 ( .A1(n16), .A2(n50), .ZN(ab_10__21_) );
  NOR2_X1 U679 ( .A1(n17), .A2(n50), .ZN(ab_10__20_) );
  NOR2_X1 U680 ( .A1(n18), .A2(n50), .ZN(ab_10__1_) );
  NOR2_X1 U681 ( .A1(n19), .A2(n50), .ZN(ab_10__19_) );
  NOR2_X1 U682 ( .A1(n20), .A2(n50), .ZN(ab_10__18_) );
  NOR2_X1 U683 ( .A1(n21), .A2(n50), .ZN(ab_10__17_) );
  NOR2_X1 U684 ( .A1(n22), .A2(n50), .ZN(ab_10__16_) );
  NOR2_X1 U685 ( .A1(n23), .A2(n50), .ZN(ab_10__15_) );
  NOR2_X1 U686 ( .A1(n24), .A2(n50), .ZN(ab_10__14_) );
  NOR2_X1 U687 ( .A1(n25), .A2(n50), .ZN(ab_10__13_) );
  NOR2_X1 U688 ( .A1(n26), .A2(n50), .ZN(ab_10__12_) );
  NOR2_X1 U689 ( .A1(n27), .A2(n50), .ZN(ab_10__11_) );
  NOR2_X1 U690 ( .A1(n28), .A2(n50), .ZN(ab_10__10_) );
  NOR2_X1 U691 ( .A1(n29), .A2(n50), .ZN(ab_10__0_) );
  NOR2_X1 U692 ( .A1(n7), .A2(n51), .ZN(ab_0__9_) );
  NOR2_X1 U693 ( .A1(n8), .A2(n51), .ZN(ab_0__8_) );
  NOR2_X1 U694 ( .A1(n9), .A2(n51), .ZN(ab_0__7_) );
  NOR2_X1 U695 ( .A1(n10), .A2(n51), .ZN(ab_0__6_) );
  NOR2_X1 U696 ( .A1(n11), .A2(n51), .ZN(ab_0__5_) );
  NOR2_X1 U697 ( .A1(n12), .A2(n51), .ZN(ab_0__4_) );
  NOR2_X1 U698 ( .A1(n13), .A2(n51), .ZN(ab_0__3_) );
  NOR2_X1 U699 ( .A1(n14), .A2(n51), .ZN(ab_0__2_) );
  NOR2_X1 U700 ( .A1(A[0]), .A2(n1), .ZN(ab_0__23_) );
  NOR2_X1 U701 ( .A1(n15), .A2(n51), .ZN(ab_0__22_) );
  NOR2_X1 U702 ( .A1(n16), .A2(n51), .ZN(ab_0__21_) );
  NOR2_X1 U703 ( .A1(n17), .A2(n51), .ZN(ab_0__20_) );
  NOR2_X1 U704 ( .A1(n19), .A2(n51), .ZN(ab_0__19_) );
  NOR2_X1 U705 ( .A1(n20), .A2(n51), .ZN(ab_0__18_) );
  NOR2_X1 U706 ( .A1(n21), .A2(n51), .ZN(ab_0__17_) );
  NOR2_X1 U707 ( .A1(n22), .A2(n51), .ZN(ab_0__16_) );
  NOR2_X1 U708 ( .A1(n23), .A2(n51), .ZN(ab_0__15_) );
  NOR2_X1 U709 ( .A1(n24), .A2(n51), .ZN(ab_0__14_) );
  NOR2_X1 U710 ( .A1(n25), .A2(n51), .ZN(ab_0__13_) );
  NOR2_X1 U711 ( .A1(n26), .A2(n51), .ZN(ab_0__12_) );
  NOR2_X1 U712 ( .A1(n27), .A2(n51), .ZN(ab_0__11_) );
  NOR2_X1 U713 ( .A1(n28), .A2(n51), .ZN(ab_0__10_) );
  INV_X1 U714 ( .A(B[23]), .ZN(QB) );
  INV_X1 U715 ( .A(A[23]), .ZN(QA) );
  AND3_X1 U716 ( .A1(ab_1__1_), .A2(B[0]), .A3(A[0]), .ZN(CARRYB_1__0_) );
  NOR2_X1 U717 ( .A1(n40), .A2(n18), .ZN(ab_1__1_) );
  INV_X1 U719 ( .A(CARRYB_23__23_), .ZN(A1_45_) );
endmodule


module iir_filter_DW01_add_5 ( A, B, CI, SUM, CO );
  input [45:0] A;
  input [45:0] B;
  output [45:0] SUM;
  input CI;
  output CO;
  wire   A_21_, A_20_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112;
  assign SUM[21] = A_21_;
  assign A_21_ = A[21];
  assign SUM[20] = A_20_;
  assign A_20_ = A[20];

  XOR2_X1 U2 ( .A(n1), .B(n2), .Z(SUM[45]) );
  XOR2_X1 U3 ( .A(B[45]), .B(A[45]), .Z(n2) );
  OAI21_X1 U4 ( .B1(n3), .B2(n4), .A(n5), .ZN(n1) );
  OAI21_X1 U5 ( .B1(A[44]), .B2(n6), .A(B[44]), .ZN(n5) );
  INV_X1 U6 ( .A(n3), .ZN(n6) );
  INV_X1 U7 ( .A(A[44]), .ZN(n4) );
  AOI21_X1 U8 ( .B1(A[43]), .B2(B[43]), .A(n7), .ZN(n3) );
  INV_X1 U9 ( .A(n8), .ZN(n7) );
  OAI22_X1 U10 ( .A1(n9), .A2(n10), .B1(A[43]), .B2(B[43]), .ZN(n8) );
  AOI21_X1 U11 ( .B1(n11), .B2(n12), .A(n13), .ZN(n9) );
  NAND3_X1 U12 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n12) );
  AOI21_X1 U13 ( .B1(n17), .B2(n16), .A(n18), .ZN(n11) );
  INV_X1 U14 ( .A(n19), .ZN(n18) );
  XOR2_X1 U15 ( .A(n20), .B(n21), .Z(SUM[42]) );
  NOR2_X1 U16 ( .A1(n10), .A2(n13), .ZN(n21) );
  NOR2_X1 U17 ( .A1(B[42]), .A2(A[42]), .ZN(n13) );
  AND2_X1 U18 ( .A1(B[42]), .A2(A[42]), .ZN(n10) );
  OAI21_X1 U19 ( .B1(n22), .B2(n23), .A(n19), .ZN(n20) );
  XOR2_X1 U20 ( .A(n24), .B(n23), .Z(SUM[41]) );
  AOI21_X1 U21 ( .B1(n15), .B2(n14), .A(n17), .ZN(n23) );
  INV_X1 U22 ( .A(n25), .ZN(n15) );
  NAND2_X1 U23 ( .A1(n16), .A2(n19), .ZN(n24) );
  NAND2_X1 U24 ( .A1(B[41]), .A2(A[41]), .ZN(n19) );
  INV_X1 U25 ( .A(n22), .ZN(n16) );
  NOR2_X1 U26 ( .A1(B[41]), .A2(A[41]), .ZN(n22) );
  XOR2_X1 U27 ( .A(n14), .B(n26), .Z(SUM[40]) );
  NOR2_X1 U28 ( .A1(n17), .A2(n25), .ZN(n26) );
  NOR2_X1 U29 ( .A1(B[40]), .A2(A[40]), .ZN(n25) );
  AND2_X1 U30 ( .A1(B[40]), .A2(A[40]), .ZN(n17) );
  OAI21_X1 U31 ( .B1(n27), .B2(n28), .A(n29), .ZN(n14) );
  XOR2_X1 U32 ( .A(n30), .B(n28), .Z(SUM[39]) );
  AOI21_X1 U33 ( .B1(n31), .B2(n32), .A(n33), .ZN(n28) );
  INV_X1 U34 ( .A(n34), .ZN(n31) );
  NAND2_X1 U35 ( .A1(n35), .A2(n29), .ZN(n30) );
  NAND2_X1 U36 ( .A1(B[39]), .A2(A[39]), .ZN(n29) );
  INV_X1 U37 ( .A(n27), .ZN(n35) );
  NOR2_X1 U38 ( .A1(B[39]), .A2(A[39]), .ZN(n27) );
  XOR2_X1 U39 ( .A(n32), .B(n36), .Z(SUM[38]) );
  NOR2_X1 U40 ( .A1(n33), .A2(n34), .ZN(n36) );
  NOR2_X1 U41 ( .A1(B[38]), .A2(A[38]), .ZN(n34) );
  AND2_X1 U42 ( .A1(B[38]), .A2(A[38]), .ZN(n33) );
  OAI21_X1 U43 ( .B1(n37), .B2(n38), .A(n39), .ZN(n32) );
  XOR2_X1 U44 ( .A(n40), .B(n38), .Z(SUM[37]) );
  AOI21_X1 U45 ( .B1(n41), .B2(n42), .A(n43), .ZN(n38) );
  INV_X1 U46 ( .A(n44), .ZN(n41) );
  NAND2_X1 U47 ( .A1(n45), .A2(n39), .ZN(n40) );
  NAND2_X1 U48 ( .A1(B[37]), .A2(A[37]), .ZN(n39) );
  INV_X1 U49 ( .A(n37), .ZN(n45) );
  NOR2_X1 U50 ( .A1(B[37]), .A2(A[37]), .ZN(n37) );
  XOR2_X1 U51 ( .A(n42), .B(n46), .Z(SUM[36]) );
  NOR2_X1 U52 ( .A1(n43), .A2(n44), .ZN(n46) );
  NOR2_X1 U53 ( .A1(B[36]), .A2(A[36]), .ZN(n44) );
  AND2_X1 U54 ( .A1(B[36]), .A2(A[36]), .ZN(n43) );
  OAI21_X1 U55 ( .B1(n47), .B2(n48), .A(n49), .ZN(n42) );
  XOR2_X1 U56 ( .A(n50), .B(n48), .Z(SUM[35]) );
  AOI21_X1 U57 ( .B1(n51), .B2(n52), .A(n53), .ZN(n48) );
  INV_X1 U58 ( .A(n54), .ZN(n51) );
  NAND2_X1 U59 ( .A1(n55), .A2(n49), .ZN(n50) );
  NAND2_X1 U60 ( .A1(B[35]), .A2(A[35]), .ZN(n49) );
  INV_X1 U61 ( .A(n47), .ZN(n55) );
  NOR2_X1 U62 ( .A1(B[35]), .A2(A[35]), .ZN(n47) );
  XOR2_X1 U63 ( .A(n52), .B(n56), .Z(SUM[34]) );
  NOR2_X1 U64 ( .A1(n53), .A2(n54), .ZN(n56) );
  NOR2_X1 U65 ( .A1(B[34]), .A2(A[34]), .ZN(n54) );
  AND2_X1 U66 ( .A1(B[34]), .A2(A[34]), .ZN(n53) );
  OAI21_X1 U67 ( .B1(n57), .B2(n58), .A(n59), .ZN(n52) );
  XOR2_X1 U68 ( .A(n60), .B(n58), .Z(SUM[33]) );
  AOI21_X1 U69 ( .B1(n61), .B2(n62), .A(n63), .ZN(n58) );
  INV_X1 U70 ( .A(n64), .ZN(n61) );
  NAND2_X1 U71 ( .A1(n65), .A2(n59), .ZN(n60) );
  NAND2_X1 U72 ( .A1(B[33]), .A2(A[33]), .ZN(n59) );
  INV_X1 U73 ( .A(n57), .ZN(n65) );
  NOR2_X1 U74 ( .A1(B[33]), .A2(A[33]), .ZN(n57) );
  XOR2_X1 U75 ( .A(n62), .B(n66), .Z(SUM[32]) );
  NOR2_X1 U76 ( .A1(n63), .A2(n64), .ZN(n66) );
  NOR2_X1 U77 ( .A1(B[32]), .A2(A[32]), .ZN(n64) );
  AND2_X1 U78 ( .A1(B[32]), .A2(A[32]), .ZN(n63) );
  OAI21_X1 U79 ( .B1(n67), .B2(n68), .A(n69), .ZN(n62) );
  XOR2_X1 U80 ( .A(n70), .B(n68), .Z(SUM[31]) );
  AOI21_X1 U81 ( .B1(n71), .B2(n72), .A(n73), .ZN(n68) );
  INV_X1 U82 ( .A(n74), .ZN(n71) );
  NAND2_X1 U83 ( .A1(n75), .A2(n69), .ZN(n70) );
  NAND2_X1 U84 ( .A1(B[31]), .A2(A[31]), .ZN(n69) );
  INV_X1 U85 ( .A(n67), .ZN(n75) );
  NOR2_X1 U86 ( .A1(B[31]), .A2(A[31]), .ZN(n67) );
  XOR2_X1 U87 ( .A(n72), .B(n76), .Z(SUM[30]) );
  NOR2_X1 U88 ( .A1(n73), .A2(n74), .ZN(n76) );
  NOR2_X1 U89 ( .A1(B[30]), .A2(A[30]), .ZN(n74) );
  AND2_X1 U90 ( .A1(B[30]), .A2(A[30]), .ZN(n73) );
  OAI21_X1 U91 ( .B1(n77), .B2(n78), .A(n79), .ZN(n72) );
  XOR2_X1 U92 ( .A(n80), .B(n78), .Z(SUM[29]) );
  AOI21_X1 U93 ( .B1(n81), .B2(n82), .A(n83), .ZN(n78) );
  INV_X1 U94 ( .A(n84), .ZN(n81) );
  NAND2_X1 U95 ( .A1(n85), .A2(n79), .ZN(n80) );
  NAND2_X1 U96 ( .A1(B[29]), .A2(A[29]), .ZN(n79) );
  INV_X1 U97 ( .A(n77), .ZN(n85) );
  NOR2_X1 U98 ( .A1(B[29]), .A2(A[29]), .ZN(n77) );
  XOR2_X1 U99 ( .A(n82), .B(n86), .Z(SUM[28]) );
  NOR2_X1 U100 ( .A1(n83), .A2(n84), .ZN(n86) );
  NOR2_X1 U101 ( .A1(B[28]), .A2(A[28]), .ZN(n84) );
  AND2_X1 U102 ( .A1(B[28]), .A2(A[28]), .ZN(n83) );
  OAI21_X1 U103 ( .B1(n87), .B2(n88), .A(n89), .ZN(n82) );
  XOR2_X1 U104 ( .A(n90), .B(n88), .Z(SUM[27]) );
  AOI21_X1 U105 ( .B1(n91), .B2(n92), .A(n93), .ZN(n88) );
  INV_X1 U106 ( .A(n94), .ZN(n92) );
  NAND2_X1 U107 ( .A1(n95), .A2(n89), .ZN(n90) );
  NAND2_X1 U108 ( .A1(B[27]), .A2(A[27]), .ZN(n89) );
  INV_X1 U109 ( .A(n87), .ZN(n95) );
  NOR2_X1 U110 ( .A1(B[27]), .A2(A[27]), .ZN(n87) );
  XOR2_X1 U111 ( .A(n91), .B(n96), .Z(SUM[26]) );
  NOR2_X1 U112 ( .A1(n93), .A2(n94), .ZN(n96) );
  NOR2_X1 U113 ( .A1(B[26]), .A2(A[26]), .ZN(n94) );
  AND2_X1 U114 ( .A1(B[26]), .A2(A[26]), .ZN(n93) );
  OAI21_X1 U115 ( .B1(n97), .B2(n98), .A(n99), .ZN(n91) );
  XOR2_X1 U116 ( .A(n100), .B(n98), .Z(SUM[25]) );
  AOI21_X1 U117 ( .B1(n101), .B2(n102), .A(n103), .ZN(n98) );
  INV_X1 U118 ( .A(n104), .ZN(n101) );
  NAND2_X1 U119 ( .A1(n105), .A2(n99), .ZN(n100) );
  NAND2_X1 U120 ( .A1(B[25]), .A2(A[25]), .ZN(n99) );
  INV_X1 U121 ( .A(n97), .ZN(n105) );
  NOR2_X1 U122 ( .A1(B[25]), .A2(A[25]), .ZN(n97) );
  XOR2_X1 U123 ( .A(n102), .B(n106), .Z(SUM[24]) );
  NOR2_X1 U124 ( .A1(n103), .A2(n104), .ZN(n106) );
  NOR2_X1 U125 ( .A1(B[24]), .A2(A[24]), .ZN(n104) );
  AND2_X1 U126 ( .A1(B[24]), .A2(A[24]), .ZN(n103) );
  OAI21_X1 U127 ( .B1(n107), .B2(n108), .A(n109), .ZN(n102) );
  XOR2_X1 U128 ( .A(n108), .B(n110), .Z(SUM[23]) );
  NAND2_X1 U129 ( .A1(n111), .A2(n109), .ZN(n110) );
  NAND2_X1 U130 ( .A1(B[23]), .A2(A[23]), .ZN(n109) );
  INV_X1 U131 ( .A(n107), .ZN(n111) );
  NOR2_X1 U132 ( .A1(B[23]), .A2(A[23]), .ZN(n107) );
  INV_X1 U133 ( .A(n112), .ZN(SUM[22]) );
  OAI21_X1 U134 ( .B1(B[22]), .B2(A[22]), .A(n108), .ZN(n112) );
  NAND2_X1 U135 ( .A1(B[22]), .A2(A[22]), .ZN(n108) );
endmodule


module iir_filter_DW02_mult_1 ( A, B, TC, PRODUCT );
  input [23:0] A;
  input [23:0] B;
  output [47:0] PRODUCT;
  input TC;
  wire   ab_23__23_, ab_23__22_, ab_23__21_, ab_23__20_, ab_23__19_,
         ab_23__18_, ab_23__17_, ab_23__16_, ab_23__15_, ab_23__14_,
         ab_23__13_, ab_23__12_, ab_23__11_, ab_23__10_, ab_23__9_, ab_23__8_,
         ab_23__7_, ab_23__6_, ab_23__5_, ab_23__4_, ab_23__3_, ab_23__2_,
         ab_23__1_, ab_23__0_, ab_22__23_, ab_22__22_, ab_22__21_, ab_22__20_,
         ab_22__19_, ab_22__18_, ab_22__17_, ab_22__16_, ab_22__15_,
         ab_22__14_, ab_22__13_, ab_22__12_, ab_22__11_, ab_22__10_, ab_22__9_,
         ab_22__8_, ab_22__7_, ab_22__6_, ab_22__5_, ab_22__4_, ab_22__3_,
         ab_22__2_, ab_22__1_, ab_22__0_, ab_21__23_, ab_21__22_, ab_21__21_,
         ab_21__20_, ab_21__19_, ab_21__18_, ab_21__17_, ab_21__16_,
         ab_21__15_, ab_21__14_, ab_21__13_, ab_21__12_, ab_21__11_,
         ab_21__10_, ab_21__9_, ab_21__8_, ab_21__7_, ab_21__6_, ab_21__5_,
         ab_21__4_, ab_21__3_, ab_21__2_, ab_21__1_, ab_21__0_, ab_20__23_,
         ab_20__22_, ab_20__21_, ab_20__20_, ab_20__19_, ab_20__18_,
         ab_20__17_, ab_20__16_, ab_20__15_, ab_20__14_, ab_20__13_,
         ab_20__12_, ab_20__11_, ab_20__10_, ab_20__9_, ab_20__8_, ab_20__7_,
         ab_20__6_, ab_20__5_, ab_20__4_, ab_20__3_, ab_20__2_, ab_20__1_,
         ab_20__0_, ab_19__23_, ab_19__22_, ab_19__21_, ab_19__20_, ab_19__19_,
         ab_19__18_, ab_19__17_, ab_19__16_, ab_19__15_, ab_19__14_,
         ab_19__13_, ab_19__12_, ab_19__11_, ab_19__10_, ab_19__9_, ab_19__8_,
         ab_19__7_, ab_19__6_, ab_19__5_, ab_19__4_, ab_19__3_, ab_19__2_,
         ab_19__1_, ab_19__0_, ab_18__23_, ab_18__22_, ab_18__21_, ab_18__20_,
         ab_18__19_, ab_18__18_, ab_18__17_, ab_18__16_, ab_18__15_,
         ab_18__14_, ab_18__13_, ab_18__12_, ab_18__11_, ab_18__10_, ab_18__9_,
         ab_18__8_, ab_18__7_, ab_18__6_, ab_18__5_, ab_18__4_, ab_18__3_,
         ab_18__2_, ab_18__1_, ab_18__0_, ab_17__23_, ab_17__22_, ab_17__21_,
         ab_17__20_, ab_17__19_, ab_17__18_, ab_17__17_, ab_17__16_,
         ab_17__15_, ab_17__14_, ab_17__13_, ab_17__12_, ab_17__11_,
         ab_17__10_, ab_17__9_, ab_17__8_, ab_17__7_, ab_17__6_, ab_17__5_,
         ab_17__4_, ab_17__3_, ab_17__2_, ab_17__1_, ab_17__0_, ab_16__23_,
         ab_16__22_, ab_16__21_, ab_16__20_, ab_16__19_, ab_16__18_,
         ab_16__17_, ab_16__16_, ab_16__15_, ab_16__14_, ab_16__13_,
         ab_16__12_, ab_16__11_, ab_16__10_, ab_16__9_, ab_16__8_, ab_16__7_,
         ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_, ab_16__1_,
         ab_16__0_, ab_15__23_, ab_15__22_, ab_15__21_, ab_15__20_, ab_15__19_,
         ab_15__18_, ab_15__17_, ab_15__16_, ab_15__15_, ab_15__14_,
         ab_15__13_, ab_15__12_, ab_15__11_, ab_15__10_, ab_15__9_, ab_15__8_,
         ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_, ab_15__3_, ab_15__2_,
         ab_15__1_, ab_15__0_, ab_14__23_, ab_14__22_, ab_14__21_, ab_14__20_,
         ab_14__19_, ab_14__18_, ab_14__17_, ab_14__16_, ab_14__15_,
         ab_14__14_, ab_14__13_, ab_14__12_, ab_14__11_, ab_14__10_, ab_14__9_,
         ab_14__8_, ab_14__7_, ab_14__6_, ab_14__5_, ab_14__4_, ab_14__3_,
         ab_14__2_, ab_14__1_, ab_14__0_, ab_13__23_, ab_13__22_, ab_13__21_,
         ab_13__20_, ab_13__19_, ab_13__18_, ab_13__17_, ab_13__16_,
         ab_13__15_, ab_13__14_, ab_13__13_, ab_13__12_, ab_13__11_,
         ab_13__10_, ab_13__9_, ab_13__8_, ab_13__7_, ab_13__6_, ab_13__5_,
         ab_13__4_, ab_13__3_, ab_13__2_, ab_13__1_, ab_13__0_, ab_12__23_,
         ab_12__22_, ab_12__21_, ab_12__20_, ab_12__19_, ab_12__18_,
         ab_12__17_, ab_12__16_, ab_12__15_, ab_12__14_, ab_12__13_,
         ab_12__12_, ab_12__11_, ab_12__10_, ab_12__9_, ab_12__8_, ab_12__7_,
         ab_12__6_, ab_12__5_, ab_12__4_, ab_12__3_, ab_12__2_, ab_12__1_,
         ab_12__0_, ab_11__23_, ab_11__22_, ab_11__21_, ab_11__20_, ab_11__19_,
         ab_11__18_, ab_11__17_, ab_11__16_, ab_11__15_, ab_11__14_,
         ab_11__13_, ab_11__12_, ab_11__11_, ab_11__10_, ab_11__9_, ab_11__8_,
         ab_11__7_, ab_11__6_, ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_,
         ab_11__1_, ab_11__0_, ab_10__23_, ab_10__22_, ab_10__21_, ab_10__20_,
         ab_10__19_, ab_10__18_, ab_10__17_, ab_10__16_, ab_10__15_,
         ab_10__14_, ab_10__13_, ab_10__12_, ab_10__11_, ab_10__10_, ab_10__9_,
         ab_10__8_, ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_,
         ab_10__2_, ab_10__1_, ab_10__0_, ab_9__23_, ab_9__22_, ab_9__21_,
         ab_9__20_, ab_9__19_, ab_9__18_, ab_9__17_, ab_9__16_, ab_9__15_,
         ab_9__14_, ab_9__13_, ab_9__12_, ab_9__11_, ab_9__10_, ab_9__9_,
         ab_9__8_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_,
         ab_9__1_, ab_9__0_, ab_8__23_, ab_8__22_, ab_8__21_, ab_8__20_,
         ab_8__19_, ab_8__18_, ab_8__17_, ab_8__16_, ab_8__15_, ab_8__14_,
         ab_8__13_, ab_8__12_, ab_8__11_, ab_8__10_, ab_8__9_, ab_8__8_,
         ab_8__7_, ab_8__6_, ab_8__5_, ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_,
         ab_8__0_, ab_7__23_, ab_7__22_, ab_7__21_, ab_7__20_, ab_7__19_,
         ab_7__18_, ab_7__17_, ab_7__16_, ab_7__15_, ab_7__14_, ab_7__13_,
         ab_7__12_, ab_7__11_, ab_7__10_, ab_7__9_, ab_7__8_, ab_7__7_,
         ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_,
         ab_6__23_, ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_, ab_6__18_,
         ab_6__17_, ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_, ab_6__12_,
         ab_6__11_, ab_6__10_, ab_6__9_, ab_6__8_, ab_6__7_, ab_6__6_,
         ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_, ab_5__23_,
         ab_5__22_, ab_5__21_, ab_5__20_, ab_5__19_, ab_5__18_, ab_5__17_,
         ab_5__16_, ab_5__15_, ab_5__14_, ab_5__13_, ab_5__12_, ab_5__11_,
         ab_5__10_, ab_5__9_, ab_5__8_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_,
         ab_5__3_, ab_5__2_, ab_5__1_, ab_5__0_, ab_4__23_, ab_4__22_,
         ab_4__21_, ab_4__20_, ab_4__19_, ab_4__18_, ab_4__17_, ab_4__16_,
         ab_4__15_, ab_4__14_, ab_4__13_, ab_4__12_, ab_4__11_, ab_4__10_,
         ab_4__9_, ab_4__8_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_,
         ab_4__2_, ab_4__1_, ab_4__0_, ab_3__23_, ab_3__22_, ab_3__21_,
         ab_3__20_, ab_3__19_, ab_3__18_, ab_3__17_, ab_3__16_, ab_3__15_,
         ab_3__14_, ab_3__13_, ab_3__12_, ab_3__11_, ab_3__10_, ab_3__9_,
         ab_3__8_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_, ab_3__2_,
         ab_3__1_, ab_3__0_, ab_2__23_, ab_2__22_, ab_2__21_, ab_2__20_,
         ab_2__19_, ab_2__18_, ab_2__17_, ab_2__16_, ab_2__15_, ab_2__14_,
         ab_2__13_, ab_2__12_, ab_2__11_, ab_2__10_, ab_2__9_, ab_2__8_,
         ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_,
         ab_2__0_, ab_1__23_, ab_1__22_, ab_1__21_, ab_1__20_, ab_1__19_,
         ab_1__18_, ab_1__17_, ab_1__16_, ab_1__15_, ab_1__14_, ab_1__13_,
         ab_1__12_, ab_1__11_, ab_1__10_, ab_1__9_, ab_1__8_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_0__23_,
         ab_0__22_, ab_0__21_, ab_0__20_, ab_0__19_, ab_0__18_, ab_0__17_,
         ab_0__16_, ab_0__15_, ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_,
         ab_0__10_, ab_0__9_, ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_23__23_, CARRYB_23__22_, CARRYB_23__21_,
         CARRYB_23__20_, CARRYB_23__19_, CARRYB_23__18_, CARRYB_23__17_,
         CARRYB_23__16_, CARRYB_23__15_, CARRYB_23__14_, CARRYB_23__13_,
         CARRYB_23__12_, CARRYB_23__11_, CARRYB_23__10_, CARRYB_23__9_,
         CARRYB_23__8_, CARRYB_23__7_, CARRYB_23__6_, CARRYB_23__5_,
         CARRYB_23__4_, CARRYB_23__3_, CARRYB_23__2_, CARRYB_23__1_,
         CARRYB_23__0_, CARRYB_22__22_, CARRYB_22__21_, CARRYB_22__20_,
         CARRYB_22__19_, CARRYB_22__18_, CARRYB_22__17_, CARRYB_22__16_,
         CARRYB_22__15_, CARRYB_22__14_, CARRYB_22__13_, CARRYB_22__12_,
         CARRYB_22__11_, CARRYB_22__10_, CARRYB_22__9_, CARRYB_22__8_,
         CARRYB_22__7_, CARRYB_22__6_, CARRYB_22__5_, CARRYB_22__4_,
         CARRYB_22__3_, CARRYB_22__2_, CARRYB_22__1_, CARRYB_22__0_,
         CARRYB_21__22_, CARRYB_21__21_, CARRYB_21__20_, CARRYB_21__19_,
         CARRYB_21__18_, CARRYB_21__17_, CARRYB_21__16_, CARRYB_21__15_,
         CARRYB_21__14_, CARRYB_21__13_, CARRYB_21__12_, CARRYB_21__11_,
         CARRYB_21__10_, CARRYB_21__9_, CARRYB_21__8_, CARRYB_21__7_,
         CARRYB_21__6_, CARRYB_21__5_, CARRYB_21__4_, CARRYB_21__3_,
         CARRYB_21__2_, CARRYB_21__1_, CARRYB_21__0_, CARRYB_20__22_,
         CARRYB_20__21_, CARRYB_20__20_, CARRYB_20__19_, CARRYB_20__18_,
         CARRYB_20__17_, CARRYB_20__16_, CARRYB_20__15_, CARRYB_20__14_,
         CARRYB_20__13_, CARRYB_20__12_, CARRYB_20__11_, CARRYB_20__10_,
         CARRYB_20__9_, CARRYB_20__8_, CARRYB_20__7_, CARRYB_20__6_,
         CARRYB_20__5_, CARRYB_20__4_, CARRYB_20__3_, CARRYB_20__2_,
         CARRYB_20__1_, CARRYB_20__0_, CARRYB_19__22_, CARRYB_19__21_,
         CARRYB_19__20_, CARRYB_19__19_, CARRYB_19__18_, CARRYB_19__17_,
         CARRYB_19__16_, CARRYB_19__15_, CARRYB_19__14_, CARRYB_19__13_,
         CARRYB_19__12_, CARRYB_19__11_, CARRYB_19__10_, CARRYB_19__9_,
         CARRYB_19__8_, CARRYB_19__7_, CARRYB_19__6_, CARRYB_19__5_,
         CARRYB_19__4_, CARRYB_19__3_, CARRYB_19__2_, CARRYB_19__1_,
         CARRYB_19__0_, CARRYB_18__22_, CARRYB_18__21_, CARRYB_18__20_,
         CARRYB_18__19_, CARRYB_18__18_, CARRYB_18__17_, CARRYB_18__16_,
         CARRYB_18__15_, CARRYB_18__14_, CARRYB_18__13_, CARRYB_18__12_,
         CARRYB_18__11_, CARRYB_18__10_, CARRYB_18__9_, CARRYB_18__8_,
         CARRYB_18__7_, CARRYB_18__6_, CARRYB_18__5_, CARRYB_18__4_,
         CARRYB_18__3_, CARRYB_18__2_, CARRYB_18__1_, CARRYB_18__0_,
         CARRYB_17__22_, CARRYB_17__21_, CARRYB_17__20_, CARRYB_17__19_,
         CARRYB_17__18_, CARRYB_17__17_, CARRYB_17__16_, CARRYB_17__15_,
         CARRYB_17__14_, CARRYB_17__13_, CARRYB_17__12_, CARRYB_17__11_,
         CARRYB_17__10_, CARRYB_17__9_, CARRYB_17__8_, CARRYB_17__7_,
         CARRYB_17__6_, CARRYB_17__5_, CARRYB_17__4_, CARRYB_17__3_,
         CARRYB_17__2_, CARRYB_17__1_, CARRYB_17__0_, CARRYB_16__22_,
         CARRYB_16__21_, CARRYB_16__20_, CARRYB_16__19_, CARRYB_16__18_,
         CARRYB_16__17_, CARRYB_16__16_, CARRYB_16__15_, CARRYB_16__14_,
         CARRYB_16__13_, CARRYB_16__12_, CARRYB_16__11_, CARRYB_16__10_,
         CARRYB_16__9_, CARRYB_16__8_, CARRYB_16__7_, CARRYB_16__6_,
         CARRYB_16__5_, CARRYB_16__4_, CARRYB_16__3_, CARRYB_16__2_,
         CARRYB_16__1_, CARRYB_16__0_, CARRYB_15__22_, CARRYB_15__21_,
         CARRYB_15__20_, CARRYB_15__19_, CARRYB_15__18_, CARRYB_15__17_,
         CARRYB_15__16_, CARRYB_15__15_, CARRYB_15__14_, CARRYB_15__13_,
         CARRYB_15__12_, CARRYB_15__11_, CARRYB_15__10_, CARRYB_15__9_,
         CARRYB_15__8_, CARRYB_15__7_, CARRYB_15__6_, CARRYB_15__5_,
         CARRYB_15__4_, CARRYB_15__3_, CARRYB_15__2_, CARRYB_15__1_,
         CARRYB_15__0_, CARRYB_14__22_, CARRYB_14__21_, CARRYB_14__20_,
         CARRYB_14__19_, CARRYB_14__18_, CARRYB_14__17_, CARRYB_14__16_,
         CARRYB_14__15_, CARRYB_14__14_, CARRYB_14__13_, CARRYB_14__12_,
         CARRYB_14__11_, CARRYB_14__10_, CARRYB_14__9_, CARRYB_14__8_,
         CARRYB_14__7_, CARRYB_14__6_, CARRYB_14__5_, CARRYB_14__4_,
         CARRYB_14__3_, CARRYB_14__2_, CARRYB_14__1_, CARRYB_14__0_,
         CARRYB_13__22_, CARRYB_13__21_, CARRYB_13__20_, CARRYB_13__19_,
         CARRYB_13__18_, CARRYB_13__17_, CARRYB_13__16_, CARRYB_13__15_,
         CARRYB_13__14_, CARRYB_13__13_, CARRYB_13__12_, CARRYB_13__11_,
         CARRYB_13__10_, CARRYB_13__9_, CARRYB_13__8_, CARRYB_13__7_,
         CARRYB_13__6_, CARRYB_13__5_, CARRYB_13__4_, CARRYB_13__3_,
         CARRYB_13__2_, CARRYB_13__1_, CARRYB_13__0_, CARRYB_12__22_,
         CARRYB_12__21_, CARRYB_12__20_, CARRYB_12__19_, CARRYB_12__18_,
         CARRYB_12__17_, CARRYB_12__16_, CARRYB_12__15_, CARRYB_12__14_,
         CARRYB_12__13_, CARRYB_12__12_, CARRYB_12__11_, CARRYB_12__10_,
         CARRYB_12__9_, CARRYB_12__8_, CARRYB_12__7_, CARRYB_12__6_,
         CARRYB_12__5_, CARRYB_12__4_, CARRYB_12__3_, CARRYB_12__2_,
         CARRYB_12__1_, CARRYB_12__0_, CARRYB_11__22_, CARRYB_11__21_,
         CARRYB_11__20_, CARRYB_11__19_, CARRYB_11__18_, CARRYB_11__17_,
         CARRYB_11__16_, CARRYB_11__15_, CARRYB_11__14_, CARRYB_11__13_,
         CARRYB_11__12_, CARRYB_11__11_, CARRYB_11__10_, CARRYB_11__9_,
         CARRYB_11__8_, CARRYB_11__7_, CARRYB_11__6_, CARRYB_11__5_,
         CARRYB_11__4_, CARRYB_11__3_, CARRYB_11__2_, CARRYB_11__1_,
         CARRYB_11__0_, CARRYB_10__22_, CARRYB_10__21_, CARRYB_10__20_,
         CARRYB_10__19_, CARRYB_10__18_, CARRYB_10__17_, CARRYB_10__16_,
         CARRYB_10__15_, CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_,
         CARRYB_10__11_, CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_,
         CARRYB_10__7_, CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_,
         CARRYB_10__3_, CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_,
         CARRYB_9__22_, CARRYB_9__21_, CARRYB_9__20_, CARRYB_9__19_,
         CARRYB_9__18_, CARRYB_9__17_, CARRYB_9__16_, CARRYB_9__15_,
         CARRYB_9__14_, CARRYB_9__13_, CARRYB_9__12_, CARRYB_9__11_,
         CARRYB_9__10_, CARRYB_9__9_, CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_,
         CARRYB_9__5_, CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_,
         CARRYB_9__0_, CARRYB_8__22_, CARRYB_8__21_, CARRYB_8__20_,
         CARRYB_8__19_, CARRYB_8__18_, CARRYB_8__17_, CARRYB_8__16_,
         CARRYB_8__15_, CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_,
         CARRYB_8__11_, CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_,
         CARRYB_8__7_, CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_,
         CARRYB_8__2_, CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__22_,
         CARRYB_7__21_, CARRYB_7__20_, CARRYB_7__19_, CARRYB_7__18_,
         CARRYB_7__17_, CARRYB_7__16_, CARRYB_7__15_, CARRYB_7__14_,
         CARRYB_7__13_, CARRYB_7__12_, CARRYB_7__11_, CARRYB_7__10_,
         CARRYB_7__9_, CARRYB_7__8_, CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_,
         CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_,
         CARRYB_6__22_, CARRYB_6__21_, CARRYB_6__20_, CARRYB_6__19_,
         CARRYB_6__18_, CARRYB_6__17_, CARRYB_6__16_, CARRYB_6__15_,
         CARRYB_6__14_, CARRYB_6__13_, CARRYB_6__12_, CARRYB_6__11_,
         CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_, CARRYB_6__7_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__22_, CARRYB_5__21_, CARRYB_5__20_,
         CARRYB_5__19_, CARRYB_5__18_, CARRYB_5__17_, CARRYB_5__16_,
         CARRYB_5__15_, CARRYB_5__14_, CARRYB_5__13_, CARRYB_5__12_,
         CARRYB_5__11_, CARRYB_5__10_, CARRYB_5__9_, CARRYB_5__8_,
         CARRYB_5__7_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__22_,
         CARRYB_4__21_, CARRYB_4__20_, CARRYB_4__19_, CARRYB_4__18_,
         CARRYB_4__17_, CARRYB_4__16_, CARRYB_4__15_, CARRYB_4__14_,
         CARRYB_4__13_, CARRYB_4__12_, CARRYB_4__11_, CARRYB_4__10_,
         CARRYB_4__9_, CARRYB_4__8_, CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__22_, CARRYB_3__21_, CARRYB_3__20_, CARRYB_3__19_,
         CARRYB_3__18_, CARRYB_3__17_, CARRYB_3__16_, CARRYB_3__15_,
         CARRYB_3__14_, CARRYB_3__13_, CARRYB_3__12_, CARRYB_3__11_,
         CARRYB_3__10_, CARRYB_3__9_, CARRYB_3__8_, CARRYB_3__7_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__22_, CARRYB_2__21_, CARRYB_2__20_,
         CARRYB_2__19_, CARRYB_2__18_, CARRYB_2__17_, CARRYB_2__16_,
         CARRYB_2__15_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__22_,
         CARRYB_1__21_, CARRYB_1__20_, CARRYB_1__19_, CARRYB_1__18_,
         CARRYB_1__17_, CARRYB_1__16_, CARRYB_1__15_, CARRYB_1__14_,
         CARRYB_1__13_, CARRYB_1__12_, CARRYB_1__11_, CARRYB_1__10_,
         CARRYB_1__9_, CARRYB_1__8_, CARRYB_1__7_, CARRYB_1__6_, CARRYB_1__5_,
         CARRYB_1__4_, CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_,
         SUMB_23__23_, SUMB_23__22_, SUMB_23__21_, SUMB_23__20_, SUMB_23__19_,
         SUMB_23__18_, SUMB_23__17_, SUMB_23__16_, SUMB_23__15_, SUMB_23__14_,
         SUMB_23__13_, SUMB_23__12_, SUMB_23__11_, SUMB_23__10_, SUMB_23__9_,
         SUMB_23__8_, SUMB_23__7_, SUMB_23__6_, SUMB_23__5_, SUMB_23__4_,
         SUMB_23__3_, SUMB_23__2_, SUMB_23__1_, SUMB_23__0_, SUMB_22__22_,
         SUMB_22__21_, SUMB_22__20_, SUMB_22__19_, SUMB_22__18_, SUMB_22__17_,
         SUMB_22__16_, SUMB_22__15_, SUMB_22__14_, SUMB_22__13_, SUMB_22__12_,
         SUMB_22__11_, SUMB_22__10_, SUMB_22__9_, SUMB_22__8_, SUMB_22__7_,
         SUMB_22__6_, SUMB_22__5_, SUMB_22__4_, SUMB_22__3_, SUMB_22__2_,
         SUMB_22__1_, SUMB_21__22_, SUMB_21__21_, SUMB_21__20_, SUMB_21__19_,
         SUMB_21__18_, SUMB_21__17_, SUMB_21__16_, SUMB_21__15_, SUMB_21__14_,
         SUMB_21__13_, SUMB_21__12_, SUMB_21__11_, SUMB_21__10_, SUMB_21__9_,
         SUMB_21__8_, SUMB_21__7_, SUMB_21__6_, SUMB_21__5_, SUMB_21__4_,
         SUMB_21__3_, SUMB_21__2_, SUMB_21__1_, SUMB_20__22_, SUMB_20__21_,
         SUMB_20__20_, SUMB_20__19_, SUMB_20__18_, SUMB_20__17_, SUMB_20__16_,
         SUMB_20__15_, SUMB_20__14_, SUMB_20__13_, SUMB_20__12_, SUMB_20__11_,
         SUMB_20__10_, SUMB_20__9_, SUMB_20__8_, SUMB_20__7_, SUMB_20__6_,
         SUMB_20__5_, SUMB_20__4_, SUMB_20__3_, SUMB_20__2_, SUMB_20__1_,
         SUMB_19__22_, SUMB_19__21_, SUMB_19__20_, SUMB_19__19_, SUMB_19__18_,
         SUMB_19__17_, SUMB_19__16_, SUMB_19__15_, SUMB_19__14_, SUMB_19__13_,
         SUMB_19__12_, SUMB_19__11_, SUMB_19__10_, SUMB_19__9_, SUMB_19__8_,
         SUMB_19__7_, SUMB_19__6_, SUMB_19__5_, SUMB_19__4_, SUMB_19__3_,
         SUMB_19__2_, SUMB_19__1_, SUMB_18__22_, SUMB_18__21_, SUMB_18__20_,
         SUMB_18__19_, SUMB_18__18_, SUMB_18__17_, SUMB_18__16_, SUMB_18__15_,
         SUMB_18__14_, SUMB_18__13_, SUMB_18__12_, SUMB_18__11_, SUMB_18__10_,
         SUMB_18__9_, SUMB_18__8_, SUMB_18__7_, SUMB_18__6_, SUMB_18__5_,
         SUMB_18__4_, SUMB_18__3_, SUMB_18__2_, SUMB_18__1_, SUMB_17__22_,
         SUMB_17__21_, SUMB_17__20_, SUMB_17__19_, SUMB_17__18_, SUMB_17__17_,
         SUMB_17__16_, SUMB_17__15_, SUMB_17__14_, SUMB_17__13_, SUMB_17__12_,
         SUMB_17__11_, SUMB_17__10_, SUMB_17__9_, SUMB_17__8_, SUMB_17__7_,
         SUMB_17__6_, SUMB_17__5_, SUMB_17__4_, SUMB_17__3_, SUMB_17__2_,
         SUMB_17__1_, SUMB_16__22_, SUMB_16__21_, SUMB_16__20_, SUMB_16__19_,
         SUMB_16__18_, SUMB_16__17_, SUMB_16__16_, SUMB_16__15_, SUMB_16__14_,
         SUMB_16__13_, SUMB_16__12_, SUMB_16__11_, SUMB_16__10_, SUMB_16__9_,
         SUMB_16__8_, SUMB_16__7_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_,
         SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, SUMB_15__22_, SUMB_15__21_,
         SUMB_15__20_, SUMB_15__19_, SUMB_15__18_, SUMB_15__17_, SUMB_15__16_,
         SUMB_15__15_, SUMB_15__14_, SUMB_15__13_, SUMB_15__12_, SUMB_15__11_,
         SUMB_15__10_, SUMB_15__9_, SUMB_15__8_, SUMB_15__7_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_14__22_, SUMB_14__21_, SUMB_14__20_, SUMB_14__19_, SUMB_14__18_,
         SUMB_14__17_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_, SUMB_14__13_,
         SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_, SUMB_14__8_,
         SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_,
         SUMB_14__2_, SUMB_14__1_, SUMB_13__22_, SUMB_13__21_, SUMB_13__20_,
         SUMB_13__19_, SUMB_13__18_, SUMB_13__17_, SUMB_13__16_, SUMB_13__15_,
         SUMB_13__14_, SUMB_13__13_, SUMB_13__12_, SUMB_13__11_, SUMB_13__10_,
         SUMB_13__9_, SUMB_13__8_, SUMB_13__7_, SUMB_13__6_, SUMB_13__5_,
         SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_, SUMB_12__22_,
         SUMB_12__21_, SUMB_12__20_, SUMB_12__19_, SUMB_12__18_, SUMB_12__17_,
         SUMB_12__16_, SUMB_12__15_, SUMB_12__14_, SUMB_12__13_, SUMB_12__12_,
         SUMB_12__11_, SUMB_12__10_, SUMB_12__9_, SUMB_12__8_, SUMB_12__7_,
         SUMB_12__6_, SUMB_12__5_, SUMB_12__4_, SUMB_12__3_, SUMB_12__2_,
         SUMB_12__1_, SUMB_11__22_, SUMB_11__21_, SUMB_11__20_, SUMB_11__19_,
         SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_, SUMB_11__14_,
         SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_, SUMB_11__9_,
         SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_, SUMB_11__4_,
         SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__22_, SUMB_10__21_,
         SUMB_10__20_, SUMB_10__19_, SUMB_10__18_, SUMB_10__17_, SUMB_10__16_,
         SUMB_10__15_, SUMB_10__14_, SUMB_10__13_, SUMB_10__12_, SUMB_10__11_,
         SUMB_10__10_, SUMB_10__9_, SUMB_10__8_, SUMB_10__7_, SUMB_10__6_,
         SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_,
         SUMB_9__22_, SUMB_9__21_, SUMB_9__20_, SUMB_9__19_, SUMB_9__18_,
         SUMB_9__17_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_, SUMB_9__13_,
         SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_, SUMB_9__8_,
         SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_,
         SUMB_9__2_, SUMB_9__1_, SUMB_8__22_, SUMB_8__21_, SUMB_8__20_,
         SUMB_8__19_, SUMB_8__18_, SUMB_8__17_, SUMB_8__16_, SUMB_8__15_,
         SUMB_8__14_, SUMB_8__13_, SUMB_8__12_, SUMB_8__11_, SUMB_8__10_,
         SUMB_8__9_, SUMB_8__8_, SUMB_8__7_, SUMB_8__6_, SUMB_8__5_,
         SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_, SUMB_7__22_,
         SUMB_7__21_, SUMB_7__20_, SUMB_7__19_, SUMB_7__18_, SUMB_7__17_,
         SUMB_7__16_, SUMB_7__15_, SUMB_7__14_, SUMB_7__13_, SUMB_7__12_,
         SUMB_7__11_, SUMB_7__10_, SUMB_7__9_, SUMB_7__8_, SUMB_7__7_,
         SUMB_7__6_, SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_,
         SUMB_7__1_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_, SUMB_6__19_,
         SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_, SUMB_6__14_,
         SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_, SUMB_6__9_,
         SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_,
         SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__22_, SUMB_5__21_,
         SUMB_5__20_, SUMB_5__19_, SUMB_5__18_, SUMB_5__17_, SUMB_5__16_,
         SUMB_5__15_, SUMB_5__14_, SUMB_5__13_, SUMB_5__12_, SUMB_5__11_,
         SUMB_5__10_, SUMB_5__9_, SUMB_5__8_, SUMB_5__7_, SUMB_5__6_,
         SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_,
         SUMB_4__22_, SUMB_4__21_, SUMB_4__20_, SUMB_4__19_, SUMB_4__18_,
         SUMB_4__17_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_, SUMB_4__13_,
         SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_, SUMB_4__8_,
         SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_,
         SUMB_4__2_, SUMB_4__1_, SUMB_3__22_, SUMB_3__21_, SUMB_3__20_,
         SUMB_3__19_, SUMB_3__18_, SUMB_3__17_, SUMB_3__16_, SUMB_3__15_,
         SUMB_3__14_, SUMB_3__13_, SUMB_3__12_, SUMB_3__11_, SUMB_3__10_,
         SUMB_3__9_, SUMB_3__8_, SUMB_3__7_, SUMB_3__6_, SUMB_3__5_,
         SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_, SUMB_2__22_,
         SUMB_2__21_, SUMB_2__20_, SUMB_2__19_, SUMB_2__18_, SUMB_2__17_,
         SUMB_2__16_, SUMB_2__15_, SUMB_2__14_, SUMB_2__13_, SUMB_2__12_,
         SUMB_2__11_, SUMB_2__10_, SUMB_2__9_, SUMB_2__8_, SUMB_2__7_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__22_, SUMB_1__21_, SUMB_1__20_, SUMB_1__19_,
         SUMB_1__18_, SUMB_1__17_, SUMB_1__16_, SUMB_1__15_, SUMB_1__14_,
         SUMB_1__13_, SUMB_1__12_, SUMB_1__11_, SUMB_1__10_, SUMB_1__9_,
         SUMB_1__8_, SUMB_1__7_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_,
         SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, QA, QB, A1_45_, A1_44_, A1_43_,
         A1_42_, A1_41_, A1_40_, A1_39_, A1_38_, A1_37_, A1_36_, A1_35_,
         A1_34_, A1_33_, A1_32_, A1_31_, A1_30_, A1_29_, A1_28_, A1_27_,
         A1_26_, A1_25_, A1_24_, A1_23_, A1_22_, A1_21_, A1_20_, A1_19_,
         A1_18_, A1_17_, A1_16_, A1_15_, A1_14_, A1_13_, A1_12_, A1_11_,
         A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_,
         A1_0_, A2_45_, A2_44_, A2_43_, A2_42_, A2_41_, A2_40_, A2_39_, A2_38_,
         A2_37_, A2_36_, A2_35_, A2_34_, A2_33_, A2_32_, A2_31_, A2_30_,
         A2_29_, A2_28_, A2_27_, A2_26_, A2_25_, A2_24_, A2_23_, A2_22_, n1,
         n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21;

  FA_X1 S14_23_0 ( .A(A[23]), .B(B[23]), .CI(SUMB_23__0_), .CO(A2_22_), .S(
        A1_21_) );
  FA_X1 S4_0 ( .A(ab_23__0_), .B(CARRYB_22__0_), .CI(SUMB_22__1_), .CO(
        CARRYB_23__0_), .S(SUMB_23__0_) );
  FA_X1 S4_1 ( .A(ab_23__1_), .B(CARRYB_22__1_), .CI(SUMB_22__2_), .CO(
        CARRYB_23__1_), .S(SUMB_23__1_) );
  FA_X1 S4_2 ( .A(ab_23__2_), .B(CARRYB_22__2_), .CI(SUMB_22__3_), .CO(
        CARRYB_23__2_), .S(SUMB_23__2_) );
  FA_X1 S4_3 ( .A(ab_23__3_), .B(CARRYB_22__3_), .CI(SUMB_22__4_), .CO(
        CARRYB_23__3_), .S(SUMB_23__3_) );
  FA_X1 S4_4 ( .A(ab_23__4_), .B(CARRYB_22__4_), .CI(SUMB_22__5_), .CO(
        CARRYB_23__4_), .S(SUMB_23__4_) );
  FA_X1 S4_5 ( .A(ab_23__5_), .B(CARRYB_22__5_), .CI(SUMB_22__6_), .CO(
        CARRYB_23__5_), .S(SUMB_23__5_) );
  FA_X1 S4_6 ( .A(ab_23__6_), .B(CARRYB_22__6_), .CI(SUMB_22__7_), .CO(
        CARRYB_23__6_), .S(SUMB_23__6_) );
  FA_X1 S4_7 ( .A(ab_23__7_), .B(CARRYB_22__7_), .CI(SUMB_22__8_), .CO(
        CARRYB_23__7_), .S(SUMB_23__7_) );
  FA_X1 S4_8 ( .A(ab_23__8_), .B(CARRYB_22__8_), .CI(SUMB_22__9_), .CO(
        CARRYB_23__8_), .S(SUMB_23__8_) );
  FA_X1 S4_9 ( .A(ab_23__9_), .B(CARRYB_22__9_), .CI(SUMB_22__10_), .CO(
        CARRYB_23__9_), .S(SUMB_23__9_) );
  FA_X1 S4_10 ( .A(ab_23__10_), .B(CARRYB_22__10_), .CI(SUMB_22__11_), .CO(
        CARRYB_23__10_), .S(SUMB_23__10_) );
  FA_X1 S4_11 ( .A(ab_23__11_), .B(CARRYB_22__11_), .CI(SUMB_22__12_), .CO(
        CARRYB_23__11_), .S(SUMB_23__11_) );
  FA_X1 S4_12 ( .A(ab_23__12_), .B(CARRYB_22__12_), .CI(SUMB_22__13_), .CO(
        CARRYB_23__12_), .S(SUMB_23__12_) );
  FA_X1 S4_13 ( .A(ab_23__13_), .B(CARRYB_22__13_), .CI(SUMB_22__14_), .CO(
        CARRYB_23__13_), .S(SUMB_23__13_) );
  FA_X1 S4_14 ( .A(ab_23__14_), .B(CARRYB_22__14_), .CI(SUMB_22__15_), .CO(
        CARRYB_23__14_), .S(SUMB_23__14_) );
  FA_X1 S4_15 ( .A(ab_23__15_), .B(CARRYB_22__15_), .CI(SUMB_22__16_), .CO(
        CARRYB_23__15_), .S(SUMB_23__15_) );
  FA_X1 S4_16 ( .A(ab_23__16_), .B(CARRYB_22__16_), .CI(SUMB_22__17_), .CO(
        CARRYB_23__16_), .S(SUMB_23__16_) );
  FA_X1 S4_17 ( .A(ab_23__17_), .B(CARRYB_22__17_), .CI(SUMB_22__18_), .CO(
        CARRYB_23__17_), .S(SUMB_23__17_) );
  FA_X1 S4_18 ( .A(ab_23__18_), .B(CARRYB_22__18_), .CI(SUMB_22__19_), .CO(
        CARRYB_23__18_), .S(SUMB_23__18_) );
  FA_X1 S4_19 ( .A(ab_23__19_), .B(CARRYB_22__19_), .CI(SUMB_22__20_), .CO(
        CARRYB_23__19_), .S(SUMB_23__19_) );
  FA_X1 S4_20 ( .A(ab_23__20_), .B(CARRYB_22__20_), .CI(SUMB_22__21_), .CO(
        CARRYB_23__20_), .S(SUMB_23__20_) );
  FA_X1 S4_21 ( .A(ab_23__21_), .B(CARRYB_22__21_), .CI(SUMB_22__22_), .CO(
        CARRYB_23__21_), .S(SUMB_23__21_) );
  FA_X1 S5_22 ( .A(ab_23__22_), .B(CARRYB_22__22_), .CI(ab_22__23_), .CO(
        CARRYB_23__22_), .S(SUMB_23__22_) );
  FA_X1 S14_23 ( .A(n3), .B(n1), .CI(ab_23__23_), .CO(CARRYB_23__23_), .S(
        SUMB_23__23_) );
  FA_X1 S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), .CO(
        CARRYB_22__0_), .S(A1_20_) );
  FA_X1 S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), .CO(
        CARRYB_22__1_), .S(SUMB_22__1_) );
  FA_X1 S2_22_2 ( .A(ab_22__2_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), .CO(
        CARRYB_22__2_), .S(SUMB_22__2_) );
  FA_X1 S2_22_3 ( .A(ab_22__3_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), .CO(
        CARRYB_22__3_), .S(SUMB_22__3_) );
  FA_X1 S2_22_4 ( .A(ab_22__4_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), .CO(
        CARRYB_22__4_), .S(SUMB_22__4_) );
  FA_X1 S2_22_5 ( .A(ab_22__5_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), .CO(
        CARRYB_22__5_), .S(SUMB_22__5_) );
  FA_X1 S2_22_6 ( .A(ab_22__6_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), .CO(
        CARRYB_22__6_), .S(SUMB_22__6_) );
  FA_X1 S2_22_7 ( .A(ab_22__7_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), .CO(
        CARRYB_22__7_), .S(SUMB_22__7_) );
  FA_X1 S2_22_8 ( .A(ab_22__8_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), .CO(
        CARRYB_22__8_), .S(SUMB_22__8_) );
  FA_X1 S2_22_9 ( .A(ab_22__9_), .B(CARRYB_21__9_), .CI(SUMB_21__10_), .CO(
        CARRYB_22__9_), .S(SUMB_22__9_) );
  FA_X1 S2_22_10 ( .A(ab_22__10_), .B(CARRYB_21__10_), .CI(SUMB_21__11_), .CO(
        CARRYB_22__10_), .S(SUMB_22__10_) );
  FA_X1 S2_22_11 ( .A(ab_22__11_), .B(CARRYB_21__11_), .CI(SUMB_21__12_), .CO(
        CARRYB_22__11_), .S(SUMB_22__11_) );
  FA_X1 S2_22_12 ( .A(ab_22__12_), .B(CARRYB_21__12_), .CI(SUMB_21__13_), .CO(
        CARRYB_22__12_), .S(SUMB_22__12_) );
  FA_X1 S2_22_13 ( .A(ab_22__13_), .B(CARRYB_21__13_), .CI(SUMB_21__14_), .CO(
        CARRYB_22__13_), .S(SUMB_22__13_) );
  FA_X1 S2_22_14 ( .A(ab_22__14_), .B(CARRYB_21__14_), .CI(SUMB_21__15_), .CO(
        CARRYB_22__14_), .S(SUMB_22__14_) );
  FA_X1 S2_22_15 ( .A(ab_22__15_), .B(CARRYB_21__15_), .CI(SUMB_21__16_), .CO(
        CARRYB_22__15_), .S(SUMB_22__15_) );
  FA_X1 S2_22_16 ( .A(ab_22__16_), .B(CARRYB_21__16_), .CI(SUMB_21__17_), .CO(
        CARRYB_22__16_), .S(SUMB_22__16_) );
  FA_X1 S2_22_17 ( .A(ab_22__17_), .B(CARRYB_21__17_), .CI(SUMB_21__18_), .CO(
        CARRYB_22__17_), .S(SUMB_22__17_) );
  FA_X1 S2_22_18 ( .A(ab_22__18_), .B(CARRYB_21__18_), .CI(SUMB_21__19_), .CO(
        CARRYB_22__18_), .S(SUMB_22__18_) );
  FA_X1 S2_22_19 ( .A(ab_22__19_), .B(CARRYB_21__19_), .CI(SUMB_21__20_), .CO(
        CARRYB_22__19_), .S(SUMB_22__19_) );
  FA_X1 S2_22_20 ( .A(ab_22__20_), .B(CARRYB_21__20_), .CI(SUMB_21__21_), .CO(
        CARRYB_22__20_), .S(SUMB_22__20_) );
  FA_X1 S2_22_21 ( .A(ab_22__21_), .B(CARRYB_21__21_), .CI(SUMB_21__22_), .CO(
        CARRYB_22__21_), .S(SUMB_22__21_) );
  FA_X1 S3_22_22 ( .A(ab_22__22_), .B(CARRYB_21__22_), .CI(ab_21__23_), .CO(
        CARRYB_22__22_), .S(SUMB_22__22_) );
  FA_X1 S1_21_0 ( .A(ab_21__0_), .B(CARRYB_20__0_), .CI(SUMB_20__1_), .CO(
        CARRYB_21__0_), .S(A1_19_) );
  FA_X1 S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), .CO(
        CARRYB_21__1_), .S(SUMB_21__1_) );
  FA_X1 S2_21_2 ( .A(ab_21__2_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), .CO(
        CARRYB_21__2_), .S(SUMB_21__2_) );
  FA_X1 S2_21_3 ( .A(ab_21__3_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), .CO(
        CARRYB_21__3_), .S(SUMB_21__3_) );
  FA_X1 S2_21_4 ( .A(ab_21__4_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), .CO(
        CARRYB_21__4_), .S(SUMB_21__4_) );
  FA_X1 S2_21_5 ( .A(ab_21__5_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), .CO(
        CARRYB_21__5_), .S(SUMB_21__5_) );
  FA_X1 S2_21_6 ( .A(ab_21__6_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), .CO(
        CARRYB_21__6_), .S(SUMB_21__6_) );
  FA_X1 S2_21_7 ( .A(ab_21__7_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), .CO(
        CARRYB_21__7_), .S(SUMB_21__7_) );
  FA_X1 S2_21_8 ( .A(ab_21__8_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), .CO(
        CARRYB_21__8_), .S(SUMB_21__8_) );
  FA_X1 S2_21_9 ( .A(ab_21__9_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), .CO(
        CARRYB_21__9_), .S(SUMB_21__9_) );
  FA_X1 S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .CI(SUMB_20__11_), .CO(
        CARRYB_21__10_), .S(SUMB_21__10_) );
  FA_X1 S2_21_11 ( .A(ab_21__11_), .B(CARRYB_20__11_), .CI(SUMB_20__12_), .CO(
        CARRYB_21__11_), .S(SUMB_21__11_) );
  FA_X1 S2_21_12 ( .A(ab_21__12_), .B(CARRYB_20__12_), .CI(SUMB_20__13_), .CO(
        CARRYB_21__12_), .S(SUMB_21__12_) );
  FA_X1 S2_21_13 ( .A(ab_21__13_), .B(CARRYB_20__13_), .CI(SUMB_20__14_), .CO(
        CARRYB_21__13_), .S(SUMB_21__13_) );
  FA_X1 S2_21_14 ( .A(ab_21__14_), .B(CARRYB_20__14_), .CI(SUMB_20__15_), .CO(
        CARRYB_21__14_), .S(SUMB_21__14_) );
  FA_X1 S2_21_15 ( .A(ab_21__15_), .B(CARRYB_20__15_), .CI(SUMB_20__16_), .CO(
        CARRYB_21__15_), .S(SUMB_21__15_) );
  FA_X1 S2_21_16 ( .A(ab_21__16_), .B(CARRYB_20__16_), .CI(SUMB_20__17_), .CO(
        CARRYB_21__16_), .S(SUMB_21__16_) );
  FA_X1 S2_21_17 ( .A(ab_21__17_), .B(CARRYB_20__17_), .CI(SUMB_20__18_), .CO(
        CARRYB_21__17_), .S(SUMB_21__17_) );
  FA_X1 S2_21_18 ( .A(ab_21__18_), .B(CARRYB_20__18_), .CI(SUMB_20__19_), .CO(
        CARRYB_21__18_), .S(SUMB_21__18_) );
  FA_X1 S2_21_19 ( .A(ab_21__19_), .B(CARRYB_20__19_), .CI(SUMB_20__20_), .CO(
        CARRYB_21__19_), .S(SUMB_21__19_) );
  FA_X1 S2_21_20 ( .A(ab_21__20_), .B(CARRYB_20__20_), .CI(SUMB_20__21_), .CO(
        CARRYB_21__20_), .S(SUMB_21__20_) );
  FA_X1 S2_21_21 ( .A(ab_21__21_), .B(CARRYB_20__21_), .CI(SUMB_20__22_), .CO(
        CARRYB_21__21_), .S(SUMB_21__21_) );
  FA_X1 S3_21_22 ( .A(ab_21__22_), .B(CARRYB_20__22_), .CI(ab_20__23_), .CO(
        CARRYB_21__22_), .S(SUMB_21__22_) );
  FA_X1 S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), .CO(
        CARRYB_20__0_), .S(A1_18_) );
  FA_X1 S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), .CO(
        CARRYB_20__1_), .S(SUMB_20__1_) );
  FA_X1 S2_20_2 ( .A(ab_20__2_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), .CO(
        CARRYB_20__2_), .S(SUMB_20__2_) );
  FA_X1 S2_20_3 ( .A(ab_20__3_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), .CO(
        CARRYB_20__3_), .S(SUMB_20__3_) );
  FA_X1 S2_20_4 ( .A(ab_20__4_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), .CO(
        CARRYB_20__4_), .S(SUMB_20__4_) );
  FA_X1 S2_20_5 ( .A(ab_20__5_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), .CO(
        CARRYB_20__5_), .S(SUMB_20__5_) );
  FA_X1 S2_20_6 ( .A(ab_20__6_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), .CO(
        CARRYB_20__6_), .S(SUMB_20__6_) );
  FA_X1 S2_20_7 ( .A(ab_20__7_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), .CO(
        CARRYB_20__7_), .S(SUMB_20__7_) );
  FA_X1 S2_20_8 ( .A(ab_20__8_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), .CO(
        CARRYB_20__8_), .S(SUMB_20__8_) );
  FA_X1 S2_20_9 ( .A(ab_20__9_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), .CO(
        CARRYB_20__9_), .S(SUMB_20__9_) );
  FA_X1 S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), .CO(
        CARRYB_20__10_), .S(SUMB_20__10_) );
  FA_X1 S2_20_11 ( .A(ab_20__11_), .B(CARRYB_19__11_), .CI(SUMB_19__12_), .CO(
        CARRYB_20__11_), .S(SUMB_20__11_) );
  FA_X1 S2_20_12 ( .A(ab_20__12_), .B(CARRYB_19__12_), .CI(SUMB_19__13_), .CO(
        CARRYB_20__12_), .S(SUMB_20__12_) );
  FA_X1 S2_20_13 ( .A(ab_20__13_), .B(CARRYB_19__13_), .CI(SUMB_19__14_), .CO(
        CARRYB_20__13_), .S(SUMB_20__13_) );
  FA_X1 S2_20_14 ( .A(ab_20__14_), .B(CARRYB_19__14_), .CI(SUMB_19__15_), .CO(
        CARRYB_20__14_), .S(SUMB_20__14_) );
  FA_X1 S2_20_15 ( .A(ab_20__15_), .B(CARRYB_19__15_), .CI(SUMB_19__16_), .CO(
        CARRYB_20__15_), .S(SUMB_20__15_) );
  FA_X1 S2_20_16 ( .A(ab_20__16_), .B(CARRYB_19__16_), .CI(SUMB_19__17_), .CO(
        CARRYB_20__16_), .S(SUMB_20__16_) );
  FA_X1 S2_20_17 ( .A(ab_20__17_), .B(CARRYB_19__17_), .CI(SUMB_19__18_), .CO(
        CARRYB_20__17_), .S(SUMB_20__17_) );
  FA_X1 S2_20_18 ( .A(ab_20__18_), .B(CARRYB_19__18_), .CI(SUMB_19__19_), .CO(
        CARRYB_20__18_), .S(SUMB_20__18_) );
  FA_X1 S2_20_19 ( .A(ab_20__19_), .B(CARRYB_19__19_), .CI(SUMB_19__20_), .CO(
        CARRYB_20__19_), .S(SUMB_20__19_) );
  FA_X1 S2_20_20 ( .A(ab_20__20_), .B(CARRYB_19__20_), .CI(SUMB_19__21_), .CO(
        CARRYB_20__20_), .S(SUMB_20__20_) );
  FA_X1 S2_20_21 ( .A(ab_20__21_), .B(CARRYB_19__21_), .CI(SUMB_19__22_), .CO(
        CARRYB_20__21_), .S(SUMB_20__21_) );
  FA_X1 S3_20_22 ( .A(ab_20__22_), .B(CARRYB_19__22_), .CI(ab_19__23_), .CO(
        CARRYB_20__22_), .S(SUMB_20__22_) );
  FA_X1 S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), .CO(
        CARRYB_19__0_), .S(A1_17_) );
  FA_X1 S2_19_1 ( .A(ab_19__1_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), .CO(
        CARRYB_19__1_), .S(SUMB_19__1_) );
  FA_X1 S2_19_2 ( .A(ab_19__2_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), .CO(
        CARRYB_19__2_), .S(SUMB_19__2_) );
  FA_X1 S2_19_3 ( .A(ab_19__3_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), .CO(
        CARRYB_19__3_), .S(SUMB_19__3_) );
  FA_X1 S2_19_4 ( .A(ab_19__4_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), .CO(
        CARRYB_19__4_), .S(SUMB_19__4_) );
  FA_X1 S2_19_5 ( .A(ab_19__5_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), .CO(
        CARRYB_19__5_), .S(SUMB_19__5_) );
  FA_X1 S2_19_6 ( .A(ab_19__6_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), .CO(
        CARRYB_19__6_), .S(SUMB_19__6_) );
  FA_X1 S2_19_7 ( .A(ab_19__7_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), .CO(
        CARRYB_19__7_), .S(SUMB_19__7_) );
  FA_X1 S2_19_8 ( .A(ab_19__8_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), .CO(
        CARRYB_19__8_), .S(SUMB_19__8_) );
  FA_X1 S2_19_9 ( .A(ab_19__9_), .B(CARRYB_18__9_), .CI(SUMB_18__10_), .CO(
        CARRYB_19__9_), .S(SUMB_19__9_) );
  FA_X1 S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), .CO(
        CARRYB_19__10_), .S(SUMB_19__10_) );
  FA_X1 S2_19_11 ( .A(ab_19__11_), .B(CARRYB_18__11_), .CI(SUMB_18__12_), .CO(
        CARRYB_19__11_), .S(SUMB_19__11_) );
  FA_X1 S2_19_12 ( .A(ab_19__12_), .B(CARRYB_18__12_), .CI(SUMB_18__13_), .CO(
        CARRYB_19__12_), .S(SUMB_19__12_) );
  FA_X1 S2_19_13 ( .A(ab_19__13_), .B(CARRYB_18__13_), .CI(SUMB_18__14_), .CO(
        CARRYB_19__13_), .S(SUMB_19__13_) );
  FA_X1 S2_19_14 ( .A(ab_19__14_), .B(CARRYB_18__14_), .CI(SUMB_18__15_), .CO(
        CARRYB_19__14_), .S(SUMB_19__14_) );
  FA_X1 S2_19_15 ( .A(ab_19__15_), .B(CARRYB_18__15_), .CI(SUMB_18__16_), .CO(
        CARRYB_19__15_), .S(SUMB_19__15_) );
  FA_X1 S2_19_16 ( .A(ab_19__16_), .B(CARRYB_18__16_), .CI(SUMB_18__17_), .CO(
        CARRYB_19__16_), .S(SUMB_19__16_) );
  FA_X1 S2_19_17 ( .A(ab_19__17_), .B(CARRYB_18__17_), .CI(SUMB_18__18_), .CO(
        CARRYB_19__17_), .S(SUMB_19__17_) );
  FA_X1 S2_19_18 ( .A(ab_19__18_), .B(CARRYB_18__18_), .CI(SUMB_18__19_), .CO(
        CARRYB_19__18_), .S(SUMB_19__18_) );
  FA_X1 S2_19_19 ( .A(ab_19__19_), .B(CARRYB_18__19_), .CI(SUMB_18__20_), .CO(
        CARRYB_19__19_), .S(SUMB_19__19_) );
  FA_X1 S2_19_20 ( .A(ab_19__20_), .B(CARRYB_18__20_), .CI(SUMB_18__21_), .CO(
        CARRYB_19__20_), .S(SUMB_19__20_) );
  FA_X1 S2_19_21 ( .A(ab_19__21_), .B(CARRYB_18__21_), .CI(SUMB_18__22_), .CO(
        CARRYB_19__21_), .S(SUMB_19__21_) );
  FA_X1 S3_19_22 ( .A(ab_19__22_), .B(CARRYB_18__22_), .CI(ab_18__23_), .CO(
        CARRYB_19__22_), .S(SUMB_19__22_) );
  FA_X1 S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), .CO(
        CARRYB_18__0_), .S(A1_16_) );
  FA_X1 S2_18_1 ( .A(ab_18__1_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), .CO(
        CARRYB_18__1_), .S(SUMB_18__1_) );
  FA_X1 S2_18_2 ( .A(ab_18__2_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), .CO(
        CARRYB_18__2_), .S(SUMB_18__2_) );
  FA_X1 S2_18_3 ( .A(ab_18__3_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), .CO(
        CARRYB_18__3_), .S(SUMB_18__3_) );
  FA_X1 S2_18_4 ( .A(ab_18__4_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), .CO(
        CARRYB_18__4_), .S(SUMB_18__4_) );
  FA_X1 S2_18_5 ( .A(ab_18__5_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), .CO(
        CARRYB_18__5_), .S(SUMB_18__5_) );
  FA_X1 S2_18_6 ( .A(ab_18__6_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), .CO(
        CARRYB_18__6_), .S(SUMB_18__6_) );
  FA_X1 S2_18_7 ( .A(ab_18__7_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), .CO(
        CARRYB_18__7_), .S(SUMB_18__7_) );
  FA_X1 S2_18_8 ( .A(ab_18__8_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), .CO(
        CARRYB_18__8_), .S(SUMB_18__8_) );
  FA_X1 S2_18_9 ( .A(ab_18__9_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), .CO(
        CARRYB_18__9_), .S(SUMB_18__9_) );
  FA_X1 S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), .CO(
        CARRYB_18__10_), .S(SUMB_18__10_) );
  FA_X1 S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), .CO(
        CARRYB_18__11_), .S(SUMB_18__11_) );
  FA_X1 S2_18_12 ( .A(ab_18__12_), .B(CARRYB_17__12_), .CI(SUMB_17__13_), .CO(
        CARRYB_18__12_), .S(SUMB_18__12_) );
  FA_X1 S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .CI(SUMB_17__14_), .CO(
        CARRYB_18__13_), .S(SUMB_18__13_) );
  FA_X1 S2_18_14 ( .A(ab_18__14_), .B(CARRYB_17__14_), .CI(SUMB_17__15_), .CO(
        CARRYB_18__14_), .S(SUMB_18__14_) );
  FA_X1 S2_18_15 ( .A(ab_18__15_), .B(CARRYB_17__15_), .CI(SUMB_17__16_), .CO(
        CARRYB_18__15_), .S(SUMB_18__15_) );
  FA_X1 S2_18_16 ( .A(ab_18__16_), .B(CARRYB_17__16_), .CI(SUMB_17__17_), .CO(
        CARRYB_18__16_), .S(SUMB_18__16_) );
  FA_X1 S2_18_17 ( .A(ab_18__17_), .B(CARRYB_17__17_), .CI(SUMB_17__18_), .CO(
        CARRYB_18__17_), .S(SUMB_18__17_) );
  FA_X1 S2_18_18 ( .A(ab_18__18_), .B(CARRYB_17__18_), .CI(SUMB_17__19_), .CO(
        CARRYB_18__18_), .S(SUMB_18__18_) );
  FA_X1 S2_18_19 ( .A(ab_18__19_), .B(CARRYB_17__19_), .CI(SUMB_17__20_), .CO(
        CARRYB_18__19_), .S(SUMB_18__19_) );
  FA_X1 S2_18_20 ( .A(ab_18__20_), .B(CARRYB_17__20_), .CI(SUMB_17__21_), .CO(
        CARRYB_18__20_), .S(SUMB_18__20_) );
  FA_X1 S2_18_21 ( .A(ab_18__21_), .B(CARRYB_17__21_), .CI(SUMB_17__22_), .CO(
        CARRYB_18__21_), .S(SUMB_18__21_) );
  FA_X1 S3_18_22 ( .A(ab_18__22_), .B(CARRYB_17__22_), .CI(ab_17__23_), .CO(
        CARRYB_18__22_), .S(SUMB_18__22_) );
  FA_X1 S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), .CO(
        CARRYB_17__0_), .S(A1_15_) );
  FA_X1 S2_17_1 ( .A(ab_17__1_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), .CO(
        CARRYB_17__1_), .S(SUMB_17__1_) );
  FA_X1 S2_17_2 ( .A(ab_17__2_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), .CO(
        CARRYB_17__2_), .S(SUMB_17__2_) );
  FA_X1 S2_17_3 ( .A(ab_17__3_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), .CO(
        CARRYB_17__3_), .S(SUMB_17__3_) );
  FA_X1 S2_17_4 ( .A(ab_17__4_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), .CO(
        CARRYB_17__4_), .S(SUMB_17__4_) );
  FA_X1 S2_17_5 ( .A(ab_17__5_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), .CO(
        CARRYB_17__5_), .S(SUMB_17__5_) );
  FA_X1 S2_17_6 ( .A(ab_17__6_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), .CO(
        CARRYB_17__6_), .S(SUMB_17__6_) );
  FA_X1 S2_17_7 ( .A(ab_17__7_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), .CO(
        CARRYB_17__7_), .S(SUMB_17__7_) );
  FA_X1 S2_17_8 ( .A(ab_17__8_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), .CO(
        CARRYB_17__8_), .S(SUMB_17__8_) );
  FA_X1 S2_17_9 ( .A(ab_17__9_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), .CO(
        CARRYB_17__9_), .S(SUMB_17__9_) );
  FA_X1 S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), .CO(
        CARRYB_17__10_), .S(SUMB_17__10_) );
  FA_X1 S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), .CO(
        CARRYB_17__11_), .S(SUMB_17__11_) );
  FA_X1 S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), .CO(
        CARRYB_17__12_), .S(SUMB_17__12_) );
  FA_X1 S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), .CO(
        CARRYB_17__13_), .S(SUMB_17__13_) );
  FA_X1 S2_17_14 ( .A(ab_17__14_), .B(CARRYB_16__14_), .CI(SUMB_16__15_), .CO(
        CARRYB_17__14_), .S(SUMB_17__14_) );
  FA_X1 S2_17_15 ( .A(ab_17__15_), .B(CARRYB_16__15_), .CI(SUMB_16__16_), .CO(
        CARRYB_17__15_), .S(SUMB_17__15_) );
  FA_X1 S2_17_16 ( .A(ab_17__16_), .B(CARRYB_16__16_), .CI(SUMB_16__17_), .CO(
        CARRYB_17__16_), .S(SUMB_17__16_) );
  FA_X1 S2_17_17 ( .A(ab_17__17_), .B(CARRYB_16__17_), .CI(SUMB_16__18_), .CO(
        CARRYB_17__17_), .S(SUMB_17__17_) );
  FA_X1 S2_17_18 ( .A(ab_17__18_), .B(CARRYB_16__18_), .CI(SUMB_16__19_), .CO(
        CARRYB_17__18_), .S(SUMB_17__18_) );
  FA_X1 S2_17_19 ( .A(ab_17__19_), .B(CARRYB_16__19_), .CI(SUMB_16__20_), .CO(
        CARRYB_17__19_), .S(SUMB_17__19_) );
  FA_X1 S2_17_20 ( .A(ab_17__20_), .B(CARRYB_16__20_), .CI(SUMB_16__21_), .CO(
        CARRYB_17__20_), .S(SUMB_17__20_) );
  FA_X1 S2_17_21 ( .A(ab_17__21_), .B(CARRYB_16__21_), .CI(SUMB_16__22_), .CO(
        CARRYB_17__21_), .S(SUMB_17__21_) );
  FA_X1 S3_17_22 ( .A(ab_17__22_), .B(CARRYB_16__22_), .CI(ab_16__23_), .CO(
        CARRYB_17__22_), .S(SUMB_17__22_) );
  FA_X1 S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(A1_14_) );
  FA_X1 S2_16_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  FA_X1 S2_16_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  FA_X1 S2_16_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  FA_X1 S2_16_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  FA_X1 S2_16_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  FA_X1 S2_16_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  FA_X1 S2_16_7 ( .A(ab_16__7_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), .CO(
        CARRYB_16__7_), .S(SUMB_16__7_) );
  FA_X1 S2_16_8 ( .A(ab_16__8_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), .CO(
        CARRYB_16__8_), .S(SUMB_16__8_) );
  FA_X1 S2_16_9 ( .A(ab_16__9_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), .CO(
        CARRYB_16__9_), .S(SUMB_16__9_) );
  FA_X1 S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), .CO(
        CARRYB_16__10_), .S(SUMB_16__10_) );
  FA_X1 S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), .CO(
        CARRYB_16__11_), .S(SUMB_16__11_) );
  FA_X1 S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), .CO(
        CARRYB_16__12_), .S(SUMB_16__12_) );
  FA_X1 S2_16_13 ( .A(ab_16__13_), .B(CARRYB_15__13_), .CI(SUMB_15__14_), .CO(
        CARRYB_16__13_), .S(SUMB_16__13_) );
  FA_X1 S2_16_14 ( .A(ab_16__14_), .B(CARRYB_15__14_), .CI(SUMB_15__15_), .CO(
        CARRYB_16__14_), .S(SUMB_16__14_) );
  FA_X1 S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .CI(SUMB_15__16_), .CO(
        CARRYB_16__15_), .S(SUMB_16__15_) );
  FA_X1 S2_16_16 ( .A(ab_16__16_), .B(CARRYB_15__16_), .CI(SUMB_15__17_), .CO(
        CARRYB_16__16_), .S(SUMB_16__16_) );
  FA_X1 S2_16_17 ( .A(ab_16__17_), .B(CARRYB_15__17_), .CI(SUMB_15__18_), .CO(
        CARRYB_16__17_), .S(SUMB_16__17_) );
  FA_X1 S2_16_18 ( .A(ab_16__18_), .B(CARRYB_15__18_), .CI(SUMB_15__19_), .CO(
        CARRYB_16__18_), .S(SUMB_16__18_) );
  FA_X1 S2_16_19 ( .A(ab_16__19_), .B(CARRYB_15__19_), .CI(SUMB_15__20_), .CO(
        CARRYB_16__19_), .S(SUMB_16__19_) );
  FA_X1 S2_16_20 ( .A(ab_16__20_), .B(CARRYB_15__20_), .CI(SUMB_15__21_), .CO(
        CARRYB_16__20_), .S(SUMB_16__20_) );
  FA_X1 S2_16_21 ( .A(ab_16__21_), .B(CARRYB_15__21_), .CI(SUMB_15__22_), .CO(
        CARRYB_16__21_), .S(SUMB_16__21_) );
  FA_X1 S3_16_22 ( .A(ab_16__22_), .B(CARRYB_15__22_), .CI(ab_15__23_), .CO(
        CARRYB_16__22_), .S(SUMB_16__22_) );
  FA_X1 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  FA_X1 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  FA_X1 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  FA_X1 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  FA_X1 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  FA_X1 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  FA_X1 S2_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  FA_X1 S2_15_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), .CO(
        CARRYB_15__7_), .S(SUMB_15__7_) );
  FA_X1 S2_15_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), .CO(
        CARRYB_15__8_), .S(SUMB_15__8_) );
  FA_X1 S2_15_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), .CO(
        CARRYB_15__9_), .S(SUMB_15__9_) );
  FA_X1 S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), .CO(
        CARRYB_15__10_), .S(SUMB_15__10_) );
  FA_X1 S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), .CO(
        CARRYB_15__11_), .S(SUMB_15__11_) );
  FA_X1 S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), .CO(
        CARRYB_15__12_), .S(SUMB_15__12_) );
  FA_X1 S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), .CO(
        CARRYB_15__13_), .S(SUMB_15__13_) );
  FA_X1 S2_15_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), .CO(
        CARRYB_15__14_), .S(SUMB_15__14_) );
  FA_X1 S2_15_15 ( .A(ab_15__15_), .B(CARRYB_14__15_), .CI(SUMB_14__16_), .CO(
        CARRYB_15__15_), .S(SUMB_15__15_) );
  FA_X1 S2_15_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .CI(SUMB_14__17_), .CO(
        CARRYB_15__16_), .S(SUMB_15__16_) );
  FA_X1 S2_15_17 ( .A(ab_15__17_), .B(CARRYB_14__17_), .CI(SUMB_14__18_), .CO(
        CARRYB_15__17_), .S(SUMB_15__17_) );
  FA_X1 S2_15_18 ( .A(ab_15__18_), .B(CARRYB_14__18_), .CI(SUMB_14__19_), .CO(
        CARRYB_15__18_), .S(SUMB_15__18_) );
  FA_X1 S2_15_19 ( .A(ab_15__19_), .B(CARRYB_14__19_), .CI(SUMB_14__20_), .CO(
        CARRYB_15__19_), .S(SUMB_15__19_) );
  FA_X1 S2_15_20 ( .A(ab_15__20_), .B(CARRYB_14__20_), .CI(SUMB_14__21_), .CO(
        CARRYB_15__20_), .S(SUMB_15__20_) );
  FA_X1 S2_15_21 ( .A(ab_15__21_), .B(CARRYB_14__21_), .CI(SUMB_14__22_), .CO(
        CARRYB_15__21_), .S(SUMB_15__21_) );
  FA_X1 S3_15_22 ( .A(ab_15__22_), .B(CARRYB_14__22_), .CI(ab_14__23_), .CO(
        CARRYB_15__22_), .S(SUMB_15__22_) );
  FA_X1 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  FA_X1 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  FA_X1 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  FA_X1 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  FA_X1 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  FA_X1 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  FA_X1 S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  FA_X1 S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), .CO(
        CARRYB_14__7_), .S(SUMB_14__7_) );
  FA_X1 S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), .CO(
        CARRYB_14__8_), .S(SUMB_14__8_) );
  FA_X1 S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), .CO(
        CARRYB_14__9_), .S(SUMB_14__9_) );
  FA_X1 S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), .CO(
        CARRYB_14__10_), .S(SUMB_14__10_) );
  FA_X1 S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), .CO(
        CARRYB_14__11_), .S(SUMB_14__11_) );
  FA_X1 S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), .CO(
        CARRYB_14__12_), .S(SUMB_14__12_) );
  FA_X1 S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), .CO(
        CARRYB_14__13_), .S(SUMB_14__13_) );
  FA_X1 S2_14_14 ( .A(ab_14__14_), .B(CARRYB_13__14_), .CI(SUMB_13__15_), .CO(
        CARRYB_14__14_), .S(SUMB_14__14_) );
  FA_X1 S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), .CO(
        CARRYB_14__15_), .S(SUMB_14__15_) );
  FA_X1 S2_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), .CO(
        CARRYB_14__16_), .S(SUMB_14__16_) );
  FA_X1 S2_14_17 ( .A(ab_14__17_), .B(CARRYB_13__17_), .CI(SUMB_13__18_), .CO(
        CARRYB_14__17_), .S(SUMB_14__17_) );
  FA_X1 S2_14_18 ( .A(ab_14__18_), .B(CARRYB_13__18_), .CI(SUMB_13__19_), .CO(
        CARRYB_14__18_), .S(SUMB_14__18_) );
  FA_X1 S2_14_19 ( .A(ab_14__19_), .B(CARRYB_13__19_), .CI(SUMB_13__20_), .CO(
        CARRYB_14__19_), .S(SUMB_14__19_) );
  FA_X1 S2_14_20 ( .A(ab_14__20_), .B(CARRYB_13__20_), .CI(SUMB_13__21_), .CO(
        CARRYB_14__20_), .S(SUMB_14__20_) );
  FA_X1 S2_14_21 ( .A(ab_14__21_), .B(CARRYB_13__21_), .CI(SUMB_13__22_), .CO(
        CARRYB_14__21_), .S(SUMB_14__21_) );
  FA_X1 S3_14_22 ( .A(ab_14__22_), .B(CARRYB_13__22_), .CI(ab_13__23_), .CO(
        CARRYB_14__22_), .S(SUMB_14__22_) );
  FA_X1 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  FA_X1 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  FA_X1 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  FA_X1 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  FA_X1 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  FA_X1 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  FA_X1 S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  FA_X1 S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), .CO(
        CARRYB_13__7_), .S(SUMB_13__7_) );
  FA_X1 S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), .CO(
        CARRYB_13__8_), .S(SUMB_13__8_) );
  FA_X1 S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), .CO(
        CARRYB_13__9_), .S(SUMB_13__9_) );
  FA_X1 S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), .CO(
        CARRYB_13__10_), .S(SUMB_13__10_) );
  FA_X1 S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), .CO(
        CARRYB_13__11_), .S(SUMB_13__11_) );
  FA_X1 S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), .CO(
        CARRYB_13__12_), .S(SUMB_13__12_) );
  FA_X1 S2_13_13 ( .A(ab_13__13_), .B(CARRYB_12__13_), .CI(SUMB_12__14_), .CO(
        CARRYB_13__13_), .S(SUMB_13__13_) );
  FA_X1 S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), .CO(
        CARRYB_13__14_), .S(SUMB_13__14_) );
  FA_X1 S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), .CO(
        CARRYB_13__15_), .S(SUMB_13__15_) );
  FA_X1 S2_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), .CO(
        CARRYB_13__16_), .S(SUMB_13__16_) );
  FA_X1 S2_13_17 ( .A(ab_13__17_), .B(CARRYB_12__17_), .CI(SUMB_12__18_), .CO(
        CARRYB_13__17_), .S(SUMB_13__17_) );
  FA_X1 S2_13_18 ( .A(ab_13__18_), .B(CARRYB_12__18_), .CI(SUMB_12__19_), .CO(
        CARRYB_13__18_), .S(SUMB_13__18_) );
  FA_X1 S2_13_19 ( .A(ab_13__19_), .B(CARRYB_12__19_), .CI(SUMB_12__20_), .CO(
        CARRYB_13__19_), .S(SUMB_13__19_) );
  FA_X1 S2_13_20 ( .A(ab_13__20_), .B(CARRYB_12__20_), .CI(SUMB_12__21_), .CO(
        CARRYB_13__20_), .S(SUMB_13__20_) );
  FA_X1 S2_13_21 ( .A(ab_13__21_), .B(CARRYB_12__21_), .CI(SUMB_12__22_), .CO(
        CARRYB_13__21_), .S(SUMB_13__21_) );
  FA_X1 S3_13_22 ( .A(ab_13__22_), .B(CARRYB_12__22_), .CI(ab_12__23_), .CO(
        CARRYB_13__22_), .S(SUMB_13__22_) );
  FA_X1 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  FA_X1 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  FA_X1 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  FA_X1 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  FA_X1 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  FA_X1 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  FA_X1 S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  FA_X1 S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), .CO(
        CARRYB_12__7_), .S(SUMB_12__7_) );
  FA_X1 S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), .CO(
        CARRYB_12__8_), .S(SUMB_12__8_) );
  FA_X1 S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), .CO(
        CARRYB_12__9_), .S(SUMB_12__9_) );
  FA_X1 S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), .CO(
        CARRYB_12__10_), .S(SUMB_12__10_) );
  FA_X1 S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), .CO(
        CARRYB_12__11_), .S(SUMB_12__11_) );
  FA_X1 S2_12_12 ( .A(ab_12__12_), .B(CARRYB_11__12_), .CI(SUMB_11__13_), .CO(
        CARRYB_12__12_), .S(SUMB_12__12_) );
  FA_X1 S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), .CO(
        CARRYB_12__13_), .S(SUMB_12__13_) );
  FA_X1 S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), .CO(
        CARRYB_12__14_), .S(SUMB_12__14_) );
  FA_X1 S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), .CO(
        CARRYB_12__15_), .S(SUMB_12__15_) );
  FA_X1 S2_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), .CO(
        CARRYB_12__16_), .S(SUMB_12__16_) );
  FA_X1 S2_12_17 ( .A(ab_12__17_), .B(CARRYB_11__17_), .CI(SUMB_11__18_), .CO(
        CARRYB_12__17_), .S(SUMB_12__17_) );
  FA_X1 S2_12_18 ( .A(ab_12__18_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), .CO(
        CARRYB_12__18_), .S(SUMB_12__18_) );
  FA_X1 S2_12_19 ( .A(ab_12__19_), .B(CARRYB_11__19_), .CI(SUMB_11__20_), .CO(
        CARRYB_12__19_), .S(SUMB_12__19_) );
  FA_X1 S2_12_20 ( .A(ab_12__20_), .B(CARRYB_11__20_), .CI(SUMB_11__21_), .CO(
        CARRYB_12__20_), .S(SUMB_12__20_) );
  FA_X1 S2_12_21 ( .A(ab_12__21_), .B(CARRYB_11__21_), .CI(SUMB_11__22_), .CO(
        CARRYB_12__21_), .S(SUMB_12__21_) );
  FA_X1 S3_12_22 ( .A(ab_12__22_), .B(CARRYB_11__22_), .CI(ab_11__23_), .CO(
        CARRYB_12__22_), .S(SUMB_12__22_) );
  FA_X1 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  FA_X1 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  FA_X1 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  FA_X1 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  FA_X1 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  FA_X1 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  FA_X1 S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  FA_X1 S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), .CO(
        CARRYB_11__7_), .S(SUMB_11__7_) );
  FA_X1 S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), .CO(
        CARRYB_11__8_), .S(SUMB_11__8_) );
  FA_X1 S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), .CO(
        CARRYB_11__9_), .S(SUMB_11__9_) );
  FA_X1 S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), .CO(
        CARRYB_11__10_), .S(SUMB_11__10_) );
  FA_X1 S2_11_11 ( .A(ab_11__11_), .B(CARRYB_10__11_), .CI(SUMB_10__12_), .CO(
        CARRYB_11__11_), .S(SUMB_11__11_) );
  FA_X1 S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), .CO(
        CARRYB_11__12_), .S(SUMB_11__12_) );
  FA_X1 S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), .CO(
        CARRYB_11__13_), .S(SUMB_11__13_) );
  FA_X1 S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), .CO(
        CARRYB_11__14_), .S(SUMB_11__14_) );
  FA_X1 S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), .CO(
        CARRYB_11__15_), .S(SUMB_11__15_) );
  FA_X1 S2_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(SUMB_10__17_), .CO(
        CARRYB_11__16_), .S(SUMB_11__16_) );
  FA_X1 S2_11_17 ( .A(ab_11__17_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), .CO(
        CARRYB_11__17_), .S(SUMB_11__17_) );
  FA_X1 S2_11_18 ( .A(ab_11__18_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), .CO(
        CARRYB_11__18_), .S(SUMB_11__18_) );
  FA_X1 S2_11_19 ( .A(ab_11__19_), .B(CARRYB_10__19_), .CI(SUMB_10__20_), .CO(
        CARRYB_11__19_), .S(SUMB_11__19_) );
  FA_X1 S2_11_20 ( .A(ab_11__20_), .B(CARRYB_10__20_), .CI(SUMB_10__21_), .CO(
        CARRYB_11__20_), .S(SUMB_11__20_) );
  FA_X1 S2_11_21 ( .A(ab_11__21_), .B(CARRYB_10__21_), .CI(SUMB_10__22_), .CO(
        CARRYB_11__21_), .S(SUMB_11__21_) );
  FA_X1 S3_11_22 ( .A(ab_11__22_), .B(CARRYB_10__22_), .CI(ab_10__23_), .CO(
        CARRYB_11__22_), .S(SUMB_11__22_) );
  FA_X1 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  FA_X1 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  FA_X1 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  FA_X1 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  FA_X1 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  FA_X1 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  FA_X1 S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  FA_X1 S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  FA_X1 S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  FA_X1 S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  FA_X1 S2_10_10 ( .A(ab_10__10_), .B(CARRYB_9__10_), .CI(SUMB_9__11_), .CO(
        CARRYB_10__10_), .S(SUMB_10__10_) );
  FA_X1 S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), .CO(
        CARRYB_10__11_), .S(SUMB_10__11_) );
  FA_X1 S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), .CO(
        CARRYB_10__12_), .S(SUMB_10__12_) );
  FA_X1 S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), .CO(
        CARRYB_10__13_), .S(SUMB_10__13_) );
  FA_X1 S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), .CO(
        CARRYB_10__14_), .S(SUMB_10__14_) );
  FA_X1 S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), .CO(
        CARRYB_10__15_), .S(SUMB_10__15_) );
  FA_X1 S2_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), .CO(
        CARRYB_10__16_), .S(SUMB_10__16_) );
  FA_X1 S2_10_17 ( .A(ab_10__17_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), .CO(
        CARRYB_10__17_), .S(SUMB_10__17_) );
  FA_X1 S2_10_18 ( .A(ab_10__18_), .B(CARRYB_9__18_), .CI(SUMB_9__19_), .CO(
        CARRYB_10__18_), .S(SUMB_10__18_) );
  FA_X1 S2_10_19 ( .A(ab_10__19_), .B(CARRYB_9__19_), .CI(SUMB_9__20_), .CO(
        CARRYB_10__19_), .S(SUMB_10__19_) );
  FA_X1 S2_10_20 ( .A(ab_10__20_), .B(CARRYB_9__20_), .CI(SUMB_9__21_), .CO(
        CARRYB_10__20_), .S(SUMB_10__20_) );
  FA_X1 S2_10_21 ( .A(ab_10__21_), .B(CARRYB_9__21_), .CI(SUMB_9__22_), .CO(
        CARRYB_10__21_), .S(SUMB_10__21_) );
  FA_X1 S3_10_22 ( .A(ab_10__22_), .B(CARRYB_9__22_), .CI(ab_9__23_), .CO(
        CARRYB_10__22_), .S(SUMB_10__22_) );
  FA_X1 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  FA_X1 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  FA_X1 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  FA_X1 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  FA_X1 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  FA_X1 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  FA_X1 S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  FA_X1 S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  FA_X1 S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  FA_X1 S2_9_9 ( .A(ab_9__9_), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  FA_X1 S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), .CO(
        CARRYB_9__10_), .S(SUMB_9__10_) );
  FA_X1 S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), .CO(
        CARRYB_9__11_), .S(SUMB_9__11_) );
  FA_X1 S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), .CO(
        CARRYB_9__12_), .S(SUMB_9__12_) );
  FA_X1 S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), .CO(
        CARRYB_9__13_), .S(SUMB_9__13_) );
  FA_X1 S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), .CO(
        CARRYB_9__14_), .S(SUMB_9__14_) );
  FA_X1 S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), .CO(
        CARRYB_9__15_), .S(SUMB_9__15_) );
  FA_X1 S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), .CO(
        CARRYB_9__16_), .S(SUMB_9__16_) );
  FA_X1 S2_9_17 ( .A(ab_9__17_), .B(CARRYB_8__17_), .CI(SUMB_8__18_), .CO(
        CARRYB_9__17_), .S(SUMB_9__17_) );
  FA_X1 S2_9_18 ( .A(ab_9__18_), .B(CARRYB_8__18_), .CI(SUMB_8__19_), .CO(
        CARRYB_9__18_), .S(SUMB_9__18_) );
  FA_X1 S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), .CO(
        CARRYB_9__19_), .S(SUMB_9__19_) );
  FA_X1 S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(SUMB_8__21_), .CO(
        CARRYB_9__20_), .S(SUMB_9__20_) );
  FA_X1 S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), .CO(
        CARRYB_9__21_), .S(SUMB_9__21_) );
  FA_X1 S3_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .CI(ab_8__23_), .CO(
        CARRYB_9__22_), .S(SUMB_9__22_) );
  FA_X1 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  FA_X1 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  FA_X1 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  FA_X1 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  FA_X1 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  FA_X1 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  FA_X1 S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  FA_X1 S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  FA_X1 S2_8_8 ( .A(ab_8__8_), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  FA_X1 S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  FA_X1 S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), .CO(
        CARRYB_8__10_), .S(SUMB_8__10_) );
  FA_X1 S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), .CO(
        CARRYB_8__11_), .S(SUMB_8__11_) );
  FA_X1 S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), .CO(
        CARRYB_8__12_), .S(SUMB_8__12_) );
  FA_X1 S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), .CO(
        CARRYB_8__13_), .S(SUMB_8__13_) );
  FA_X1 S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), .CO(
        CARRYB_8__14_), .S(SUMB_8__14_) );
  FA_X1 S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), .CO(
        CARRYB_8__15_), .S(SUMB_8__15_) );
  FA_X1 S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), .CO(
        CARRYB_8__16_), .S(SUMB_8__16_) );
  FA_X1 S2_8_17 ( .A(ab_8__17_), .B(CARRYB_7__17_), .CI(SUMB_7__18_), .CO(
        CARRYB_8__17_), .S(SUMB_8__17_) );
  FA_X1 S2_8_18 ( .A(ab_8__18_), .B(CARRYB_7__18_), .CI(SUMB_7__19_), .CO(
        CARRYB_8__18_), .S(SUMB_8__18_) );
  FA_X1 S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), .CO(
        CARRYB_8__19_), .S(SUMB_8__19_) );
  FA_X1 S2_8_20 ( .A(ab_8__20_), .B(CARRYB_7__20_), .CI(SUMB_7__21_), .CO(
        CARRYB_8__20_), .S(SUMB_8__20_) );
  FA_X1 S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), .CO(
        CARRYB_8__21_), .S(SUMB_8__21_) );
  FA_X1 S3_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(ab_7__23_), .CO(
        CARRYB_8__22_), .S(SUMB_8__22_) );
  FA_X1 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(A1_5_) );
  FA_X1 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S2_7_7 ( .A(ab_7__7_), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  FA_X1 S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  FA_X1 S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  FA_X1 S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), .CO(
        CARRYB_7__10_), .S(SUMB_7__10_) );
  FA_X1 S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), .CO(
        CARRYB_7__11_), .S(SUMB_7__11_) );
  FA_X1 S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), .CO(
        CARRYB_7__12_), .S(SUMB_7__12_) );
  FA_X1 S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), .CO(
        CARRYB_7__13_), .S(SUMB_7__13_) );
  FA_X1 S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), .CO(
        CARRYB_7__14_), .S(SUMB_7__14_) );
  FA_X1 S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), .CO(
        CARRYB_7__15_), .S(SUMB_7__15_) );
  FA_X1 S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), .CO(
        CARRYB_7__16_), .S(SUMB_7__16_) );
  FA_X1 S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), .CO(
        CARRYB_7__17_), .S(SUMB_7__17_) );
  FA_X1 S2_7_18 ( .A(ab_7__18_), .B(CARRYB_6__18_), .CI(SUMB_6__19_), .CO(
        CARRYB_7__18_), .S(SUMB_7__18_) );
  FA_X1 S2_7_19 ( .A(ab_7__19_), .B(CARRYB_6__19_), .CI(SUMB_6__20_), .CO(
        CARRYB_7__19_), .S(SUMB_7__19_) );
  FA_X1 S2_7_20 ( .A(ab_7__20_), .B(CARRYB_6__20_), .CI(SUMB_6__21_), .CO(
        CARRYB_7__20_), .S(SUMB_7__20_) );
  FA_X1 S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), .CO(
        CARRYB_7__21_), .S(SUMB_7__21_) );
  FA_X1 S3_7_22 ( .A(ab_7__22_), .B(CARRYB_6__22_), .CI(ab_6__23_), .CO(
        CARRYB_7__22_), .S(SUMB_7__22_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S2_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  FA_X1 S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  FA_X1 S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  FA_X1 S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), .CO(
        CARRYB_6__10_), .S(SUMB_6__10_) );
  FA_X1 S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), .CO(
        CARRYB_6__11_), .S(SUMB_6__11_) );
  FA_X1 S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), .CO(
        CARRYB_6__12_), .S(SUMB_6__12_) );
  FA_X1 S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), .CO(
        CARRYB_6__13_), .S(SUMB_6__13_) );
  FA_X1 S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), .CO(
        CARRYB_6__14_), .S(SUMB_6__14_) );
  FA_X1 S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), .CO(
        CARRYB_6__15_), .S(SUMB_6__15_) );
  FA_X1 S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), .CO(
        CARRYB_6__16_), .S(SUMB_6__16_) );
  FA_X1 S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), .CO(
        CARRYB_6__17_), .S(SUMB_6__17_) );
  FA_X1 S2_6_18 ( .A(ab_6__18_), .B(CARRYB_5__18_), .CI(SUMB_5__19_), .CO(
        CARRYB_6__18_), .S(SUMB_6__18_) );
  FA_X1 S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), .CO(
        CARRYB_6__19_), .S(SUMB_6__19_) );
  FA_X1 S2_6_20 ( .A(ab_6__20_), .B(CARRYB_5__20_), .CI(SUMB_5__21_), .CO(
        CARRYB_6__20_), .S(SUMB_6__20_) );
  FA_X1 S2_6_21 ( .A(ab_6__21_), .B(CARRYB_5__21_), .CI(SUMB_5__22_), .CO(
        CARRYB_6__21_), .S(SUMB_6__21_) );
  FA_X1 S3_6_22 ( .A(ab_6__22_), .B(CARRYB_5__22_), .CI(ab_5__23_), .CO(
        CARRYB_6__22_), .S(SUMB_6__22_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  FA_X1 S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  FA_X1 S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  FA_X1 S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), .CO(
        CARRYB_5__10_), .S(SUMB_5__10_) );
  FA_X1 S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), .CO(
        CARRYB_5__11_), .S(SUMB_5__11_) );
  FA_X1 S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), .CO(
        CARRYB_5__12_), .S(SUMB_5__12_) );
  FA_X1 S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), .CO(
        CARRYB_5__13_), .S(SUMB_5__13_) );
  FA_X1 S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), .CO(
        CARRYB_5__14_), .S(SUMB_5__14_) );
  FA_X1 S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), .CO(
        CARRYB_5__15_), .S(SUMB_5__15_) );
  FA_X1 S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), .CO(
        CARRYB_5__16_), .S(SUMB_5__16_) );
  FA_X1 S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), .CO(
        CARRYB_5__17_), .S(SUMB_5__17_) );
  FA_X1 S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), .CO(
        CARRYB_5__18_), .S(SUMB_5__18_) );
  FA_X1 S2_5_19 ( .A(ab_5__19_), .B(CARRYB_4__19_), .CI(SUMB_4__20_), .CO(
        CARRYB_5__19_), .S(SUMB_5__19_) );
  FA_X1 S2_5_20 ( .A(ab_5__20_), .B(CARRYB_4__20_), .CI(SUMB_4__21_), .CO(
        CARRYB_5__20_), .S(SUMB_5__20_) );
  FA_X1 S2_5_21 ( .A(ab_5__21_), .B(CARRYB_4__21_), .CI(SUMB_4__22_), .CO(
        CARRYB_5__21_), .S(SUMB_5__21_) );
  FA_X1 S3_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(ab_4__23_), .CO(
        CARRYB_5__22_), .S(SUMB_5__22_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  FA_X1 S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  FA_X1 S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  FA_X1 S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), .CO(
        CARRYB_4__10_), .S(SUMB_4__10_) );
  FA_X1 S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), .CO(
        CARRYB_4__11_), .S(SUMB_4__11_) );
  FA_X1 S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), .CO(
        CARRYB_4__12_), .S(SUMB_4__12_) );
  FA_X1 S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), .CO(
        CARRYB_4__13_), .S(SUMB_4__13_) );
  FA_X1 S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), .CO(
        CARRYB_4__14_), .S(SUMB_4__14_) );
  FA_X1 S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), .CO(
        CARRYB_4__15_), .S(SUMB_4__15_) );
  FA_X1 S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), .CO(
        CARRYB_4__16_), .S(SUMB_4__16_) );
  FA_X1 S2_4_17 ( .A(ab_4__17_), .B(CARRYB_3__17_), .CI(SUMB_3__18_), .CO(
        CARRYB_4__17_), .S(SUMB_4__17_) );
  FA_X1 S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), .CO(
        CARRYB_4__18_), .S(SUMB_4__18_) );
  FA_X1 S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), .CO(
        CARRYB_4__19_), .S(SUMB_4__19_) );
  FA_X1 S2_4_20 ( .A(ab_4__20_), .B(CARRYB_3__20_), .CI(SUMB_3__21_), .CO(
        CARRYB_4__20_), .S(SUMB_4__20_) );
  FA_X1 S2_4_21 ( .A(ab_4__21_), .B(CARRYB_3__21_), .CI(SUMB_3__22_), .CO(
        CARRYB_4__21_), .S(SUMB_4__21_) );
  FA_X1 S3_4_22 ( .A(ab_4__22_), .B(CARRYB_3__22_), .CI(ab_3__23_), .CO(
        CARRYB_4__22_), .S(SUMB_4__22_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  FA_X1 S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  FA_X1 S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  FA_X1 S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), .CO(
        CARRYB_3__10_), .S(SUMB_3__10_) );
  FA_X1 S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), .CO(
        CARRYB_3__11_), .S(SUMB_3__11_) );
  FA_X1 S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), .CO(
        CARRYB_3__12_), .S(SUMB_3__12_) );
  FA_X1 S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), .CO(
        CARRYB_3__13_), .S(SUMB_3__13_) );
  FA_X1 S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), .CO(
        CARRYB_3__14_), .S(SUMB_3__14_) );
  FA_X1 S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), .CO(
        CARRYB_3__15_), .S(SUMB_3__15_) );
  FA_X1 S2_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(SUMB_2__17_), .CO(
        CARRYB_3__16_), .S(SUMB_3__16_) );
  FA_X1 S2_3_17 ( .A(ab_3__17_), .B(CARRYB_2__17_), .CI(SUMB_2__18_), .CO(
        CARRYB_3__17_), .S(SUMB_3__17_) );
  FA_X1 S2_3_18 ( .A(ab_3__18_), .B(CARRYB_2__18_), .CI(SUMB_2__19_), .CO(
        CARRYB_3__18_), .S(SUMB_3__18_) );
  FA_X1 S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), .CO(
        CARRYB_3__19_), .S(SUMB_3__19_) );
  FA_X1 S2_3_20 ( .A(ab_3__20_), .B(CARRYB_2__20_), .CI(SUMB_2__21_), .CO(
        CARRYB_3__20_), .S(SUMB_3__20_) );
  FA_X1 S2_3_21 ( .A(ab_3__21_), .B(CARRYB_2__21_), .CI(SUMB_2__22_), .CO(
        CARRYB_3__21_), .S(SUMB_3__21_) );
  FA_X1 S3_3_22 ( .A(ab_3__22_), .B(CARRYB_2__22_), .CI(ab_2__23_), .CO(
        CARRYB_3__22_), .S(SUMB_3__22_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S2_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(SUMB_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  FA_X1 S2_2_7 ( .A(ab_2__7_), .B(CARRYB_1__7_), .CI(SUMB_1__8_), .CO(
        CARRYB_2__7_), .S(SUMB_2__7_) );
  FA_X1 S2_2_8 ( .A(ab_2__8_), .B(CARRYB_1__8_), .CI(SUMB_1__9_), .CO(
        CARRYB_2__8_), .S(SUMB_2__8_) );
  FA_X1 S2_2_9 ( .A(ab_2__9_), .B(CARRYB_1__9_), .CI(SUMB_1__10_), .CO(
        CARRYB_2__9_), .S(SUMB_2__9_) );
  FA_X1 S2_2_10 ( .A(ab_2__10_), .B(CARRYB_1__10_), .CI(SUMB_1__11_), .CO(
        CARRYB_2__10_), .S(SUMB_2__10_) );
  FA_X1 S2_2_11 ( .A(ab_2__11_), .B(CARRYB_1__11_), .CI(SUMB_1__12_), .CO(
        CARRYB_2__11_), .S(SUMB_2__11_) );
  FA_X1 S2_2_12 ( .A(ab_2__12_), .B(CARRYB_1__12_), .CI(SUMB_1__13_), .CO(
        CARRYB_2__12_), .S(SUMB_2__12_) );
  FA_X1 S2_2_13 ( .A(ab_2__13_), .B(CARRYB_1__13_), .CI(SUMB_1__14_), .CO(
        CARRYB_2__13_), .S(SUMB_2__13_) );
  FA_X1 S2_2_14 ( .A(ab_2__14_), .B(CARRYB_1__14_), .CI(SUMB_1__15_), .CO(
        CARRYB_2__14_), .S(SUMB_2__14_) );
  FA_X1 S2_2_15 ( .A(ab_2__15_), .B(CARRYB_1__15_), .CI(SUMB_1__16_), .CO(
        CARRYB_2__15_), .S(SUMB_2__15_) );
  FA_X1 S2_2_16 ( .A(ab_2__16_), .B(CARRYB_1__16_), .CI(SUMB_1__17_), .CO(
        CARRYB_2__16_), .S(SUMB_2__16_) );
  FA_X1 S2_2_17 ( .A(ab_2__17_), .B(CARRYB_1__17_), .CI(SUMB_1__18_), .CO(
        CARRYB_2__17_), .S(SUMB_2__17_) );
  FA_X1 S2_2_18 ( .A(ab_2__18_), .B(CARRYB_1__18_), .CI(SUMB_1__19_), .CO(
        CARRYB_2__18_), .S(SUMB_2__18_) );
  FA_X1 S2_2_19 ( .A(ab_2__19_), .B(CARRYB_1__19_), .CI(SUMB_1__20_), .CO(
        CARRYB_2__19_), .S(SUMB_2__19_) );
  FA_X1 S2_2_20 ( .A(ab_2__20_), .B(CARRYB_1__20_), .CI(SUMB_1__21_), .CO(
        CARRYB_2__20_), .S(SUMB_2__20_) );
  FA_X1 S2_2_21 ( .A(ab_2__21_), .B(CARRYB_1__21_), .CI(SUMB_1__22_), .CO(
        CARRYB_2__21_), .S(SUMB_2__21_) );
  FA_X1 S3_2_22 ( .A(ab_2__22_), .B(CARRYB_1__22_), .CI(ab_1__23_), .CO(
        CARRYB_2__22_), .S(SUMB_2__22_) );
  iir_filter_DW01_add_5 FS_1 ( .A({A1_45_, A1_44_, A1_43_, A1_42_, A1_41_, 
        A1_40_, A1_39_, A1_38_, A1_37_, A1_36_, A1_35_, A1_34_, A1_33_, A1_32_, 
        A1_31_, A1_30_, A1_29_, A1_28_, A1_27_, A1_26_, A1_25_, A1_24_, A1_23_, 
        A1_22_, A1_21_, A1_20_, A1_19_, A1_18_, A1_17_, A1_16_, A1_15_, A1_14_, 
        A1_13_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, A1_5_, 
        A1_4_, A1_3_, A1_2_, A1_1_, A1_0_}), .B({A2_45_, A2_44_, A2_43_, 
        A2_42_, A2_41_, A2_40_, A2_39_, A2_38_, A2_37_, A2_36_, A2_35_, A2_34_, 
        A2_33_, A2_32_, A2_31_, A2_30_, A2_29_, A2_28_, A2_27_, A2_26_, A2_25_, 
        A2_24_, A2_23_, A2_22_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({PRODUCT[47], SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, PRODUCT[44:22], SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21}) );
  BUF_X1 U2 ( .A(QB), .Z(n1) );
  BUF_X1 U3 ( .A(QB), .Z(n2) );
  BUF_X1 U4 ( .A(QA), .Z(n3) );
  BUF_X1 U5 ( .A(QA), .Z(n4) );
  INV_X1 U6 ( .A(A[2]), .ZN(n36) );
  INV_X1 U7 ( .A(A[3]), .ZN(n35) );
  INV_X1 U8 ( .A(A[4]), .ZN(n34) );
  INV_X1 U9 ( .A(A[5]), .ZN(n33) );
  INV_X1 U10 ( .A(A[6]), .ZN(n32) );
  INV_X1 U11 ( .A(B[1]), .ZN(n18) );
  INV_X1 U12 ( .A(A[1]), .ZN(n40) );
  INV_X1 U13 ( .A(B[0]), .ZN(n29) );
  INV_X1 U14 ( .A(A[0]), .ZN(n51) );
  INV_X1 U15 ( .A(B[22]), .ZN(n15) );
  INV_X1 U16 ( .A(B[21]), .ZN(n16) );
  INV_X1 U17 ( .A(B[20]), .ZN(n17) );
  INV_X1 U18 ( .A(B[19]), .ZN(n19) );
  INV_X1 U19 ( .A(B[18]), .ZN(n20) );
  INV_X1 U20 ( .A(B[17]), .ZN(n21) );
  INV_X1 U21 ( .A(B[16]), .ZN(n22) );
  INV_X1 U22 ( .A(B[15]), .ZN(n23) );
  INV_X1 U23 ( .A(B[14]), .ZN(n24) );
  INV_X1 U24 ( .A(B[13]), .ZN(n25) );
  INV_X1 U25 ( .A(B[12]), .ZN(n26) );
  INV_X1 U26 ( .A(B[11]), .ZN(n27) );
  INV_X1 U27 ( .A(B[10]), .ZN(n28) );
  INV_X1 U28 ( .A(B[9]), .ZN(n7) );
  INV_X1 U29 ( .A(B[8]), .ZN(n8) );
  INV_X1 U30 ( .A(B[7]), .ZN(n9) );
  INV_X1 U31 ( .A(B[6]), .ZN(n10) );
  INV_X1 U32 ( .A(B[5]), .ZN(n11) );
  INV_X1 U33 ( .A(B[4]), .ZN(n12) );
  INV_X1 U34 ( .A(B[3]), .ZN(n13) );
  INV_X1 U35 ( .A(B[2]), .ZN(n14) );
  INV_X1 U36 ( .A(A[7]), .ZN(n31) );
  INV_X1 U37 ( .A(A[8]), .ZN(n30) );
  INV_X1 U38 ( .A(A[10]), .ZN(n50) );
  INV_X1 U39 ( .A(A[11]), .ZN(n49) );
  INV_X1 U40 ( .A(A[12]), .ZN(n48) );
  INV_X1 U41 ( .A(A[13]), .ZN(n47) );
  INV_X1 U42 ( .A(A[14]), .ZN(n46) );
  INV_X1 U43 ( .A(A[9]), .ZN(n6) );
  INV_X1 U44 ( .A(A[22]), .ZN(n37) );
  INV_X1 U45 ( .A(A[15]), .ZN(n45) );
  INV_X1 U46 ( .A(A[16]), .ZN(n44) );
  INV_X1 U47 ( .A(A[17]), .ZN(n43) );
  INV_X1 U48 ( .A(A[18]), .ZN(n42) );
  INV_X1 U49 ( .A(A[19]), .ZN(n41) );
  INV_X1 U50 ( .A(A[20]), .ZN(n39) );
  INV_X1 U51 ( .A(A[21]), .ZN(n38) );
  AND2_X1 U52 ( .A1(SUMB_23__23_), .A2(CARRYB_23__22_), .ZN(A2_45_) );
  XOR2_X1 U53 ( .A(CARRYB_23__22_), .B(SUMB_23__23_), .Z(A1_44_) );
  AND2_X1 U54 ( .A1(SUMB_23__22_), .A2(CARRYB_23__21_), .ZN(A2_44_) );
  XOR2_X1 U55 ( .A(CARRYB_23__21_), .B(SUMB_23__22_), .Z(A1_43_) );
  AND2_X1 U56 ( .A1(SUMB_23__21_), .A2(CARRYB_23__20_), .ZN(A2_43_) );
  XOR2_X1 U57 ( .A(CARRYB_23__20_), .B(SUMB_23__21_), .Z(A1_42_) );
  AND2_X1 U58 ( .A1(SUMB_23__20_), .A2(CARRYB_23__19_), .ZN(A2_42_) );
  XOR2_X1 U59 ( .A(CARRYB_23__19_), .B(SUMB_23__20_), .Z(A1_41_) );
  AND2_X1 U60 ( .A1(SUMB_23__19_), .A2(CARRYB_23__18_), .ZN(A2_41_) );
  XOR2_X1 U61 ( .A(CARRYB_23__18_), .B(SUMB_23__19_), .Z(A1_40_) );
  AND2_X1 U62 ( .A1(SUMB_23__18_), .A2(CARRYB_23__17_), .ZN(A2_40_) );
  XOR2_X1 U63 ( .A(CARRYB_23__17_), .B(SUMB_23__18_), .Z(A1_39_) );
  AND2_X1 U64 ( .A1(SUMB_23__17_), .A2(CARRYB_23__16_), .ZN(A2_39_) );
  XOR2_X1 U65 ( .A(CARRYB_23__16_), .B(SUMB_23__17_), .Z(A1_38_) );
  AND2_X1 U66 ( .A1(SUMB_23__16_), .A2(CARRYB_23__15_), .ZN(A2_38_) );
  XOR2_X1 U67 ( .A(CARRYB_23__15_), .B(SUMB_23__16_), .Z(A1_37_) );
  AND2_X1 U68 ( .A1(SUMB_23__15_), .A2(CARRYB_23__14_), .ZN(A2_37_) );
  XOR2_X1 U69 ( .A(CARRYB_23__14_), .B(SUMB_23__15_), .Z(A1_36_) );
  AND2_X1 U70 ( .A1(SUMB_23__14_), .A2(CARRYB_23__13_), .ZN(A2_36_) );
  XOR2_X1 U71 ( .A(CARRYB_23__13_), .B(SUMB_23__14_), .Z(A1_35_) );
  AND2_X1 U72 ( .A1(SUMB_23__13_), .A2(CARRYB_23__12_), .ZN(A2_35_) );
  XOR2_X1 U73 ( .A(CARRYB_23__12_), .B(SUMB_23__13_), .Z(A1_34_) );
  AND2_X1 U74 ( .A1(SUMB_23__12_), .A2(CARRYB_23__11_), .ZN(A2_34_) );
  XOR2_X1 U75 ( .A(CARRYB_23__11_), .B(SUMB_23__12_), .Z(A1_33_) );
  AND2_X1 U76 ( .A1(SUMB_23__11_), .A2(CARRYB_23__10_), .ZN(A2_33_) );
  XOR2_X1 U77 ( .A(CARRYB_23__10_), .B(SUMB_23__11_), .Z(A1_32_) );
  AND2_X1 U78 ( .A1(SUMB_23__10_), .A2(CARRYB_23__9_), .ZN(A2_32_) );
  XOR2_X1 U79 ( .A(CARRYB_23__9_), .B(SUMB_23__10_), .Z(A1_31_) );
  AND2_X1 U80 ( .A1(SUMB_23__9_), .A2(CARRYB_23__8_), .ZN(A2_31_) );
  XOR2_X1 U81 ( .A(CARRYB_23__8_), .B(SUMB_23__9_), .Z(A1_30_) );
  AND2_X1 U82 ( .A1(SUMB_23__8_), .A2(CARRYB_23__7_), .ZN(A2_30_) );
  XOR2_X1 U83 ( .A(CARRYB_23__7_), .B(SUMB_23__8_), .Z(A1_29_) );
  AND2_X1 U84 ( .A1(SUMB_23__7_), .A2(CARRYB_23__6_), .ZN(A2_29_) );
  XOR2_X1 U85 ( .A(CARRYB_23__6_), .B(SUMB_23__7_), .Z(A1_28_) );
  AND2_X1 U86 ( .A1(SUMB_23__6_), .A2(CARRYB_23__5_), .ZN(A2_28_) );
  XOR2_X1 U87 ( .A(CARRYB_23__5_), .B(SUMB_23__6_), .Z(A1_27_) );
  AND2_X1 U88 ( .A1(SUMB_23__5_), .A2(CARRYB_23__4_), .ZN(A2_27_) );
  XOR2_X1 U89 ( .A(CARRYB_23__4_), .B(SUMB_23__5_), .Z(A1_26_) );
  AND2_X1 U90 ( .A1(SUMB_23__4_), .A2(CARRYB_23__3_), .ZN(A2_26_) );
  XOR2_X1 U91 ( .A(CARRYB_23__3_), .B(SUMB_23__4_), .Z(A1_25_) );
  AND2_X1 U92 ( .A1(SUMB_23__3_), .A2(CARRYB_23__2_), .ZN(A2_25_) );
  XOR2_X1 U93 ( .A(CARRYB_23__2_), .B(SUMB_23__3_), .Z(A1_24_) );
  AND2_X1 U94 ( .A1(SUMB_23__2_), .A2(CARRYB_23__1_), .ZN(A2_24_) );
  XOR2_X1 U95 ( .A(CARRYB_23__1_), .B(SUMB_23__2_), .Z(A1_23_) );
  AND2_X1 U96 ( .A1(SUMB_23__1_), .A2(CARRYB_23__0_), .ZN(A2_23_) );
  XOR2_X1 U97 ( .A(CARRYB_23__0_), .B(SUMB_23__1_), .Z(A1_22_) );
  AND2_X1 U98 ( .A1(ab_1__22_), .A2(ab_0__23_), .ZN(CARRYB_1__22_) );
  XOR2_X1 U99 ( .A(ab_1__22_), .B(ab_0__23_), .Z(SUMB_1__22_) );
  AND2_X1 U100 ( .A1(ab_1__21_), .A2(ab_0__22_), .ZN(CARRYB_1__21_) );
  XOR2_X1 U101 ( .A(ab_1__21_), .B(ab_0__22_), .Z(SUMB_1__21_) );
  AND2_X1 U102 ( .A1(ab_1__20_), .A2(ab_0__21_), .ZN(CARRYB_1__20_) );
  XOR2_X1 U103 ( .A(ab_1__20_), .B(ab_0__21_), .Z(SUMB_1__20_) );
  AND2_X1 U104 ( .A1(ab_1__19_), .A2(ab_0__20_), .ZN(CARRYB_1__19_) );
  XOR2_X1 U105 ( .A(ab_1__19_), .B(ab_0__20_), .Z(SUMB_1__19_) );
  AND2_X1 U106 ( .A1(ab_1__18_), .A2(ab_0__19_), .ZN(CARRYB_1__18_) );
  XOR2_X1 U107 ( .A(ab_1__18_), .B(ab_0__19_), .Z(SUMB_1__18_) );
  AND2_X1 U108 ( .A1(ab_1__17_), .A2(ab_0__18_), .ZN(CARRYB_1__17_) );
  XOR2_X1 U109 ( .A(ab_1__17_), .B(ab_0__18_), .Z(SUMB_1__17_) );
  AND2_X1 U110 ( .A1(ab_1__16_), .A2(ab_0__17_), .ZN(CARRYB_1__16_) );
  XOR2_X1 U111 ( .A(ab_1__16_), .B(ab_0__17_), .Z(SUMB_1__16_) );
  AND2_X1 U112 ( .A1(ab_1__15_), .A2(ab_0__16_), .ZN(CARRYB_1__15_) );
  XOR2_X1 U113 ( .A(ab_1__15_), .B(ab_0__16_), .Z(SUMB_1__15_) );
  AND2_X1 U114 ( .A1(ab_1__14_), .A2(ab_0__15_), .ZN(CARRYB_1__14_) );
  XOR2_X1 U115 ( .A(ab_1__14_), .B(ab_0__15_), .Z(SUMB_1__14_) );
  AND2_X1 U116 ( .A1(ab_1__13_), .A2(ab_0__14_), .ZN(CARRYB_1__13_) );
  XOR2_X1 U117 ( .A(ab_1__13_), .B(ab_0__14_), .Z(SUMB_1__13_) );
  AND2_X1 U118 ( .A1(ab_1__12_), .A2(ab_0__13_), .ZN(CARRYB_1__12_) );
  XOR2_X1 U119 ( .A(ab_1__12_), .B(ab_0__13_), .Z(SUMB_1__12_) );
  AND2_X1 U120 ( .A1(ab_1__11_), .A2(ab_0__12_), .ZN(CARRYB_1__11_) );
  XOR2_X1 U121 ( .A(ab_1__11_), .B(ab_0__12_), .Z(SUMB_1__11_) );
  AND2_X1 U122 ( .A1(ab_1__10_), .A2(ab_0__11_), .ZN(CARRYB_1__10_) );
  XOR2_X1 U123 ( .A(ab_1__10_), .B(ab_0__11_), .Z(SUMB_1__10_) );
  AND2_X1 U124 ( .A1(ab_1__9_), .A2(ab_0__10_), .ZN(CARRYB_1__9_) );
  XOR2_X1 U125 ( .A(ab_1__9_), .B(ab_0__10_), .Z(SUMB_1__9_) );
  AND2_X1 U126 ( .A1(ab_1__8_), .A2(ab_0__9_), .ZN(CARRYB_1__8_) );
  XOR2_X1 U127 ( .A(ab_1__8_), .B(ab_0__9_), .Z(SUMB_1__8_) );
  AND2_X1 U128 ( .A1(ab_1__7_), .A2(ab_0__8_), .ZN(CARRYB_1__7_) );
  XOR2_X1 U129 ( .A(ab_1__7_), .B(ab_0__8_), .Z(SUMB_1__7_) );
  AND2_X1 U130 ( .A1(ab_1__6_), .A2(ab_0__7_), .ZN(CARRYB_1__6_) );
  XOR2_X1 U131 ( .A(ab_1__6_), .B(ab_0__7_), .Z(SUMB_1__6_) );
  AND2_X1 U132 ( .A1(ab_1__5_), .A2(ab_0__6_), .ZN(CARRYB_1__5_) );
  XOR2_X1 U133 ( .A(ab_1__5_), .B(ab_0__6_), .Z(SUMB_1__5_) );
  AND2_X1 U134 ( .A1(ab_1__4_), .A2(ab_0__5_), .ZN(CARRYB_1__4_) );
  XOR2_X1 U135 ( .A(ab_1__4_), .B(ab_0__5_), .Z(SUMB_1__4_) );
  AND2_X1 U136 ( .A1(ab_1__3_), .A2(ab_0__4_), .ZN(CARRYB_1__3_) );
  XOR2_X1 U137 ( .A(ab_1__3_), .B(ab_0__4_), .Z(SUMB_1__3_) );
  AND2_X1 U138 ( .A1(ab_1__2_), .A2(ab_0__3_), .ZN(CARRYB_1__2_) );
  XOR2_X1 U139 ( .A(ab_1__2_), .B(ab_0__3_), .Z(SUMB_1__2_) );
  AND2_X1 U140 ( .A1(ab_1__1_), .A2(ab_0__2_), .ZN(CARRYB_1__1_) );
  XOR2_X1 U141 ( .A(ab_1__1_), .B(ab_0__2_), .Z(SUMB_1__1_) );
  NOR2_X1 U142 ( .A1(n6), .A2(n7), .ZN(ab_9__9_) );
  NOR2_X1 U143 ( .A1(n6), .A2(n8), .ZN(ab_9__8_) );
  NOR2_X1 U144 ( .A1(n6), .A2(n9), .ZN(ab_9__7_) );
  NOR2_X1 U145 ( .A1(n6), .A2(n10), .ZN(ab_9__6_) );
  NOR2_X1 U146 ( .A1(n6), .A2(n11), .ZN(ab_9__5_) );
  NOR2_X1 U147 ( .A1(n6), .A2(n12), .ZN(ab_9__4_) );
  NOR2_X1 U148 ( .A1(n6), .A2(n13), .ZN(ab_9__3_) );
  NOR2_X1 U149 ( .A1(n6), .A2(n14), .ZN(ab_9__2_) );
  NOR2_X1 U150 ( .A1(A[9]), .A2(n1), .ZN(ab_9__23_) );
  NOR2_X1 U151 ( .A1(n6), .A2(n15), .ZN(ab_9__22_) );
  NOR2_X1 U152 ( .A1(n6), .A2(n16), .ZN(ab_9__21_) );
  NOR2_X1 U153 ( .A1(n6), .A2(n17), .ZN(ab_9__20_) );
  NOR2_X1 U154 ( .A1(n6), .A2(n18), .ZN(ab_9__1_) );
  NOR2_X1 U155 ( .A1(n6), .A2(n19), .ZN(ab_9__19_) );
  NOR2_X1 U156 ( .A1(n6), .A2(n20), .ZN(ab_9__18_) );
  NOR2_X1 U157 ( .A1(n6), .A2(n21), .ZN(ab_9__17_) );
  NOR2_X1 U158 ( .A1(n6), .A2(n22), .ZN(ab_9__16_) );
  NOR2_X1 U159 ( .A1(n6), .A2(n23), .ZN(ab_9__15_) );
  NOR2_X1 U160 ( .A1(n6), .A2(n24), .ZN(ab_9__14_) );
  NOR2_X1 U161 ( .A1(n6), .A2(n25), .ZN(ab_9__13_) );
  NOR2_X1 U162 ( .A1(n6), .A2(n26), .ZN(ab_9__12_) );
  NOR2_X1 U163 ( .A1(n6), .A2(n27), .ZN(ab_9__11_) );
  NOR2_X1 U164 ( .A1(n6), .A2(n28), .ZN(ab_9__10_) );
  NOR2_X1 U165 ( .A1(n6), .A2(n29), .ZN(ab_9__0_) );
  NOR2_X1 U166 ( .A1(n7), .A2(n30), .ZN(ab_8__9_) );
  NOR2_X1 U167 ( .A1(n8), .A2(n30), .ZN(ab_8__8_) );
  NOR2_X1 U168 ( .A1(n9), .A2(n30), .ZN(ab_8__7_) );
  NOR2_X1 U169 ( .A1(n10), .A2(n30), .ZN(ab_8__6_) );
  NOR2_X1 U170 ( .A1(n11), .A2(n30), .ZN(ab_8__5_) );
  NOR2_X1 U171 ( .A1(n12), .A2(n30), .ZN(ab_8__4_) );
  NOR2_X1 U172 ( .A1(n13), .A2(n30), .ZN(ab_8__3_) );
  NOR2_X1 U173 ( .A1(n14), .A2(n30), .ZN(ab_8__2_) );
  NOR2_X1 U174 ( .A1(A[8]), .A2(n1), .ZN(ab_8__23_) );
  NOR2_X1 U175 ( .A1(n15), .A2(n30), .ZN(ab_8__22_) );
  NOR2_X1 U176 ( .A1(n16), .A2(n30), .ZN(ab_8__21_) );
  NOR2_X1 U177 ( .A1(n17), .A2(n30), .ZN(ab_8__20_) );
  NOR2_X1 U178 ( .A1(n18), .A2(n30), .ZN(ab_8__1_) );
  NOR2_X1 U179 ( .A1(n19), .A2(n30), .ZN(ab_8__19_) );
  NOR2_X1 U180 ( .A1(n20), .A2(n30), .ZN(ab_8__18_) );
  NOR2_X1 U181 ( .A1(n21), .A2(n30), .ZN(ab_8__17_) );
  NOR2_X1 U182 ( .A1(n22), .A2(n30), .ZN(ab_8__16_) );
  NOR2_X1 U183 ( .A1(n23), .A2(n30), .ZN(ab_8__15_) );
  NOR2_X1 U184 ( .A1(n24), .A2(n30), .ZN(ab_8__14_) );
  NOR2_X1 U185 ( .A1(n25), .A2(n30), .ZN(ab_8__13_) );
  NOR2_X1 U186 ( .A1(n26), .A2(n30), .ZN(ab_8__12_) );
  NOR2_X1 U187 ( .A1(n27), .A2(n30), .ZN(ab_8__11_) );
  NOR2_X1 U188 ( .A1(n28), .A2(n30), .ZN(ab_8__10_) );
  NOR2_X1 U189 ( .A1(n29), .A2(n30), .ZN(ab_8__0_) );
  NOR2_X1 U190 ( .A1(n7), .A2(n31), .ZN(ab_7__9_) );
  NOR2_X1 U191 ( .A1(n8), .A2(n31), .ZN(ab_7__8_) );
  NOR2_X1 U192 ( .A1(n9), .A2(n31), .ZN(ab_7__7_) );
  NOR2_X1 U193 ( .A1(n10), .A2(n31), .ZN(ab_7__6_) );
  NOR2_X1 U194 ( .A1(n11), .A2(n31), .ZN(ab_7__5_) );
  NOR2_X1 U195 ( .A1(n12), .A2(n31), .ZN(ab_7__4_) );
  NOR2_X1 U196 ( .A1(n13), .A2(n31), .ZN(ab_7__3_) );
  NOR2_X1 U197 ( .A1(n14), .A2(n31), .ZN(ab_7__2_) );
  NOR2_X1 U198 ( .A1(A[7]), .A2(n1), .ZN(ab_7__23_) );
  NOR2_X1 U199 ( .A1(n15), .A2(n31), .ZN(ab_7__22_) );
  NOR2_X1 U200 ( .A1(n16), .A2(n31), .ZN(ab_7__21_) );
  NOR2_X1 U201 ( .A1(n17), .A2(n31), .ZN(ab_7__20_) );
  NOR2_X1 U202 ( .A1(n18), .A2(n31), .ZN(ab_7__1_) );
  NOR2_X1 U203 ( .A1(n19), .A2(n31), .ZN(ab_7__19_) );
  NOR2_X1 U204 ( .A1(n20), .A2(n31), .ZN(ab_7__18_) );
  NOR2_X1 U205 ( .A1(n21), .A2(n31), .ZN(ab_7__17_) );
  NOR2_X1 U206 ( .A1(n22), .A2(n31), .ZN(ab_7__16_) );
  NOR2_X1 U207 ( .A1(n23), .A2(n31), .ZN(ab_7__15_) );
  NOR2_X1 U208 ( .A1(n24), .A2(n31), .ZN(ab_7__14_) );
  NOR2_X1 U209 ( .A1(n25), .A2(n31), .ZN(ab_7__13_) );
  NOR2_X1 U210 ( .A1(n26), .A2(n31), .ZN(ab_7__12_) );
  NOR2_X1 U211 ( .A1(n27), .A2(n31), .ZN(ab_7__11_) );
  NOR2_X1 U212 ( .A1(n28), .A2(n31), .ZN(ab_7__10_) );
  NOR2_X1 U213 ( .A1(n29), .A2(n31), .ZN(ab_7__0_) );
  NOR2_X1 U214 ( .A1(n7), .A2(n32), .ZN(ab_6__9_) );
  NOR2_X1 U215 ( .A1(n8), .A2(n32), .ZN(ab_6__8_) );
  NOR2_X1 U216 ( .A1(n9), .A2(n32), .ZN(ab_6__7_) );
  NOR2_X1 U217 ( .A1(n10), .A2(n32), .ZN(ab_6__6_) );
  NOR2_X1 U218 ( .A1(n11), .A2(n32), .ZN(ab_6__5_) );
  NOR2_X1 U219 ( .A1(n12), .A2(n32), .ZN(ab_6__4_) );
  NOR2_X1 U220 ( .A1(n13), .A2(n32), .ZN(ab_6__3_) );
  NOR2_X1 U221 ( .A1(n14), .A2(n32), .ZN(ab_6__2_) );
  NOR2_X1 U222 ( .A1(A[6]), .A2(n1), .ZN(ab_6__23_) );
  NOR2_X1 U223 ( .A1(n15), .A2(n32), .ZN(ab_6__22_) );
  NOR2_X1 U224 ( .A1(n16), .A2(n32), .ZN(ab_6__21_) );
  NOR2_X1 U225 ( .A1(n17), .A2(n32), .ZN(ab_6__20_) );
  NOR2_X1 U226 ( .A1(n18), .A2(n32), .ZN(ab_6__1_) );
  NOR2_X1 U227 ( .A1(n19), .A2(n32), .ZN(ab_6__19_) );
  NOR2_X1 U228 ( .A1(n20), .A2(n32), .ZN(ab_6__18_) );
  NOR2_X1 U229 ( .A1(n21), .A2(n32), .ZN(ab_6__17_) );
  NOR2_X1 U230 ( .A1(n22), .A2(n32), .ZN(ab_6__16_) );
  NOR2_X1 U231 ( .A1(n23), .A2(n32), .ZN(ab_6__15_) );
  NOR2_X1 U232 ( .A1(n24), .A2(n32), .ZN(ab_6__14_) );
  NOR2_X1 U233 ( .A1(n25), .A2(n32), .ZN(ab_6__13_) );
  NOR2_X1 U234 ( .A1(n26), .A2(n32), .ZN(ab_6__12_) );
  NOR2_X1 U235 ( .A1(n27), .A2(n32), .ZN(ab_6__11_) );
  NOR2_X1 U236 ( .A1(n28), .A2(n32), .ZN(ab_6__10_) );
  NOR2_X1 U237 ( .A1(n29), .A2(n32), .ZN(ab_6__0_) );
  NOR2_X1 U238 ( .A1(n7), .A2(n33), .ZN(ab_5__9_) );
  NOR2_X1 U239 ( .A1(n8), .A2(n33), .ZN(ab_5__8_) );
  NOR2_X1 U240 ( .A1(n9), .A2(n33), .ZN(ab_5__7_) );
  NOR2_X1 U241 ( .A1(n10), .A2(n33), .ZN(ab_5__6_) );
  NOR2_X1 U242 ( .A1(n11), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U243 ( .A1(n12), .A2(n33), .ZN(ab_5__4_) );
  NOR2_X1 U244 ( .A1(n13), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U245 ( .A1(n14), .A2(n33), .ZN(ab_5__2_) );
  NOR2_X1 U246 ( .A1(A[5]), .A2(n1), .ZN(ab_5__23_) );
  NOR2_X1 U247 ( .A1(n15), .A2(n33), .ZN(ab_5__22_) );
  NOR2_X1 U248 ( .A1(n16), .A2(n33), .ZN(ab_5__21_) );
  NOR2_X1 U249 ( .A1(n17), .A2(n33), .ZN(ab_5__20_) );
  NOR2_X1 U250 ( .A1(n18), .A2(n33), .ZN(ab_5__1_) );
  NOR2_X1 U251 ( .A1(n19), .A2(n33), .ZN(ab_5__19_) );
  NOR2_X1 U252 ( .A1(n20), .A2(n33), .ZN(ab_5__18_) );
  NOR2_X1 U253 ( .A1(n21), .A2(n33), .ZN(ab_5__17_) );
  NOR2_X1 U254 ( .A1(n22), .A2(n33), .ZN(ab_5__16_) );
  NOR2_X1 U255 ( .A1(n23), .A2(n33), .ZN(ab_5__15_) );
  NOR2_X1 U256 ( .A1(n24), .A2(n33), .ZN(ab_5__14_) );
  NOR2_X1 U257 ( .A1(n25), .A2(n33), .ZN(ab_5__13_) );
  NOR2_X1 U258 ( .A1(n26), .A2(n33), .ZN(ab_5__12_) );
  NOR2_X1 U259 ( .A1(n27), .A2(n33), .ZN(ab_5__11_) );
  NOR2_X1 U260 ( .A1(n28), .A2(n33), .ZN(ab_5__10_) );
  NOR2_X1 U261 ( .A1(n29), .A2(n33), .ZN(ab_5__0_) );
  NOR2_X1 U262 ( .A1(n7), .A2(n34), .ZN(ab_4__9_) );
  NOR2_X1 U263 ( .A1(n8), .A2(n34), .ZN(ab_4__8_) );
  NOR2_X1 U264 ( .A1(n9), .A2(n34), .ZN(ab_4__7_) );
  NOR2_X1 U265 ( .A1(n10), .A2(n34), .ZN(ab_4__6_) );
  NOR2_X1 U266 ( .A1(n11), .A2(n34), .ZN(ab_4__5_) );
  NOR2_X1 U267 ( .A1(n12), .A2(n34), .ZN(ab_4__4_) );
  NOR2_X1 U268 ( .A1(n13), .A2(n34), .ZN(ab_4__3_) );
  NOR2_X1 U269 ( .A1(n14), .A2(n34), .ZN(ab_4__2_) );
  NOR2_X1 U270 ( .A1(A[4]), .A2(n1), .ZN(ab_4__23_) );
  NOR2_X1 U271 ( .A1(n15), .A2(n34), .ZN(ab_4__22_) );
  NOR2_X1 U272 ( .A1(n16), .A2(n34), .ZN(ab_4__21_) );
  NOR2_X1 U273 ( .A1(n17), .A2(n34), .ZN(ab_4__20_) );
  NOR2_X1 U274 ( .A1(n18), .A2(n34), .ZN(ab_4__1_) );
  NOR2_X1 U275 ( .A1(n19), .A2(n34), .ZN(ab_4__19_) );
  NOR2_X1 U276 ( .A1(n20), .A2(n34), .ZN(ab_4__18_) );
  NOR2_X1 U277 ( .A1(n21), .A2(n34), .ZN(ab_4__17_) );
  NOR2_X1 U278 ( .A1(n22), .A2(n34), .ZN(ab_4__16_) );
  NOR2_X1 U279 ( .A1(n23), .A2(n34), .ZN(ab_4__15_) );
  NOR2_X1 U280 ( .A1(n24), .A2(n34), .ZN(ab_4__14_) );
  NOR2_X1 U281 ( .A1(n25), .A2(n34), .ZN(ab_4__13_) );
  NOR2_X1 U282 ( .A1(n26), .A2(n34), .ZN(ab_4__12_) );
  NOR2_X1 U283 ( .A1(n27), .A2(n34), .ZN(ab_4__11_) );
  NOR2_X1 U284 ( .A1(n28), .A2(n34), .ZN(ab_4__10_) );
  NOR2_X1 U285 ( .A1(n29), .A2(n34), .ZN(ab_4__0_) );
  NOR2_X1 U286 ( .A1(n7), .A2(n35), .ZN(ab_3__9_) );
  NOR2_X1 U287 ( .A1(n8), .A2(n35), .ZN(ab_3__8_) );
  NOR2_X1 U288 ( .A1(n9), .A2(n35), .ZN(ab_3__7_) );
  NOR2_X1 U289 ( .A1(n10), .A2(n35), .ZN(ab_3__6_) );
  NOR2_X1 U290 ( .A1(n11), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U291 ( .A1(n12), .A2(n35), .ZN(ab_3__4_) );
  NOR2_X1 U292 ( .A1(n13), .A2(n35), .ZN(ab_3__3_) );
  NOR2_X1 U293 ( .A1(n14), .A2(n35), .ZN(ab_3__2_) );
  NOR2_X1 U294 ( .A1(A[3]), .A2(n1), .ZN(ab_3__23_) );
  NOR2_X1 U295 ( .A1(n15), .A2(n35), .ZN(ab_3__22_) );
  NOR2_X1 U296 ( .A1(n16), .A2(n35), .ZN(ab_3__21_) );
  NOR2_X1 U297 ( .A1(n17), .A2(n35), .ZN(ab_3__20_) );
  NOR2_X1 U298 ( .A1(n18), .A2(n35), .ZN(ab_3__1_) );
  NOR2_X1 U299 ( .A1(n19), .A2(n35), .ZN(ab_3__19_) );
  NOR2_X1 U300 ( .A1(n20), .A2(n35), .ZN(ab_3__18_) );
  NOR2_X1 U301 ( .A1(n21), .A2(n35), .ZN(ab_3__17_) );
  NOR2_X1 U302 ( .A1(n22), .A2(n35), .ZN(ab_3__16_) );
  NOR2_X1 U303 ( .A1(n23), .A2(n35), .ZN(ab_3__15_) );
  NOR2_X1 U304 ( .A1(n24), .A2(n35), .ZN(ab_3__14_) );
  NOR2_X1 U305 ( .A1(n25), .A2(n35), .ZN(ab_3__13_) );
  NOR2_X1 U306 ( .A1(n26), .A2(n35), .ZN(ab_3__12_) );
  NOR2_X1 U307 ( .A1(n27), .A2(n35), .ZN(ab_3__11_) );
  NOR2_X1 U308 ( .A1(n28), .A2(n35), .ZN(ab_3__10_) );
  NOR2_X1 U309 ( .A1(n29), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U310 ( .A1(n7), .A2(n36), .ZN(ab_2__9_) );
  NOR2_X1 U311 ( .A1(n8), .A2(n36), .ZN(ab_2__8_) );
  NOR2_X1 U312 ( .A1(n9), .A2(n36), .ZN(ab_2__7_) );
  NOR2_X1 U313 ( .A1(n10), .A2(n36), .ZN(ab_2__6_) );
  NOR2_X1 U314 ( .A1(n11), .A2(n36), .ZN(ab_2__5_) );
  NOR2_X1 U315 ( .A1(n12), .A2(n36), .ZN(ab_2__4_) );
  NOR2_X1 U316 ( .A1(n13), .A2(n36), .ZN(ab_2__3_) );
  NOR2_X1 U317 ( .A1(n14), .A2(n36), .ZN(ab_2__2_) );
  NOR2_X1 U318 ( .A1(A[2]), .A2(n1), .ZN(ab_2__23_) );
  NOR2_X1 U319 ( .A1(n15), .A2(n36), .ZN(ab_2__22_) );
  NOR2_X1 U320 ( .A1(n16), .A2(n36), .ZN(ab_2__21_) );
  NOR2_X1 U321 ( .A1(n17), .A2(n36), .ZN(ab_2__20_) );
  NOR2_X1 U322 ( .A1(n18), .A2(n36), .ZN(ab_2__1_) );
  NOR2_X1 U323 ( .A1(n19), .A2(n36), .ZN(ab_2__19_) );
  NOR2_X1 U324 ( .A1(n20), .A2(n36), .ZN(ab_2__18_) );
  NOR2_X1 U325 ( .A1(n21), .A2(n36), .ZN(ab_2__17_) );
  NOR2_X1 U326 ( .A1(n22), .A2(n36), .ZN(ab_2__16_) );
  NOR2_X1 U327 ( .A1(n23), .A2(n36), .ZN(ab_2__15_) );
  NOR2_X1 U328 ( .A1(n24), .A2(n36), .ZN(ab_2__14_) );
  NOR2_X1 U329 ( .A1(n25), .A2(n36), .ZN(ab_2__13_) );
  NOR2_X1 U330 ( .A1(n26), .A2(n36), .ZN(ab_2__12_) );
  NOR2_X1 U331 ( .A1(n27), .A2(n36), .ZN(ab_2__11_) );
  NOR2_X1 U332 ( .A1(n28), .A2(n36), .ZN(ab_2__10_) );
  NOR2_X1 U333 ( .A1(n29), .A2(n36), .ZN(ab_2__0_) );
  NOR2_X1 U334 ( .A1(B[9]), .A2(n4), .ZN(ab_23__9_) );
  NOR2_X1 U335 ( .A1(B[8]), .A2(n4), .ZN(ab_23__8_) );
  NOR2_X1 U336 ( .A1(B[7]), .A2(n4), .ZN(ab_23__7_) );
  NOR2_X1 U337 ( .A1(B[6]), .A2(n4), .ZN(ab_23__6_) );
  NOR2_X1 U338 ( .A1(B[5]), .A2(n3), .ZN(ab_23__5_) );
  NOR2_X1 U339 ( .A1(B[4]), .A2(n3), .ZN(ab_23__4_) );
  NOR2_X1 U340 ( .A1(B[3]), .A2(n3), .ZN(ab_23__3_) );
  NOR2_X1 U341 ( .A1(B[2]), .A2(n3), .ZN(ab_23__2_) );
  NOR2_X1 U342 ( .A1(n1), .A2(n3), .ZN(ab_23__23_) );
  NOR2_X1 U343 ( .A1(B[22]), .A2(n3), .ZN(ab_23__22_) );
  NOR2_X1 U344 ( .A1(B[21]), .A2(n3), .ZN(ab_23__21_) );
  NOR2_X1 U345 ( .A1(B[20]), .A2(n3), .ZN(ab_23__20_) );
  NOR2_X1 U346 ( .A1(B[1]), .A2(n3), .ZN(ab_23__1_) );
  NOR2_X1 U347 ( .A1(B[19]), .A2(n3), .ZN(ab_23__19_) );
  NOR2_X1 U348 ( .A1(B[18]), .A2(n3), .ZN(ab_23__18_) );
  NOR2_X1 U349 ( .A1(B[17]), .A2(n3), .ZN(ab_23__17_) );
  NOR2_X1 U350 ( .A1(B[16]), .A2(n3), .ZN(ab_23__16_) );
  NOR2_X1 U351 ( .A1(B[15]), .A2(n3), .ZN(ab_23__15_) );
  NOR2_X1 U352 ( .A1(B[14]), .A2(n3), .ZN(ab_23__14_) );
  NOR2_X1 U353 ( .A1(B[13]), .A2(n3), .ZN(ab_23__13_) );
  NOR2_X1 U354 ( .A1(B[12]), .A2(n3), .ZN(ab_23__12_) );
  NOR2_X1 U355 ( .A1(B[11]), .A2(n3), .ZN(ab_23__11_) );
  NOR2_X1 U356 ( .A1(B[10]), .A2(n3), .ZN(ab_23__10_) );
  NOR2_X1 U357 ( .A1(B[0]), .A2(n3), .ZN(ab_23__0_) );
  NOR2_X1 U358 ( .A1(n7), .A2(n37), .ZN(ab_22__9_) );
  NOR2_X1 U359 ( .A1(n8), .A2(n37), .ZN(ab_22__8_) );
  NOR2_X1 U360 ( .A1(n9), .A2(n37), .ZN(ab_22__7_) );
  NOR2_X1 U361 ( .A1(n10), .A2(n37), .ZN(ab_22__6_) );
  NOR2_X1 U362 ( .A1(n11), .A2(n37), .ZN(ab_22__5_) );
  NOR2_X1 U363 ( .A1(n12), .A2(n37), .ZN(ab_22__4_) );
  NOR2_X1 U364 ( .A1(n13), .A2(n37), .ZN(ab_22__3_) );
  NOR2_X1 U365 ( .A1(n14), .A2(n37), .ZN(ab_22__2_) );
  NOR2_X1 U366 ( .A1(A[22]), .A2(n1), .ZN(ab_22__23_) );
  NOR2_X1 U367 ( .A1(n15), .A2(n37), .ZN(ab_22__22_) );
  NOR2_X1 U368 ( .A1(n16), .A2(n37), .ZN(ab_22__21_) );
  NOR2_X1 U369 ( .A1(n17), .A2(n37), .ZN(ab_22__20_) );
  NOR2_X1 U370 ( .A1(n18), .A2(n37), .ZN(ab_22__1_) );
  NOR2_X1 U371 ( .A1(n19), .A2(n37), .ZN(ab_22__19_) );
  NOR2_X1 U372 ( .A1(n20), .A2(n37), .ZN(ab_22__18_) );
  NOR2_X1 U373 ( .A1(n21), .A2(n37), .ZN(ab_22__17_) );
  NOR2_X1 U374 ( .A1(n22), .A2(n37), .ZN(ab_22__16_) );
  NOR2_X1 U375 ( .A1(n23), .A2(n37), .ZN(ab_22__15_) );
  NOR2_X1 U376 ( .A1(n24), .A2(n37), .ZN(ab_22__14_) );
  NOR2_X1 U377 ( .A1(n25), .A2(n37), .ZN(ab_22__13_) );
  NOR2_X1 U378 ( .A1(n26), .A2(n37), .ZN(ab_22__12_) );
  NOR2_X1 U379 ( .A1(n27), .A2(n37), .ZN(ab_22__11_) );
  NOR2_X1 U380 ( .A1(n28), .A2(n37), .ZN(ab_22__10_) );
  NOR2_X1 U381 ( .A1(n29), .A2(n37), .ZN(ab_22__0_) );
  NOR2_X1 U382 ( .A1(n7), .A2(n38), .ZN(ab_21__9_) );
  NOR2_X1 U383 ( .A1(n8), .A2(n38), .ZN(ab_21__8_) );
  NOR2_X1 U384 ( .A1(n9), .A2(n38), .ZN(ab_21__7_) );
  NOR2_X1 U385 ( .A1(n10), .A2(n38), .ZN(ab_21__6_) );
  NOR2_X1 U386 ( .A1(n11), .A2(n38), .ZN(ab_21__5_) );
  NOR2_X1 U387 ( .A1(n12), .A2(n38), .ZN(ab_21__4_) );
  NOR2_X1 U388 ( .A1(n13), .A2(n38), .ZN(ab_21__3_) );
  NOR2_X1 U389 ( .A1(n14), .A2(n38), .ZN(ab_21__2_) );
  NOR2_X1 U390 ( .A1(A[21]), .A2(n1), .ZN(ab_21__23_) );
  NOR2_X1 U391 ( .A1(n15), .A2(n38), .ZN(ab_21__22_) );
  NOR2_X1 U392 ( .A1(n16), .A2(n38), .ZN(ab_21__21_) );
  NOR2_X1 U393 ( .A1(n17), .A2(n38), .ZN(ab_21__20_) );
  NOR2_X1 U394 ( .A1(n18), .A2(n38), .ZN(ab_21__1_) );
  NOR2_X1 U395 ( .A1(n19), .A2(n38), .ZN(ab_21__19_) );
  NOR2_X1 U396 ( .A1(n20), .A2(n38), .ZN(ab_21__18_) );
  NOR2_X1 U397 ( .A1(n21), .A2(n38), .ZN(ab_21__17_) );
  NOR2_X1 U398 ( .A1(n22), .A2(n38), .ZN(ab_21__16_) );
  NOR2_X1 U399 ( .A1(n23), .A2(n38), .ZN(ab_21__15_) );
  NOR2_X1 U400 ( .A1(n24), .A2(n38), .ZN(ab_21__14_) );
  NOR2_X1 U401 ( .A1(n25), .A2(n38), .ZN(ab_21__13_) );
  NOR2_X1 U402 ( .A1(n26), .A2(n38), .ZN(ab_21__12_) );
  NOR2_X1 U403 ( .A1(n27), .A2(n38), .ZN(ab_21__11_) );
  NOR2_X1 U404 ( .A1(n28), .A2(n38), .ZN(ab_21__10_) );
  NOR2_X1 U405 ( .A1(n29), .A2(n38), .ZN(ab_21__0_) );
  NOR2_X1 U406 ( .A1(n7), .A2(n39), .ZN(ab_20__9_) );
  NOR2_X1 U407 ( .A1(n8), .A2(n39), .ZN(ab_20__8_) );
  NOR2_X1 U408 ( .A1(n9), .A2(n39), .ZN(ab_20__7_) );
  NOR2_X1 U409 ( .A1(n10), .A2(n39), .ZN(ab_20__6_) );
  NOR2_X1 U410 ( .A1(n11), .A2(n39), .ZN(ab_20__5_) );
  NOR2_X1 U411 ( .A1(n12), .A2(n39), .ZN(ab_20__4_) );
  NOR2_X1 U412 ( .A1(n13), .A2(n39), .ZN(ab_20__3_) );
  NOR2_X1 U413 ( .A1(n14), .A2(n39), .ZN(ab_20__2_) );
  NOR2_X1 U414 ( .A1(A[20]), .A2(n1), .ZN(ab_20__23_) );
  NOR2_X1 U415 ( .A1(n15), .A2(n39), .ZN(ab_20__22_) );
  NOR2_X1 U416 ( .A1(n16), .A2(n39), .ZN(ab_20__21_) );
  NOR2_X1 U417 ( .A1(n17), .A2(n39), .ZN(ab_20__20_) );
  NOR2_X1 U418 ( .A1(n18), .A2(n39), .ZN(ab_20__1_) );
  NOR2_X1 U419 ( .A1(n19), .A2(n39), .ZN(ab_20__19_) );
  NOR2_X1 U420 ( .A1(n20), .A2(n39), .ZN(ab_20__18_) );
  NOR2_X1 U421 ( .A1(n21), .A2(n39), .ZN(ab_20__17_) );
  NOR2_X1 U422 ( .A1(n22), .A2(n39), .ZN(ab_20__16_) );
  NOR2_X1 U423 ( .A1(n23), .A2(n39), .ZN(ab_20__15_) );
  NOR2_X1 U424 ( .A1(n24), .A2(n39), .ZN(ab_20__14_) );
  NOR2_X1 U425 ( .A1(n25), .A2(n39), .ZN(ab_20__13_) );
  NOR2_X1 U426 ( .A1(n26), .A2(n39), .ZN(ab_20__12_) );
  NOR2_X1 U427 ( .A1(n27), .A2(n39), .ZN(ab_20__11_) );
  NOR2_X1 U428 ( .A1(n28), .A2(n39), .ZN(ab_20__10_) );
  NOR2_X1 U429 ( .A1(n29), .A2(n39), .ZN(ab_20__0_) );
  NOR2_X1 U430 ( .A1(n7), .A2(n40), .ZN(ab_1__9_) );
  NOR2_X1 U431 ( .A1(n8), .A2(n40), .ZN(ab_1__8_) );
  NOR2_X1 U432 ( .A1(n9), .A2(n40), .ZN(ab_1__7_) );
  NOR2_X1 U433 ( .A1(n10), .A2(n40), .ZN(ab_1__6_) );
  NOR2_X1 U434 ( .A1(n11), .A2(n40), .ZN(ab_1__5_) );
  NOR2_X1 U435 ( .A1(n12), .A2(n40), .ZN(ab_1__4_) );
  NOR2_X1 U436 ( .A1(n13), .A2(n40), .ZN(ab_1__3_) );
  NOR2_X1 U437 ( .A1(n14), .A2(n40), .ZN(ab_1__2_) );
  NOR2_X1 U438 ( .A1(A[1]), .A2(n1), .ZN(ab_1__23_) );
  NOR2_X1 U439 ( .A1(n15), .A2(n40), .ZN(ab_1__22_) );
  NOR2_X1 U440 ( .A1(n16), .A2(n40), .ZN(ab_1__21_) );
  NOR2_X1 U441 ( .A1(n17), .A2(n40), .ZN(ab_1__20_) );
  NOR2_X1 U442 ( .A1(n19), .A2(n40), .ZN(ab_1__19_) );
  NOR2_X1 U443 ( .A1(n20), .A2(n40), .ZN(ab_1__18_) );
  NOR2_X1 U444 ( .A1(n21), .A2(n40), .ZN(ab_1__17_) );
  NOR2_X1 U445 ( .A1(n22), .A2(n40), .ZN(ab_1__16_) );
  NOR2_X1 U446 ( .A1(n23), .A2(n40), .ZN(ab_1__15_) );
  NOR2_X1 U447 ( .A1(n24), .A2(n40), .ZN(ab_1__14_) );
  NOR2_X1 U448 ( .A1(n25), .A2(n40), .ZN(ab_1__13_) );
  NOR2_X1 U449 ( .A1(n26), .A2(n40), .ZN(ab_1__12_) );
  NOR2_X1 U450 ( .A1(n27), .A2(n40), .ZN(ab_1__11_) );
  NOR2_X1 U451 ( .A1(n28), .A2(n40), .ZN(ab_1__10_) );
  NOR2_X1 U452 ( .A1(n7), .A2(n41), .ZN(ab_19__9_) );
  NOR2_X1 U453 ( .A1(n8), .A2(n41), .ZN(ab_19__8_) );
  NOR2_X1 U454 ( .A1(n9), .A2(n41), .ZN(ab_19__7_) );
  NOR2_X1 U455 ( .A1(n10), .A2(n41), .ZN(ab_19__6_) );
  NOR2_X1 U456 ( .A1(n11), .A2(n41), .ZN(ab_19__5_) );
  NOR2_X1 U457 ( .A1(n12), .A2(n41), .ZN(ab_19__4_) );
  NOR2_X1 U458 ( .A1(n13), .A2(n41), .ZN(ab_19__3_) );
  NOR2_X1 U459 ( .A1(n14), .A2(n41), .ZN(ab_19__2_) );
  NOR2_X1 U460 ( .A1(A[19]), .A2(n1), .ZN(ab_19__23_) );
  NOR2_X1 U461 ( .A1(n15), .A2(n41), .ZN(ab_19__22_) );
  NOR2_X1 U462 ( .A1(n16), .A2(n41), .ZN(ab_19__21_) );
  NOR2_X1 U463 ( .A1(n17), .A2(n41), .ZN(ab_19__20_) );
  NOR2_X1 U464 ( .A1(n18), .A2(n41), .ZN(ab_19__1_) );
  NOR2_X1 U465 ( .A1(n19), .A2(n41), .ZN(ab_19__19_) );
  NOR2_X1 U466 ( .A1(n20), .A2(n41), .ZN(ab_19__18_) );
  NOR2_X1 U467 ( .A1(n21), .A2(n41), .ZN(ab_19__17_) );
  NOR2_X1 U468 ( .A1(n22), .A2(n41), .ZN(ab_19__16_) );
  NOR2_X1 U469 ( .A1(n23), .A2(n41), .ZN(ab_19__15_) );
  NOR2_X1 U470 ( .A1(n24), .A2(n41), .ZN(ab_19__14_) );
  NOR2_X1 U471 ( .A1(n25), .A2(n41), .ZN(ab_19__13_) );
  NOR2_X1 U472 ( .A1(n26), .A2(n41), .ZN(ab_19__12_) );
  NOR2_X1 U473 ( .A1(n27), .A2(n41), .ZN(ab_19__11_) );
  NOR2_X1 U474 ( .A1(n28), .A2(n41), .ZN(ab_19__10_) );
  NOR2_X1 U475 ( .A1(n29), .A2(n41), .ZN(ab_19__0_) );
  NOR2_X1 U476 ( .A1(n7), .A2(n42), .ZN(ab_18__9_) );
  NOR2_X1 U477 ( .A1(n8), .A2(n42), .ZN(ab_18__8_) );
  NOR2_X1 U478 ( .A1(n9), .A2(n42), .ZN(ab_18__7_) );
  NOR2_X1 U479 ( .A1(n10), .A2(n42), .ZN(ab_18__6_) );
  NOR2_X1 U480 ( .A1(n11), .A2(n42), .ZN(ab_18__5_) );
  NOR2_X1 U481 ( .A1(n12), .A2(n42), .ZN(ab_18__4_) );
  NOR2_X1 U482 ( .A1(n13), .A2(n42), .ZN(ab_18__3_) );
  NOR2_X1 U483 ( .A1(n14), .A2(n42), .ZN(ab_18__2_) );
  NOR2_X1 U484 ( .A1(A[18]), .A2(n1), .ZN(ab_18__23_) );
  NOR2_X1 U485 ( .A1(n15), .A2(n42), .ZN(ab_18__22_) );
  NOR2_X1 U486 ( .A1(n16), .A2(n42), .ZN(ab_18__21_) );
  NOR2_X1 U487 ( .A1(n17), .A2(n42), .ZN(ab_18__20_) );
  NOR2_X1 U488 ( .A1(n18), .A2(n42), .ZN(ab_18__1_) );
  NOR2_X1 U489 ( .A1(n19), .A2(n42), .ZN(ab_18__19_) );
  NOR2_X1 U490 ( .A1(n20), .A2(n42), .ZN(ab_18__18_) );
  NOR2_X1 U491 ( .A1(n21), .A2(n42), .ZN(ab_18__17_) );
  NOR2_X1 U492 ( .A1(n22), .A2(n42), .ZN(ab_18__16_) );
  NOR2_X1 U493 ( .A1(n23), .A2(n42), .ZN(ab_18__15_) );
  NOR2_X1 U494 ( .A1(n24), .A2(n42), .ZN(ab_18__14_) );
  NOR2_X1 U495 ( .A1(n25), .A2(n42), .ZN(ab_18__13_) );
  NOR2_X1 U496 ( .A1(n26), .A2(n42), .ZN(ab_18__12_) );
  NOR2_X1 U497 ( .A1(n27), .A2(n42), .ZN(ab_18__11_) );
  NOR2_X1 U498 ( .A1(n28), .A2(n42), .ZN(ab_18__10_) );
  NOR2_X1 U499 ( .A1(n29), .A2(n42), .ZN(ab_18__0_) );
  NOR2_X1 U500 ( .A1(n7), .A2(n43), .ZN(ab_17__9_) );
  NOR2_X1 U501 ( .A1(n8), .A2(n43), .ZN(ab_17__8_) );
  NOR2_X1 U502 ( .A1(n9), .A2(n43), .ZN(ab_17__7_) );
  NOR2_X1 U503 ( .A1(n10), .A2(n43), .ZN(ab_17__6_) );
  NOR2_X1 U504 ( .A1(n11), .A2(n43), .ZN(ab_17__5_) );
  NOR2_X1 U505 ( .A1(n12), .A2(n43), .ZN(ab_17__4_) );
  NOR2_X1 U506 ( .A1(n13), .A2(n43), .ZN(ab_17__3_) );
  NOR2_X1 U507 ( .A1(n14), .A2(n43), .ZN(ab_17__2_) );
  NOR2_X1 U508 ( .A1(A[17]), .A2(n1), .ZN(ab_17__23_) );
  NOR2_X1 U509 ( .A1(n15), .A2(n43), .ZN(ab_17__22_) );
  NOR2_X1 U510 ( .A1(n16), .A2(n43), .ZN(ab_17__21_) );
  NOR2_X1 U511 ( .A1(n17), .A2(n43), .ZN(ab_17__20_) );
  NOR2_X1 U512 ( .A1(n18), .A2(n43), .ZN(ab_17__1_) );
  NOR2_X1 U513 ( .A1(n19), .A2(n43), .ZN(ab_17__19_) );
  NOR2_X1 U514 ( .A1(n20), .A2(n43), .ZN(ab_17__18_) );
  NOR2_X1 U515 ( .A1(n21), .A2(n43), .ZN(ab_17__17_) );
  NOR2_X1 U516 ( .A1(n22), .A2(n43), .ZN(ab_17__16_) );
  NOR2_X1 U517 ( .A1(n23), .A2(n43), .ZN(ab_17__15_) );
  NOR2_X1 U518 ( .A1(n24), .A2(n43), .ZN(ab_17__14_) );
  NOR2_X1 U519 ( .A1(n25), .A2(n43), .ZN(ab_17__13_) );
  NOR2_X1 U520 ( .A1(n26), .A2(n43), .ZN(ab_17__12_) );
  NOR2_X1 U521 ( .A1(n27), .A2(n43), .ZN(ab_17__11_) );
  NOR2_X1 U522 ( .A1(n28), .A2(n43), .ZN(ab_17__10_) );
  NOR2_X1 U523 ( .A1(n29), .A2(n43), .ZN(ab_17__0_) );
  NOR2_X1 U524 ( .A1(n7), .A2(n44), .ZN(ab_16__9_) );
  NOR2_X1 U525 ( .A1(n8), .A2(n44), .ZN(ab_16__8_) );
  NOR2_X1 U526 ( .A1(n9), .A2(n44), .ZN(ab_16__7_) );
  NOR2_X1 U527 ( .A1(n10), .A2(n44), .ZN(ab_16__6_) );
  NOR2_X1 U528 ( .A1(n11), .A2(n44), .ZN(ab_16__5_) );
  NOR2_X1 U529 ( .A1(n12), .A2(n44), .ZN(ab_16__4_) );
  NOR2_X1 U530 ( .A1(n13), .A2(n44), .ZN(ab_16__3_) );
  NOR2_X1 U531 ( .A1(n14), .A2(n44), .ZN(ab_16__2_) );
  NOR2_X1 U532 ( .A1(A[16]), .A2(n1), .ZN(ab_16__23_) );
  NOR2_X1 U533 ( .A1(n15), .A2(n44), .ZN(ab_16__22_) );
  NOR2_X1 U534 ( .A1(n16), .A2(n44), .ZN(ab_16__21_) );
  NOR2_X1 U535 ( .A1(n17), .A2(n44), .ZN(ab_16__20_) );
  NOR2_X1 U536 ( .A1(n18), .A2(n44), .ZN(ab_16__1_) );
  NOR2_X1 U537 ( .A1(n19), .A2(n44), .ZN(ab_16__19_) );
  NOR2_X1 U538 ( .A1(n20), .A2(n44), .ZN(ab_16__18_) );
  NOR2_X1 U539 ( .A1(n21), .A2(n44), .ZN(ab_16__17_) );
  NOR2_X1 U540 ( .A1(n22), .A2(n44), .ZN(ab_16__16_) );
  NOR2_X1 U541 ( .A1(n23), .A2(n44), .ZN(ab_16__15_) );
  NOR2_X1 U542 ( .A1(n24), .A2(n44), .ZN(ab_16__14_) );
  NOR2_X1 U543 ( .A1(n25), .A2(n44), .ZN(ab_16__13_) );
  NOR2_X1 U544 ( .A1(n26), .A2(n44), .ZN(ab_16__12_) );
  NOR2_X1 U545 ( .A1(n27), .A2(n44), .ZN(ab_16__11_) );
  NOR2_X1 U546 ( .A1(n28), .A2(n44), .ZN(ab_16__10_) );
  NOR2_X1 U547 ( .A1(n29), .A2(n44), .ZN(ab_16__0_) );
  NOR2_X1 U548 ( .A1(n7), .A2(n45), .ZN(ab_15__9_) );
  NOR2_X1 U549 ( .A1(n8), .A2(n45), .ZN(ab_15__8_) );
  NOR2_X1 U550 ( .A1(n9), .A2(n45), .ZN(ab_15__7_) );
  NOR2_X1 U551 ( .A1(n10), .A2(n45), .ZN(ab_15__6_) );
  NOR2_X1 U552 ( .A1(n11), .A2(n45), .ZN(ab_15__5_) );
  NOR2_X1 U553 ( .A1(n12), .A2(n45), .ZN(ab_15__4_) );
  NOR2_X1 U554 ( .A1(n13), .A2(n45), .ZN(ab_15__3_) );
  NOR2_X1 U555 ( .A1(n14), .A2(n45), .ZN(ab_15__2_) );
  NOR2_X1 U556 ( .A1(A[15]), .A2(n1), .ZN(ab_15__23_) );
  NOR2_X1 U557 ( .A1(n15), .A2(n45), .ZN(ab_15__22_) );
  NOR2_X1 U558 ( .A1(n16), .A2(n45), .ZN(ab_15__21_) );
  NOR2_X1 U559 ( .A1(n17), .A2(n45), .ZN(ab_15__20_) );
  NOR2_X1 U560 ( .A1(n18), .A2(n45), .ZN(ab_15__1_) );
  NOR2_X1 U561 ( .A1(n19), .A2(n45), .ZN(ab_15__19_) );
  NOR2_X1 U562 ( .A1(n20), .A2(n45), .ZN(ab_15__18_) );
  NOR2_X1 U563 ( .A1(n21), .A2(n45), .ZN(ab_15__17_) );
  NOR2_X1 U564 ( .A1(n22), .A2(n45), .ZN(ab_15__16_) );
  NOR2_X1 U565 ( .A1(n23), .A2(n45), .ZN(ab_15__15_) );
  NOR2_X1 U566 ( .A1(n24), .A2(n45), .ZN(ab_15__14_) );
  NOR2_X1 U567 ( .A1(n25), .A2(n45), .ZN(ab_15__13_) );
  NOR2_X1 U568 ( .A1(n26), .A2(n45), .ZN(ab_15__12_) );
  NOR2_X1 U569 ( .A1(n27), .A2(n45), .ZN(ab_15__11_) );
  NOR2_X1 U570 ( .A1(n28), .A2(n45), .ZN(ab_15__10_) );
  NOR2_X1 U571 ( .A1(n29), .A2(n45), .ZN(ab_15__0_) );
  NOR2_X1 U572 ( .A1(n7), .A2(n46), .ZN(ab_14__9_) );
  NOR2_X1 U573 ( .A1(n8), .A2(n46), .ZN(ab_14__8_) );
  NOR2_X1 U574 ( .A1(n9), .A2(n46), .ZN(ab_14__7_) );
  NOR2_X1 U575 ( .A1(n10), .A2(n46), .ZN(ab_14__6_) );
  NOR2_X1 U576 ( .A1(n11), .A2(n46), .ZN(ab_14__5_) );
  NOR2_X1 U577 ( .A1(n12), .A2(n46), .ZN(ab_14__4_) );
  NOR2_X1 U578 ( .A1(n13), .A2(n46), .ZN(ab_14__3_) );
  NOR2_X1 U579 ( .A1(n14), .A2(n46), .ZN(ab_14__2_) );
  NOR2_X1 U580 ( .A1(A[14]), .A2(n2), .ZN(ab_14__23_) );
  NOR2_X1 U581 ( .A1(n15), .A2(n46), .ZN(ab_14__22_) );
  NOR2_X1 U582 ( .A1(n16), .A2(n46), .ZN(ab_14__21_) );
  NOR2_X1 U583 ( .A1(n17), .A2(n46), .ZN(ab_14__20_) );
  NOR2_X1 U584 ( .A1(n18), .A2(n46), .ZN(ab_14__1_) );
  NOR2_X1 U585 ( .A1(n19), .A2(n46), .ZN(ab_14__19_) );
  NOR2_X1 U586 ( .A1(n20), .A2(n46), .ZN(ab_14__18_) );
  NOR2_X1 U587 ( .A1(n21), .A2(n46), .ZN(ab_14__17_) );
  NOR2_X1 U588 ( .A1(n22), .A2(n46), .ZN(ab_14__16_) );
  NOR2_X1 U589 ( .A1(n23), .A2(n46), .ZN(ab_14__15_) );
  NOR2_X1 U590 ( .A1(n24), .A2(n46), .ZN(ab_14__14_) );
  NOR2_X1 U591 ( .A1(n25), .A2(n46), .ZN(ab_14__13_) );
  NOR2_X1 U592 ( .A1(n26), .A2(n46), .ZN(ab_14__12_) );
  NOR2_X1 U593 ( .A1(n27), .A2(n46), .ZN(ab_14__11_) );
  NOR2_X1 U594 ( .A1(n28), .A2(n46), .ZN(ab_14__10_) );
  NOR2_X1 U595 ( .A1(n29), .A2(n46), .ZN(ab_14__0_) );
  NOR2_X1 U596 ( .A1(n7), .A2(n47), .ZN(ab_13__9_) );
  NOR2_X1 U597 ( .A1(n8), .A2(n47), .ZN(ab_13__8_) );
  NOR2_X1 U598 ( .A1(n9), .A2(n47), .ZN(ab_13__7_) );
  NOR2_X1 U599 ( .A1(n10), .A2(n47), .ZN(ab_13__6_) );
  NOR2_X1 U600 ( .A1(n11), .A2(n47), .ZN(ab_13__5_) );
  NOR2_X1 U601 ( .A1(n12), .A2(n47), .ZN(ab_13__4_) );
  NOR2_X1 U602 ( .A1(n13), .A2(n47), .ZN(ab_13__3_) );
  NOR2_X1 U603 ( .A1(n14), .A2(n47), .ZN(ab_13__2_) );
  NOR2_X1 U604 ( .A1(A[13]), .A2(n2), .ZN(ab_13__23_) );
  NOR2_X1 U605 ( .A1(n15), .A2(n47), .ZN(ab_13__22_) );
  NOR2_X1 U606 ( .A1(n16), .A2(n47), .ZN(ab_13__21_) );
  NOR2_X1 U607 ( .A1(n17), .A2(n47), .ZN(ab_13__20_) );
  NOR2_X1 U608 ( .A1(n18), .A2(n47), .ZN(ab_13__1_) );
  NOR2_X1 U609 ( .A1(n19), .A2(n47), .ZN(ab_13__19_) );
  NOR2_X1 U610 ( .A1(n20), .A2(n47), .ZN(ab_13__18_) );
  NOR2_X1 U611 ( .A1(n21), .A2(n47), .ZN(ab_13__17_) );
  NOR2_X1 U612 ( .A1(n22), .A2(n47), .ZN(ab_13__16_) );
  NOR2_X1 U613 ( .A1(n23), .A2(n47), .ZN(ab_13__15_) );
  NOR2_X1 U614 ( .A1(n24), .A2(n47), .ZN(ab_13__14_) );
  NOR2_X1 U615 ( .A1(n25), .A2(n47), .ZN(ab_13__13_) );
  NOR2_X1 U616 ( .A1(n26), .A2(n47), .ZN(ab_13__12_) );
  NOR2_X1 U617 ( .A1(n27), .A2(n47), .ZN(ab_13__11_) );
  NOR2_X1 U618 ( .A1(n28), .A2(n47), .ZN(ab_13__10_) );
  NOR2_X1 U619 ( .A1(n29), .A2(n47), .ZN(ab_13__0_) );
  NOR2_X1 U620 ( .A1(n7), .A2(n48), .ZN(ab_12__9_) );
  NOR2_X1 U621 ( .A1(n8), .A2(n48), .ZN(ab_12__8_) );
  NOR2_X1 U622 ( .A1(n9), .A2(n48), .ZN(ab_12__7_) );
  NOR2_X1 U623 ( .A1(n10), .A2(n48), .ZN(ab_12__6_) );
  NOR2_X1 U624 ( .A1(n11), .A2(n48), .ZN(ab_12__5_) );
  NOR2_X1 U625 ( .A1(n12), .A2(n48), .ZN(ab_12__4_) );
  NOR2_X1 U626 ( .A1(n13), .A2(n48), .ZN(ab_12__3_) );
  NOR2_X1 U627 ( .A1(n14), .A2(n48), .ZN(ab_12__2_) );
  NOR2_X1 U628 ( .A1(A[12]), .A2(n2), .ZN(ab_12__23_) );
  NOR2_X1 U629 ( .A1(n15), .A2(n48), .ZN(ab_12__22_) );
  NOR2_X1 U630 ( .A1(n16), .A2(n48), .ZN(ab_12__21_) );
  NOR2_X1 U631 ( .A1(n17), .A2(n48), .ZN(ab_12__20_) );
  NOR2_X1 U632 ( .A1(n18), .A2(n48), .ZN(ab_12__1_) );
  NOR2_X1 U633 ( .A1(n19), .A2(n48), .ZN(ab_12__19_) );
  NOR2_X1 U634 ( .A1(n20), .A2(n48), .ZN(ab_12__18_) );
  NOR2_X1 U635 ( .A1(n21), .A2(n48), .ZN(ab_12__17_) );
  NOR2_X1 U636 ( .A1(n22), .A2(n48), .ZN(ab_12__16_) );
  NOR2_X1 U637 ( .A1(n23), .A2(n48), .ZN(ab_12__15_) );
  NOR2_X1 U638 ( .A1(n24), .A2(n48), .ZN(ab_12__14_) );
  NOR2_X1 U639 ( .A1(n25), .A2(n48), .ZN(ab_12__13_) );
  NOR2_X1 U640 ( .A1(n26), .A2(n48), .ZN(ab_12__12_) );
  NOR2_X1 U641 ( .A1(n27), .A2(n48), .ZN(ab_12__11_) );
  NOR2_X1 U642 ( .A1(n28), .A2(n48), .ZN(ab_12__10_) );
  NOR2_X1 U643 ( .A1(n29), .A2(n48), .ZN(ab_12__0_) );
  NOR2_X1 U644 ( .A1(n7), .A2(n49), .ZN(ab_11__9_) );
  NOR2_X1 U645 ( .A1(n8), .A2(n49), .ZN(ab_11__8_) );
  NOR2_X1 U646 ( .A1(n9), .A2(n49), .ZN(ab_11__7_) );
  NOR2_X1 U647 ( .A1(n10), .A2(n49), .ZN(ab_11__6_) );
  NOR2_X1 U648 ( .A1(n11), .A2(n49), .ZN(ab_11__5_) );
  NOR2_X1 U649 ( .A1(n12), .A2(n49), .ZN(ab_11__4_) );
  NOR2_X1 U650 ( .A1(n13), .A2(n49), .ZN(ab_11__3_) );
  NOR2_X1 U651 ( .A1(n14), .A2(n49), .ZN(ab_11__2_) );
  NOR2_X1 U652 ( .A1(A[11]), .A2(n2), .ZN(ab_11__23_) );
  NOR2_X1 U653 ( .A1(n15), .A2(n49), .ZN(ab_11__22_) );
  NOR2_X1 U654 ( .A1(n16), .A2(n49), .ZN(ab_11__21_) );
  NOR2_X1 U655 ( .A1(n17), .A2(n49), .ZN(ab_11__20_) );
  NOR2_X1 U656 ( .A1(n18), .A2(n49), .ZN(ab_11__1_) );
  NOR2_X1 U657 ( .A1(n19), .A2(n49), .ZN(ab_11__19_) );
  NOR2_X1 U658 ( .A1(n20), .A2(n49), .ZN(ab_11__18_) );
  NOR2_X1 U659 ( .A1(n21), .A2(n49), .ZN(ab_11__17_) );
  NOR2_X1 U660 ( .A1(n22), .A2(n49), .ZN(ab_11__16_) );
  NOR2_X1 U661 ( .A1(n23), .A2(n49), .ZN(ab_11__15_) );
  NOR2_X1 U662 ( .A1(n24), .A2(n49), .ZN(ab_11__14_) );
  NOR2_X1 U663 ( .A1(n25), .A2(n49), .ZN(ab_11__13_) );
  NOR2_X1 U664 ( .A1(n26), .A2(n49), .ZN(ab_11__12_) );
  NOR2_X1 U665 ( .A1(n27), .A2(n49), .ZN(ab_11__11_) );
  NOR2_X1 U666 ( .A1(n28), .A2(n49), .ZN(ab_11__10_) );
  NOR2_X1 U667 ( .A1(n29), .A2(n49), .ZN(ab_11__0_) );
  NOR2_X1 U668 ( .A1(n7), .A2(n50), .ZN(ab_10__9_) );
  NOR2_X1 U669 ( .A1(n8), .A2(n50), .ZN(ab_10__8_) );
  NOR2_X1 U670 ( .A1(n9), .A2(n50), .ZN(ab_10__7_) );
  NOR2_X1 U671 ( .A1(n10), .A2(n50), .ZN(ab_10__6_) );
  NOR2_X1 U672 ( .A1(n11), .A2(n50), .ZN(ab_10__5_) );
  NOR2_X1 U673 ( .A1(n12), .A2(n50), .ZN(ab_10__4_) );
  NOR2_X1 U674 ( .A1(n13), .A2(n50), .ZN(ab_10__3_) );
  NOR2_X1 U675 ( .A1(n14), .A2(n50), .ZN(ab_10__2_) );
  NOR2_X1 U676 ( .A1(A[10]), .A2(n2), .ZN(ab_10__23_) );
  NOR2_X1 U677 ( .A1(n15), .A2(n50), .ZN(ab_10__22_) );
  NOR2_X1 U678 ( .A1(n16), .A2(n50), .ZN(ab_10__21_) );
  NOR2_X1 U679 ( .A1(n17), .A2(n50), .ZN(ab_10__20_) );
  NOR2_X1 U680 ( .A1(n18), .A2(n50), .ZN(ab_10__1_) );
  NOR2_X1 U681 ( .A1(n19), .A2(n50), .ZN(ab_10__19_) );
  NOR2_X1 U682 ( .A1(n20), .A2(n50), .ZN(ab_10__18_) );
  NOR2_X1 U683 ( .A1(n21), .A2(n50), .ZN(ab_10__17_) );
  NOR2_X1 U684 ( .A1(n22), .A2(n50), .ZN(ab_10__16_) );
  NOR2_X1 U685 ( .A1(n23), .A2(n50), .ZN(ab_10__15_) );
  NOR2_X1 U686 ( .A1(n24), .A2(n50), .ZN(ab_10__14_) );
  NOR2_X1 U687 ( .A1(n25), .A2(n50), .ZN(ab_10__13_) );
  NOR2_X1 U688 ( .A1(n26), .A2(n50), .ZN(ab_10__12_) );
  NOR2_X1 U689 ( .A1(n27), .A2(n50), .ZN(ab_10__11_) );
  NOR2_X1 U690 ( .A1(n28), .A2(n50), .ZN(ab_10__10_) );
  NOR2_X1 U691 ( .A1(n29), .A2(n50), .ZN(ab_10__0_) );
  NOR2_X1 U692 ( .A1(n7), .A2(n51), .ZN(ab_0__9_) );
  NOR2_X1 U693 ( .A1(n8), .A2(n51), .ZN(ab_0__8_) );
  NOR2_X1 U694 ( .A1(n9), .A2(n51), .ZN(ab_0__7_) );
  NOR2_X1 U695 ( .A1(n10), .A2(n51), .ZN(ab_0__6_) );
  NOR2_X1 U696 ( .A1(n11), .A2(n51), .ZN(ab_0__5_) );
  NOR2_X1 U697 ( .A1(n12), .A2(n51), .ZN(ab_0__4_) );
  NOR2_X1 U698 ( .A1(n13), .A2(n51), .ZN(ab_0__3_) );
  NOR2_X1 U699 ( .A1(n14), .A2(n51), .ZN(ab_0__2_) );
  NOR2_X1 U700 ( .A1(A[0]), .A2(n1), .ZN(ab_0__23_) );
  NOR2_X1 U701 ( .A1(n15), .A2(n51), .ZN(ab_0__22_) );
  NOR2_X1 U702 ( .A1(n16), .A2(n51), .ZN(ab_0__21_) );
  NOR2_X1 U703 ( .A1(n17), .A2(n51), .ZN(ab_0__20_) );
  NOR2_X1 U704 ( .A1(n19), .A2(n51), .ZN(ab_0__19_) );
  NOR2_X1 U705 ( .A1(n20), .A2(n51), .ZN(ab_0__18_) );
  NOR2_X1 U706 ( .A1(n21), .A2(n51), .ZN(ab_0__17_) );
  NOR2_X1 U707 ( .A1(n22), .A2(n51), .ZN(ab_0__16_) );
  NOR2_X1 U708 ( .A1(n23), .A2(n51), .ZN(ab_0__15_) );
  NOR2_X1 U709 ( .A1(n24), .A2(n51), .ZN(ab_0__14_) );
  NOR2_X1 U710 ( .A1(n25), .A2(n51), .ZN(ab_0__13_) );
  NOR2_X1 U711 ( .A1(n26), .A2(n51), .ZN(ab_0__12_) );
  NOR2_X1 U712 ( .A1(n27), .A2(n51), .ZN(ab_0__11_) );
  NOR2_X1 U713 ( .A1(n28), .A2(n51), .ZN(ab_0__10_) );
  INV_X1 U714 ( .A(B[23]), .ZN(QB) );
  INV_X1 U715 ( .A(A[23]), .ZN(QA) );
  AND3_X1 U716 ( .A1(ab_1__1_), .A2(B[0]), .A3(A[0]), .ZN(CARRYB_1__0_) );
  NOR2_X1 U717 ( .A1(n40), .A2(n18), .ZN(ab_1__1_) );
  INV_X1 U719 ( .A(CARRYB_23__23_), .ZN(A1_45_) );
endmodule


module iir_filter_DW01_add_4 ( A, B, CI, SUM, CO );
  input [45:0] A;
  input [45:0] B;
  output [45:0] SUM;
  input CI;
  output CO;
  wire   A_21_, A_20_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112;
  assign SUM[21] = A_21_;
  assign A_21_ = A[21];
  assign SUM[20] = A_20_;
  assign A_20_ = A[20];

  XOR2_X1 U2 ( .A(n1), .B(n2), .Z(SUM[45]) );
  XOR2_X1 U3 ( .A(B[45]), .B(A[45]), .Z(n2) );
  OAI21_X1 U4 ( .B1(n3), .B2(n4), .A(n5), .ZN(n1) );
  OAI21_X1 U5 ( .B1(A[44]), .B2(n6), .A(B[44]), .ZN(n5) );
  INV_X1 U6 ( .A(n3), .ZN(n6) );
  INV_X1 U7 ( .A(A[44]), .ZN(n4) );
  AOI21_X1 U8 ( .B1(A[43]), .B2(B[43]), .A(n7), .ZN(n3) );
  INV_X1 U9 ( .A(n8), .ZN(n7) );
  OAI22_X1 U10 ( .A1(n9), .A2(n10), .B1(A[43]), .B2(B[43]), .ZN(n8) );
  AOI21_X1 U11 ( .B1(n11), .B2(n12), .A(n13), .ZN(n9) );
  NAND3_X1 U12 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n12) );
  AOI21_X1 U13 ( .B1(n17), .B2(n16), .A(n18), .ZN(n11) );
  INV_X1 U14 ( .A(n19), .ZN(n18) );
  XOR2_X1 U15 ( .A(n20), .B(n21), .Z(SUM[42]) );
  NOR2_X1 U16 ( .A1(n10), .A2(n13), .ZN(n21) );
  NOR2_X1 U17 ( .A1(B[42]), .A2(A[42]), .ZN(n13) );
  AND2_X1 U18 ( .A1(B[42]), .A2(A[42]), .ZN(n10) );
  OAI21_X1 U19 ( .B1(n22), .B2(n23), .A(n19), .ZN(n20) );
  XOR2_X1 U20 ( .A(n24), .B(n23), .Z(SUM[41]) );
  AOI21_X1 U21 ( .B1(n15), .B2(n14), .A(n17), .ZN(n23) );
  INV_X1 U22 ( .A(n25), .ZN(n15) );
  NAND2_X1 U23 ( .A1(n16), .A2(n19), .ZN(n24) );
  NAND2_X1 U24 ( .A1(B[41]), .A2(A[41]), .ZN(n19) );
  INV_X1 U25 ( .A(n22), .ZN(n16) );
  NOR2_X1 U26 ( .A1(B[41]), .A2(A[41]), .ZN(n22) );
  XOR2_X1 U27 ( .A(n14), .B(n26), .Z(SUM[40]) );
  NOR2_X1 U28 ( .A1(n17), .A2(n25), .ZN(n26) );
  NOR2_X1 U29 ( .A1(B[40]), .A2(A[40]), .ZN(n25) );
  AND2_X1 U30 ( .A1(B[40]), .A2(A[40]), .ZN(n17) );
  OAI21_X1 U31 ( .B1(n27), .B2(n28), .A(n29), .ZN(n14) );
  XOR2_X1 U32 ( .A(n30), .B(n28), .Z(SUM[39]) );
  AOI21_X1 U33 ( .B1(n31), .B2(n32), .A(n33), .ZN(n28) );
  INV_X1 U34 ( .A(n34), .ZN(n31) );
  NAND2_X1 U35 ( .A1(n35), .A2(n29), .ZN(n30) );
  NAND2_X1 U36 ( .A1(B[39]), .A2(A[39]), .ZN(n29) );
  INV_X1 U37 ( .A(n27), .ZN(n35) );
  NOR2_X1 U38 ( .A1(B[39]), .A2(A[39]), .ZN(n27) );
  XOR2_X1 U39 ( .A(n32), .B(n36), .Z(SUM[38]) );
  NOR2_X1 U40 ( .A1(n33), .A2(n34), .ZN(n36) );
  NOR2_X1 U41 ( .A1(B[38]), .A2(A[38]), .ZN(n34) );
  AND2_X1 U42 ( .A1(B[38]), .A2(A[38]), .ZN(n33) );
  OAI21_X1 U43 ( .B1(n37), .B2(n38), .A(n39), .ZN(n32) );
  XOR2_X1 U44 ( .A(n40), .B(n38), .Z(SUM[37]) );
  AOI21_X1 U45 ( .B1(n41), .B2(n42), .A(n43), .ZN(n38) );
  INV_X1 U46 ( .A(n44), .ZN(n41) );
  NAND2_X1 U47 ( .A1(n45), .A2(n39), .ZN(n40) );
  NAND2_X1 U48 ( .A1(B[37]), .A2(A[37]), .ZN(n39) );
  INV_X1 U49 ( .A(n37), .ZN(n45) );
  NOR2_X1 U50 ( .A1(B[37]), .A2(A[37]), .ZN(n37) );
  XOR2_X1 U51 ( .A(n42), .B(n46), .Z(SUM[36]) );
  NOR2_X1 U52 ( .A1(n43), .A2(n44), .ZN(n46) );
  NOR2_X1 U53 ( .A1(B[36]), .A2(A[36]), .ZN(n44) );
  AND2_X1 U54 ( .A1(B[36]), .A2(A[36]), .ZN(n43) );
  OAI21_X1 U55 ( .B1(n47), .B2(n48), .A(n49), .ZN(n42) );
  XOR2_X1 U56 ( .A(n50), .B(n48), .Z(SUM[35]) );
  AOI21_X1 U57 ( .B1(n51), .B2(n52), .A(n53), .ZN(n48) );
  INV_X1 U58 ( .A(n54), .ZN(n51) );
  NAND2_X1 U59 ( .A1(n55), .A2(n49), .ZN(n50) );
  NAND2_X1 U60 ( .A1(B[35]), .A2(A[35]), .ZN(n49) );
  INV_X1 U61 ( .A(n47), .ZN(n55) );
  NOR2_X1 U62 ( .A1(B[35]), .A2(A[35]), .ZN(n47) );
  XOR2_X1 U63 ( .A(n52), .B(n56), .Z(SUM[34]) );
  NOR2_X1 U64 ( .A1(n53), .A2(n54), .ZN(n56) );
  NOR2_X1 U65 ( .A1(B[34]), .A2(A[34]), .ZN(n54) );
  AND2_X1 U66 ( .A1(B[34]), .A2(A[34]), .ZN(n53) );
  OAI21_X1 U67 ( .B1(n57), .B2(n58), .A(n59), .ZN(n52) );
  XOR2_X1 U68 ( .A(n60), .B(n58), .Z(SUM[33]) );
  AOI21_X1 U69 ( .B1(n61), .B2(n62), .A(n63), .ZN(n58) );
  INV_X1 U70 ( .A(n64), .ZN(n61) );
  NAND2_X1 U71 ( .A1(n65), .A2(n59), .ZN(n60) );
  NAND2_X1 U72 ( .A1(B[33]), .A2(A[33]), .ZN(n59) );
  INV_X1 U73 ( .A(n57), .ZN(n65) );
  NOR2_X1 U74 ( .A1(B[33]), .A2(A[33]), .ZN(n57) );
  XOR2_X1 U75 ( .A(n62), .B(n66), .Z(SUM[32]) );
  NOR2_X1 U76 ( .A1(n63), .A2(n64), .ZN(n66) );
  NOR2_X1 U77 ( .A1(B[32]), .A2(A[32]), .ZN(n64) );
  AND2_X1 U78 ( .A1(B[32]), .A2(A[32]), .ZN(n63) );
  OAI21_X1 U79 ( .B1(n67), .B2(n68), .A(n69), .ZN(n62) );
  XOR2_X1 U80 ( .A(n70), .B(n68), .Z(SUM[31]) );
  AOI21_X1 U81 ( .B1(n71), .B2(n72), .A(n73), .ZN(n68) );
  INV_X1 U82 ( .A(n74), .ZN(n71) );
  NAND2_X1 U83 ( .A1(n75), .A2(n69), .ZN(n70) );
  NAND2_X1 U84 ( .A1(B[31]), .A2(A[31]), .ZN(n69) );
  INV_X1 U85 ( .A(n67), .ZN(n75) );
  NOR2_X1 U86 ( .A1(B[31]), .A2(A[31]), .ZN(n67) );
  XOR2_X1 U87 ( .A(n72), .B(n76), .Z(SUM[30]) );
  NOR2_X1 U88 ( .A1(n73), .A2(n74), .ZN(n76) );
  NOR2_X1 U89 ( .A1(B[30]), .A2(A[30]), .ZN(n74) );
  AND2_X1 U90 ( .A1(B[30]), .A2(A[30]), .ZN(n73) );
  OAI21_X1 U91 ( .B1(n77), .B2(n78), .A(n79), .ZN(n72) );
  XOR2_X1 U92 ( .A(n80), .B(n78), .Z(SUM[29]) );
  AOI21_X1 U93 ( .B1(n81), .B2(n82), .A(n83), .ZN(n78) );
  INV_X1 U94 ( .A(n84), .ZN(n81) );
  NAND2_X1 U95 ( .A1(n85), .A2(n79), .ZN(n80) );
  NAND2_X1 U96 ( .A1(B[29]), .A2(A[29]), .ZN(n79) );
  INV_X1 U97 ( .A(n77), .ZN(n85) );
  NOR2_X1 U98 ( .A1(B[29]), .A2(A[29]), .ZN(n77) );
  XOR2_X1 U99 ( .A(n82), .B(n86), .Z(SUM[28]) );
  NOR2_X1 U100 ( .A1(n83), .A2(n84), .ZN(n86) );
  NOR2_X1 U101 ( .A1(B[28]), .A2(A[28]), .ZN(n84) );
  AND2_X1 U102 ( .A1(B[28]), .A2(A[28]), .ZN(n83) );
  OAI21_X1 U103 ( .B1(n87), .B2(n88), .A(n89), .ZN(n82) );
  XOR2_X1 U104 ( .A(n90), .B(n88), .Z(SUM[27]) );
  AOI21_X1 U105 ( .B1(n91), .B2(n92), .A(n93), .ZN(n88) );
  INV_X1 U106 ( .A(n94), .ZN(n92) );
  NAND2_X1 U107 ( .A1(n95), .A2(n89), .ZN(n90) );
  NAND2_X1 U108 ( .A1(B[27]), .A2(A[27]), .ZN(n89) );
  INV_X1 U109 ( .A(n87), .ZN(n95) );
  NOR2_X1 U110 ( .A1(B[27]), .A2(A[27]), .ZN(n87) );
  XOR2_X1 U111 ( .A(n91), .B(n96), .Z(SUM[26]) );
  NOR2_X1 U112 ( .A1(n93), .A2(n94), .ZN(n96) );
  NOR2_X1 U113 ( .A1(B[26]), .A2(A[26]), .ZN(n94) );
  AND2_X1 U114 ( .A1(B[26]), .A2(A[26]), .ZN(n93) );
  OAI21_X1 U115 ( .B1(n97), .B2(n98), .A(n99), .ZN(n91) );
  XOR2_X1 U116 ( .A(n100), .B(n98), .Z(SUM[25]) );
  AOI21_X1 U117 ( .B1(n101), .B2(n102), .A(n103), .ZN(n98) );
  INV_X1 U118 ( .A(n104), .ZN(n101) );
  NAND2_X1 U119 ( .A1(n105), .A2(n99), .ZN(n100) );
  NAND2_X1 U120 ( .A1(B[25]), .A2(A[25]), .ZN(n99) );
  INV_X1 U121 ( .A(n97), .ZN(n105) );
  NOR2_X1 U122 ( .A1(B[25]), .A2(A[25]), .ZN(n97) );
  XOR2_X1 U123 ( .A(n102), .B(n106), .Z(SUM[24]) );
  NOR2_X1 U124 ( .A1(n103), .A2(n104), .ZN(n106) );
  NOR2_X1 U125 ( .A1(B[24]), .A2(A[24]), .ZN(n104) );
  AND2_X1 U126 ( .A1(B[24]), .A2(A[24]), .ZN(n103) );
  OAI21_X1 U127 ( .B1(n107), .B2(n108), .A(n109), .ZN(n102) );
  XOR2_X1 U128 ( .A(n108), .B(n110), .Z(SUM[23]) );
  NAND2_X1 U129 ( .A1(n111), .A2(n109), .ZN(n110) );
  NAND2_X1 U130 ( .A1(B[23]), .A2(A[23]), .ZN(n109) );
  INV_X1 U131 ( .A(n107), .ZN(n111) );
  NOR2_X1 U132 ( .A1(B[23]), .A2(A[23]), .ZN(n107) );
  INV_X1 U133 ( .A(n112), .ZN(SUM[22]) );
  OAI21_X1 U134 ( .B1(B[22]), .B2(A[22]), .A(n108), .ZN(n112) );
  NAND2_X1 U135 ( .A1(B[22]), .A2(A[22]), .ZN(n108) );
endmodule


module iir_filter_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [23:0] A;
  input [23:0] B;
  output [47:0] PRODUCT;
  input TC;
  wire   ab_23__23_, ab_23__22_, ab_23__21_, ab_23__20_, ab_23__19_,
         ab_23__18_, ab_23__17_, ab_23__16_, ab_23__15_, ab_23__14_,
         ab_23__13_, ab_23__12_, ab_23__11_, ab_23__10_, ab_23__9_, ab_23__8_,
         ab_23__7_, ab_23__6_, ab_23__5_, ab_23__4_, ab_23__3_, ab_23__2_,
         ab_23__1_, ab_23__0_, ab_22__23_, ab_22__22_, ab_22__21_, ab_22__20_,
         ab_22__19_, ab_22__18_, ab_22__17_, ab_22__16_, ab_22__15_,
         ab_22__14_, ab_22__13_, ab_22__12_, ab_22__11_, ab_22__10_, ab_22__9_,
         ab_22__8_, ab_22__7_, ab_22__6_, ab_22__5_, ab_22__4_, ab_22__3_,
         ab_22__2_, ab_22__1_, ab_22__0_, ab_21__23_, ab_21__22_, ab_21__21_,
         ab_21__20_, ab_21__19_, ab_21__18_, ab_21__17_, ab_21__16_,
         ab_21__15_, ab_21__14_, ab_21__13_, ab_21__12_, ab_21__11_,
         ab_21__10_, ab_21__9_, ab_21__8_, ab_21__7_, ab_21__6_, ab_21__5_,
         ab_21__4_, ab_21__3_, ab_21__2_, ab_21__1_, ab_21__0_, ab_20__23_,
         ab_20__22_, ab_20__21_, ab_20__20_, ab_20__19_, ab_20__18_,
         ab_20__17_, ab_20__16_, ab_20__15_, ab_20__14_, ab_20__13_,
         ab_20__12_, ab_20__11_, ab_20__10_, ab_20__9_, ab_20__8_, ab_20__7_,
         ab_20__6_, ab_20__5_, ab_20__4_, ab_20__3_, ab_20__2_, ab_20__1_,
         ab_20__0_, ab_19__23_, ab_19__22_, ab_19__21_, ab_19__20_, ab_19__19_,
         ab_19__18_, ab_19__17_, ab_19__16_, ab_19__15_, ab_19__14_,
         ab_19__13_, ab_19__12_, ab_19__11_, ab_19__10_, ab_19__9_, ab_19__8_,
         ab_19__7_, ab_19__6_, ab_19__5_, ab_19__4_, ab_19__3_, ab_19__2_,
         ab_19__1_, ab_19__0_, ab_18__23_, ab_18__22_, ab_18__21_, ab_18__20_,
         ab_18__19_, ab_18__18_, ab_18__17_, ab_18__16_, ab_18__15_,
         ab_18__14_, ab_18__13_, ab_18__12_, ab_18__11_, ab_18__10_, ab_18__9_,
         ab_18__8_, ab_18__7_, ab_18__6_, ab_18__5_, ab_18__4_, ab_18__3_,
         ab_18__2_, ab_18__1_, ab_18__0_, ab_17__23_, ab_17__22_, ab_17__21_,
         ab_17__20_, ab_17__19_, ab_17__18_, ab_17__17_, ab_17__16_,
         ab_17__15_, ab_17__14_, ab_17__13_, ab_17__12_, ab_17__11_,
         ab_17__10_, ab_17__9_, ab_17__8_, ab_17__7_, ab_17__6_, ab_17__5_,
         ab_17__4_, ab_17__3_, ab_17__2_, ab_17__1_, ab_17__0_, ab_16__23_,
         ab_16__22_, ab_16__21_, ab_16__20_, ab_16__19_, ab_16__18_,
         ab_16__17_, ab_16__16_, ab_16__15_, ab_16__14_, ab_16__13_,
         ab_16__12_, ab_16__11_, ab_16__10_, ab_16__9_, ab_16__8_, ab_16__7_,
         ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_, ab_16__1_,
         ab_16__0_, ab_15__23_, ab_15__22_, ab_15__21_, ab_15__20_, ab_15__19_,
         ab_15__18_, ab_15__17_, ab_15__16_, ab_15__15_, ab_15__14_,
         ab_15__13_, ab_15__12_, ab_15__11_, ab_15__10_, ab_15__9_, ab_15__8_,
         ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_, ab_15__3_, ab_15__2_,
         ab_15__1_, ab_15__0_, ab_14__23_, ab_14__22_, ab_14__21_, ab_14__20_,
         ab_14__19_, ab_14__18_, ab_14__17_, ab_14__16_, ab_14__15_,
         ab_14__14_, ab_14__13_, ab_14__12_, ab_14__11_, ab_14__10_, ab_14__9_,
         ab_14__8_, ab_14__7_, ab_14__6_, ab_14__5_, ab_14__4_, ab_14__3_,
         ab_14__2_, ab_14__1_, ab_14__0_, ab_13__23_, ab_13__22_, ab_13__21_,
         ab_13__20_, ab_13__19_, ab_13__18_, ab_13__17_, ab_13__16_,
         ab_13__15_, ab_13__14_, ab_13__13_, ab_13__12_, ab_13__11_,
         ab_13__10_, ab_13__9_, ab_13__8_, ab_13__7_, ab_13__6_, ab_13__5_,
         ab_13__4_, ab_13__3_, ab_13__2_, ab_13__1_, ab_13__0_, ab_12__23_,
         ab_12__22_, ab_12__21_, ab_12__20_, ab_12__19_, ab_12__18_,
         ab_12__17_, ab_12__16_, ab_12__15_, ab_12__14_, ab_12__13_,
         ab_12__12_, ab_12__11_, ab_12__10_, ab_12__9_, ab_12__8_, ab_12__7_,
         ab_12__6_, ab_12__5_, ab_12__4_, ab_12__3_, ab_12__2_, ab_12__1_,
         ab_12__0_, ab_11__23_, ab_11__22_, ab_11__21_, ab_11__20_, ab_11__19_,
         ab_11__18_, ab_11__17_, ab_11__16_, ab_11__15_, ab_11__14_,
         ab_11__13_, ab_11__12_, ab_11__11_, ab_11__10_, ab_11__9_, ab_11__8_,
         ab_11__7_, ab_11__6_, ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_,
         ab_11__1_, ab_11__0_, ab_10__23_, ab_10__22_, ab_10__21_, ab_10__20_,
         ab_10__19_, ab_10__18_, ab_10__17_, ab_10__16_, ab_10__15_,
         ab_10__14_, ab_10__13_, ab_10__12_, ab_10__11_, ab_10__10_, ab_10__9_,
         ab_10__8_, ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_,
         ab_10__2_, ab_10__1_, ab_10__0_, ab_9__23_, ab_9__22_, ab_9__21_,
         ab_9__20_, ab_9__19_, ab_9__18_, ab_9__17_, ab_9__16_, ab_9__15_,
         ab_9__14_, ab_9__13_, ab_9__12_, ab_9__11_, ab_9__10_, ab_9__9_,
         ab_9__8_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_,
         ab_9__1_, ab_9__0_, ab_8__23_, ab_8__22_, ab_8__21_, ab_8__20_,
         ab_8__19_, ab_8__18_, ab_8__17_, ab_8__16_, ab_8__15_, ab_8__14_,
         ab_8__13_, ab_8__12_, ab_8__11_, ab_8__10_, ab_8__9_, ab_8__8_,
         ab_8__7_, ab_8__6_, ab_8__5_, ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_,
         ab_8__0_, ab_7__23_, ab_7__22_, ab_7__21_, ab_7__20_, ab_7__19_,
         ab_7__18_, ab_7__17_, ab_7__16_, ab_7__15_, ab_7__14_, ab_7__13_,
         ab_7__12_, ab_7__11_, ab_7__10_, ab_7__9_, ab_7__8_, ab_7__7_,
         ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_,
         ab_6__23_, ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_, ab_6__18_,
         ab_6__17_, ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_, ab_6__12_,
         ab_6__11_, ab_6__10_, ab_6__9_, ab_6__8_, ab_6__7_, ab_6__6_,
         ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_, ab_5__23_,
         ab_5__22_, ab_5__21_, ab_5__20_, ab_5__19_, ab_5__18_, ab_5__17_,
         ab_5__16_, ab_5__15_, ab_5__14_, ab_5__13_, ab_5__12_, ab_5__11_,
         ab_5__10_, ab_5__9_, ab_5__8_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_,
         ab_5__3_, ab_5__2_, ab_5__1_, ab_5__0_, ab_4__23_, ab_4__22_,
         ab_4__21_, ab_4__20_, ab_4__19_, ab_4__18_, ab_4__17_, ab_4__16_,
         ab_4__15_, ab_4__14_, ab_4__13_, ab_4__12_, ab_4__11_, ab_4__10_,
         ab_4__9_, ab_4__8_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_,
         ab_4__2_, ab_4__1_, ab_4__0_, ab_3__23_, ab_3__22_, ab_3__21_,
         ab_3__20_, ab_3__19_, ab_3__18_, ab_3__17_, ab_3__16_, ab_3__15_,
         ab_3__14_, ab_3__13_, ab_3__12_, ab_3__11_, ab_3__10_, ab_3__9_,
         ab_3__8_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_, ab_3__2_,
         ab_3__1_, ab_3__0_, ab_2__23_, ab_2__22_, ab_2__21_, ab_2__20_,
         ab_2__19_, ab_2__18_, ab_2__17_, ab_2__16_, ab_2__15_, ab_2__14_,
         ab_2__13_, ab_2__12_, ab_2__11_, ab_2__10_, ab_2__9_, ab_2__8_,
         ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_,
         ab_2__0_, ab_1__23_, ab_1__22_, ab_1__21_, ab_1__20_, ab_1__19_,
         ab_1__18_, ab_1__17_, ab_1__16_, ab_1__15_, ab_1__14_, ab_1__13_,
         ab_1__12_, ab_1__11_, ab_1__10_, ab_1__9_, ab_1__8_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_0__23_,
         ab_0__22_, ab_0__21_, ab_0__20_, ab_0__19_, ab_0__18_, ab_0__17_,
         ab_0__16_, ab_0__15_, ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_,
         ab_0__10_, ab_0__9_, ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_23__23_, CARRYB_23__22_, CARRYB_23__21_,
         CARRYB_23__20_, CARRYB_23__19_, CARRYB_23__18_, CARRYB_23__17_,
         CARRYB_23__16_, CARRYB_23__15_, CARRYB_23__14_, CARRYB_23__13_,
         CARRYB_23__12_, CARRYB_23__11_, CARRYB_23__10_, CARRYB_23__9_,
         CARRYB_23__8_, CARRYB_23__7_, CARRYB_23__6_, CARRYB_23__5_,
         CARRYB_23__4_, CARRYB_23__3_, CARRYB_23__2_, CARRYB_23__1_,
         CARRYB_23__0_, CARRYB_22__22_, CARRYB_22__21_, CARRYB_22__20_,
         CARRYB_22__19_, CARRYB_22__18_, CARRYB_22__17_, CARRYB_22__16_,
         CARRYB_22__15_, CARRYB_22__14_, CARRYB_22__13_, CARRYB_22__12_,
         CARRYB_22__11_, CARRYB_22__10_, CARRYB_22__9_, CARRYB_22__8_,
         CARRYB_22__7_, CARRYB_22__6_, CARRYB_22__5_, CARRYB_22__4_,
         CARRYB_22__3_, CARRYB_22__2_, CARRYB_22__1_, CARRYB_22__0_,
         CARRYB_21__22_, CARRYB_21__21_, CARRYB_21__20_, CARRYB_21__19_,
         CARRYB_21__18_, CARRYB_21__17_, CARRYB_21__16_, CARRYB_21__15_,
         CARRYB_21__14_, CARRYB_21__13_, CARRYB_21__12_, CARRYB_21__11_,
         CARRYB_21__10_, CARRYB_21__9_, CARRYB_21__8_, CARRYB_21__7_,
         CARRYB_21__6_, CARRYB_21__5_, CARRYB_21__4_, CARRYB_21__3_,
         CARRYB_21__2_, CARRYB_21__1_, CARRYB_21__0_, CARRYB_20__22_,
         CARRYB_20__21_, CARRYB_20__20_, CARRYB_20__19_, CARRYB_20__18_,
         CARRYB_20__17_, CARRYB_20__16_, CARRYB_20__15_, CARRYB_20__14_,
         CARRYB_20__13_, CARRYB_20__12_, CARRYB_20__11_, CARRYB_20__10_,
         CARRYB_20__9_, CARRYB_20__8_, CARRYB_20__7_, CARRYB_20__6_,
         CARRYB_20__5_, CARRYB_20__4_, CARRYB_20__3_, CARRYB_20__2_,
         CARRYB_20__1_, CARRYB_20__0_, CARRYB_19__22_, CARRYB_19__21_,
         CARRYB_19__20_, CARRYB_19__19_, CARRYB_19__18_, CARRYB_19__17_,
         CARRYB_19__16_, CARRYB_19__15_, CARRYB_19__14_, CARRYB_19__13_,
         CARRYB_19__12_, CARRYB_19__11_, CARRYB_19__10_, CARRYB_19__9_,
         CARRYB_19__8_, CARRYB_19__7_, CARRYB_19__6_, CARRYB_19__5_,
         CARRYB_19__4_, CARRYB_19__3_, CARRYB_19__2_, CARRYB_19__1_,
         CARRYB_19__0_, CARRYB_18__22_, CARRYB_18__21_, CARRYB_18__20_,
         CARRYB_18__19_, CARRYB_18__18_, CARRYB_18__17_, CARRYB_18__16_,
         CARRYB_18__15_, CARRYB_18__14_, CARRYB_18__13_, CARRYB_18__12_,
         CARRYB_18__11_, CARRYB_18__10_, CARRYB_18__9_, CARRYB_18__8_,
         CARRYB_18__7_, CARRYB_18__6_, CARRYB_18__5_, CARRYB_18__4_,
         CARRYB_18__3_, CARRYB_18__2_, CARRYB_18__1_, CARRYB_18__0_,
         CARRYB_17__22_, CARRYB_17__21_, CARRYB_17__20_, CARRYB_17__19_,
         CARRYB_17__18_, CARRYB_17__17_, CARRYB_17__16_, CARRYB_17__15_,
         CARRYB_17__14_, CARRYB_17__13_, CARRYB_17__12_, CARRYB_17__11_,
         CARRYB_17__10_, CARRYB_17__9_, CARRYB_17__8_, CARRYB_17__7_,
         CARRYB_17__6_, CARRYB_17__5_, CARRYB_17__4_, CARRYB_17__3_,
         CARRYB_17__2_, CARRYB_17__1_, CARRYB_17__0_, CARRYB_16__22_,
         CARRYB_16__21_, CARRYB_16__20_, CARRYB_16__19_, CARRYB_16__18_,
         CARRYB_16__17_, CARRYB_16__16_, CARRYB_16__15_, CARRYB_16__14_,
         CARRYB_16__13_, CARRYB_16__12_, CARRYB_16__11_, CARRYB_16__10_,
         CARRYB_16__9_, CARRYB_16__8_, CARRYB_16__7_, CARRYB_16__6_,
         CARRYB_16__5_, CARRYB_16__4_, CARRYB_16__3_, CARRYB_16__2_,
         CARRYB_16__1_, CARRYB_16__0_, CARRYB_15__22_, CARRYB_15__21_,
         CARRYB_15__20_, CARRYB_15__19_, CARRYB_15__18_, CARRYB_15__17_,
         CARRYB_15__16_, CARRYB_15__15_, CARRYB_15__14_, CARRYB_15__13_,
         CARRYB_15__12_, CARRYB_15__11_, CARRYB_15__10_, CARRYB_15__9_,
         CARRYB_15__8_, CARRYB_15__7_, CARRYB_15__6_, CARRYB_15__5_,
         CARRYB_15__4_, CARRYB_15__3_, CARRYB_15__2_, CARRYB_15__1_,
         CARRYB_15__0_, CARRYB_14__22_, CARRYB_14__21_, CARRYB_14__20_,
         CARRYB_14__19_, CARRYB_14__18_, CARRYB_14__17_, CARRYB_14__16_,
         CARRYB_14__15_, CARRYB_14__14_, CARRYB_14__13_, CARRYB_14__12_,
         CARRYB_14__11_, CARRYB_14__10_, CARRYB_14__9_, CARRYB_14__8_,
         CARRYB_14__7_, CARRYB_14__6_, CARRYB_14__5_, CARRYB_14__4_,
         CARRYB_14__3_, CARRYB_14__2_, CARRYB_14__1_, CARRYB_14__0_,
         CARRYB_13__22_, CARRYB_13__21_, CARRYB_13__20_, CARRYB_13__19_,
         CARRYB_13__18_, CARRYB_13__17_, CARRYB_13__16_, CARRYB_13__15_,
         CARRYB_13__14_, CARRYB_13__13_, CARRYB_13__12_, CARRYB_13__11_,
         CARRYB_13__10_, CARRYB_13__9_, CARRYB_13__8_, CARRYB_13__7_,
         CARRYB_13__6_, CARRYB_13__5_, CARRYB_13__4_, CARRYB_13__3_,
         CARRYB_13__2_, CARRYB_13__1_, CARRYB_13__0_, CARRYB_12__22_,
         CARRYB_12__21_, CARRYB_12__20_, CARRYB_12__19_, CARRYB_12__18_,
         CARRYB_12__17_, CARRYB_12__16_, CARRYB_12__15_, CARRYB_12__14_,
         CARRYB_12__13_, CARRYB_12__12_, CARRYB_12__11_, CARRYB_12__10_,
         CARRYB_12__9_, CARRYB_12__8_, CARRYB_12__7_, CARRYB_12__6_,
         CARRYB_12__5_, CARRYB_12__4_, CARRYB_12__3_, CARRYB_12__2_,
         CARRYB_12__1_, CARRYB_12__0_, CARRYB_11__22_, CARRYB_11__21_,
         CARRYB_11__20_, CARRYB_11__19_, CARRYB_11__18_, CARRYB_11__17_,
         CARRYB_11__16_, CARRYB_11__15_, CARRYB_11__14_, CARRYB_11__13_,
         CARRYB_11__12_, CARRYB_11__11_, CARRYB_11__10_, CARRYB_11__9_,
         CARRYB_11__8_, CARRYB_11__7_, CARRYB_11__6_, CARRYB_11__5_,
         CARRYB_11__4_, CARRYB_11__3_, CARRYB_11__2_, CARRYB_11__1_,
         CARRYB_11__0_, CARRYB_10__22_, CARRYB_10__21_, CARRYB_10__20_,
         CARRYB_10__19_, CARRYB_10__18_, CARRYB_10__17_, CARRYB_10__16_,
         CARRYB_10__15_, CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_,
         CARRYB_10__11_, CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_,
         CARRYB_10__7_, CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_,
         CARRYB_10__3_, CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_,
         CARRYB_9__22_, CARRYB_9__21_, CARRYB_9__20_, CARRYB_9__19_,
         CARRYB_9__18_, CARRYB_9__17_, CARRYB_9__16_, CARRYB_9__15_,
         CARRYB_9__14_, CARRYB_9__13_, CARRYB_9__12_, CARRYB_9__11_,
         CARRYB_9__10_, CARRYB_9__9_, CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_,
         CARRYB_9__5_, CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_,
         CARRYB_9__0_, CARRYB_8__22_, CARRYB_8__21_, CARRYB_8__20_,
         CARRYB_8__19_, CARRYB_8__18_, CARRYB_8__17_, CARRYB_8__16_,
         CARRYB_8__15_, CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_,
         CARRYB_8__11_, CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_,
         CARRYB_8__7_, CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_,
         CARRYB_8__2_, CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__22_,
         CARRYB_7__21_, CARRYB_7__20_, CARRYB_7__19_, CARRYB_7__18_,
         CARRYB_7__17_, CARRYB_7__16_, CARRYB_7__15_, CARRYB_7__14_,
         CARRYB_7__13_, CARRYB_7__12_, CARRYB_7__11_, CARRYB_7__10_,
         CARRYB_7__9_, CARRYB_7__8_, CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_,
         CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_,
         CARRYB_6__22_, CARRYB_6__21_, CARRYB_6__20_, CARRYB_6__19_,
         CARRYB_6__18_, CARRYB_6__17_, CARRYB_6__16_, CARRYB_6__15_,
         CARRYB_6__14_, CARRYB_6__13_, CARRYB_6__12_, CARRYB_6__11_,
         CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_, CARRYB_6__7_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__22_, CARRYB_5__21_, CARRYB_5__20_,
         CARRYB_5__19_, CARRYB_5__18_, CARRYB_5__17_, CARRYB_5__16_,
         CARRYB_5__15_, CARRYB_5__14_, CARRYB_5__13_, CARRYB_5__12_,
         CARRYB_5__11_, CARRYB_5__10_, CARRYB_5__9_, CARRYB_5__8_,
         CARRYB_5__7_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__22_,
         CARRYB_4__21_, CARRYB_4__20_, CARRYB_4__19_, CARRYB_4__18_,
         CARRYB_4__17_, CARRYB_4__16_, CARRYB_4__15_, CARRYB_4__14_,
         CARRYB_4__13_, CARRYB_4__12_, CARRYB_4__11_, CARRYB_4__10_,
         CARRYB_4__9_, CARRYB_4__8_, CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__22_, CARRYB_3__21_, CARRYB_3__20_, CARRYB_3__19_,
         CARRYB_3__18_, CARRYB_3__17_, CARRYB_3__16_, CARRYB_3__15_,
         CARRYB_3__14_, CARRYB_3__13_, CARRYB_3__12_, CARRYB_3__11_,
         CARRYB_3__10_, CARRYB_3__9_, CARRYB_3__8_, CARRYB_3__7_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__22_, CARRYB_2__21_, CARRYB_2__20_,
         CARRYB_2__19_, CARRYB_2__18_, CARRYB_2__17_, CARRYB_2__16_,
         CARRYB_2__15_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__22_,
         CARRYB_1__21_, CARRYB_1__20_, CARRYB_1__19_, CARRYB_1__18_,
         CARRYB_1__17_, CARRYB_1__16_, CARRYB_1__15_, CARRYB_1__14_,
         CARRYB_1__13_, CARRYB_1__12_, CARRYB_1__11_, CARRYB_1__10_,
         CARRYB_1__9_, CARRYB_1__8_, CARRYB_1__7_, CARRYB_1__6_, CARRYB_1__5_,
         CARRYB_1__4_, CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_,
         SUMB_23__23_, SUMB_23__22_, SUMB_23__21_, SUMB_23__20_, SUMB_23__19_,
         SUMB_23__18_, SUMB_23__17_, SUMB_23__16_, SUMB_23__15_, SUMB_23__14_,
         SUMB_23__13_, SUMB_23__12_, SUMB_23__11_, SUMB_23__10_, SUMB_23__9_,
         SUMB_23__8_, SUMB_23__7_, SUMB_23__6_, SUMB_23__5_, SUMB_23__4_,
         SUMB_23__3_, SUMB_23__2_, SUMB_23__1_, SUMB_23__0_, SUMB_22__22_,
         SUMB_22__21_, SUMB_22__20_, SUMB_22__19_, SUMB_22__18_, SUMB_22__17_,
         SUMB_22__16_, SUMB_22__15_, SUMB_22__14_, SUMB_22__13_, SUMB_22__12_,
         SUMB_22__11_, SUMB_22__10_, SUMB_22__9_, SUMB_22__8_, SUMB_22__7_,
         SUMB_22__6_, SUMB_22__5_, SUMB_22__4_, SUMB_22__3_, SUMB_22__2_,
         SUMB_22__1_, SUMB_21__22_, SUMB_21__21_, SUMB_21__20_, SUMB_21__19_,
         SUMB_21__18_, SUMB_21__17_, SUMB_21__16_, SUMB_21__15_, SUMB_21__14_,
         SUMB_21__13_, SUMB_21__12_, SUMB_21__11_, SUMB_21__10_, SUMB_21__9_,
         SUMB_21__8_, SUMB_21__7_, SUMB_21__6_, SUMB_21__5_, SUMB_21__4_,
         SUMB_21__3_, SUMB_21__2_, SUMB_21__1_, SUMB_20__22_, SUMB_20__21_,
         SUMB_20__20_, SUMB_20__19_, SUMB_20__18_, SUMB_20__17_, SUMB_20__16_,
         SUMB_20__15_, SUMB_20__14_, SUMB_20__13_, SUMB_20__12_, SUMB_20__11_,
         SUMB_20__10_, SUMB_20__9_, SUMB_20__8_, SUMB_20__7_, SUMB_20__6_,
         SUMB_20__5_, SUMB_20__4_, SUMB_20__3_, SUMB_20__2_, SUMB_20__1_,
         SUMB_19__22_, SUMB_19__21_, SUMB_19__20_, SUMB_19__19_, SUMB_19__18_,
         SUMB_19__17_, SUMB_19__16_, SUMB_19__15_, SUMB_19__14_, SUMB_19__13_,
         SUMB_19__12_, SUMB_19__11_, SUMB_19__10_, SUMB_19__9_, SUMB_19__8_,
         SUMB_19__7_, SUMB_19__6_, SUMB_19__5_, SUMB_19__4_, SUMB_19__3_,
         SUMB_19__2_, SUMB_19__1_, SUMB_18__22_, SUMB_18__21_, SUMB_18__20_,
         SUMB_18__19_, SUMB_18__18_, SUMB_18__17_, SUMB_18__16_, SUMB_18__15_,
         SUMB_18__14_, SUMB_18__13_, SUMB_18__12_, SUMB_18__11_, SUMB_18__10_,
         SUMB_18__9_, SUMB_18__8_, SUMB_18__7_, SUMB_18__6_, SUMB_18__5_,
         SUMB_18__4_, SUMB_18__3_, SUMB_18__2_, SUMB_18__1_, SUMB_17__22_,
         SUMB_17__21_, SUMB_17__20_, SUMB_17__19_, SUMB_17__18_, SUMB_17__17_,
         SUMB_17__16_, SUMB_17__15_, SUMB_17__14_, SUMB_17__13_, SUMB_17__12_,
         SUMB_17__11_, SUMB_17__10_, SUMB_17__9_, SUMB_17__8_, SUMB_17__7_,
         SUMB_17__6_, SUMB_17__5_, SUMB_17__4_, SUMB_17__3_, SUMB_17__2_,
         SUMB_17__1_, SUMB_16__22_, SUMB_16__21_, SUMB_16__20_, SUMB_16__19_,
         SUMB_16__18_, SUMB_16__17_, SUMB_16__16_, SUMB_16__15_, SUMB_16__14_,
         SUMB_16__13_, SUMB_16__12_, SUMB_16__11_, SUMB_16__10_, SUMB_16__9_,
         SUMB_16__8_, SUMB_16__7_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_,
         SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, SUMB_15__22_, SUMB_15__21_,
         SUMB_15__20_, SUMB_15__19_, SUMB_15__18_, SUMB_15__17_, SUMB_15__16_,
         SUMB_15__15_, SUMB_15__14_, SUMB_15__13_, SUMB_15__12_, SUMB_15__11_,
         SUMB_15__10_, SUMB_15__9_, SUMB_15__8_, SUMB_15__7_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_14__22_, SUMB_14__21_, SUMB_14__20_, SUMB_14__19_, SUMB_14__18_,
         SUMB_14__17_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_, SUMB_14__13_,
         SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_, SUMB_14__8_,
         SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_,
         SUMB_14__2_, SUMB_14__1_, SUMB_13__22_, SUMB_13__21_, SUMB_13__20_,
         SUMB_13__19_, SUMB_13__18_, SUMB_13__17_, SUMB_13__16_, SUMB_13__15_,
         SUMB_13__14_, SUMB_13__13_, SUMB_13__12_, SUMB_13__11_, SUMB_13__10_,
         SUMB_13__9_, SUMB_13__8_, SUMB_13__7_, SUMB_13__6_, SUMB_13__5_,
         SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_, SUMB_12__22_,
         SUMB_12__21_, SUMB_12__20_, SUMB_12__19_, SUMB_12__18_, SUMB_12__17_,
         SUMB_12__16_, SUMB_12__15_, SUMB_12__14_, SUMB_12__13_, SUMB_12__12_,
         SUMB_12__11_, SUMB_12__10_, SUMB_12__9_, SUMB_12__8_, SUMB_12__7_,
         SUMB_12__6_, SUMB_12__5_, SUMB_12__4_, SUMB_12__3_, SUMB_12__2_,
         SUMB_12__1_, SUMB_11__22_, SUMB_11__21_, SUMB_11__20_, SUMB_11__19_,
         SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_, SUMB_11__14_,
         SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_, SUMB_11__9_,
         SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_, SUMB_11__4_,
         SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__22_, SUMB_10__21_,
         SUMB_10__20_, SUMB_10__19_, SUMB_10__18_, SUMB_10__17_, SUMB_10__16_,
         SUMB_10__15_, SUMB_10__14_, SUMB_10__13_, SUMB_10__12_, SUMB_10__11_,
         SUMB_10__10_, SUMB_10__9_, SUMB_10__8_, SUMB_10__7_, SUMB_10__6_,
         SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_,
         SUMB_9__22_, SUMB_9__21_, SUMB_9__20_, SUMB_9__19_, SUMB_9__18_,
         SUMB_9__17_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_, SUMB_9__13_,
         SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_, SUMB_9__8_,
         SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_,
         SUMB_9__2_, SUMB_9__1_, SUMB_8__22_, SUMB_8__21_, SUMB_8__20_,
         SUMB_8__19_, SUMB_8__18_, SUMB_8__17_, SUMB_8__16_, SUMB_8__15_,
         SUMB_8__14_, SUMB_8__13_, SUMB_8__12_, SUMB_8__11_, SUMB_8__10_,
         SUMB_8__9_, SUMB_8__8_, SUMB_8__7_, SUMB_8__6_, SUMB_8__5_,
         SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_, SUMB_7__22_,
         SUMB_7__21_, SUMB_7__20_, SUMB_7__19_, SUMB_7__18_, SUMB_7__17_,
         SUMB_7__16_, SUMB_7__15_, SUMB_7__14_, SUMB_7__13_, SUMB_7__12_,
         SUMB_7__11_, SUMB_7__10_, SUMB_7__9_, SUMB_7__8_, SUMB_7__7_,
         SUMB_7__6_, SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_,
         SUMB_7__1_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_, SUMB_6__19_,
         SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_, SUMB_6__14_,
         SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_, SUMB_6__9_,
         SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_,
         SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__22_, SUMB_5__21_,
         SUMB_5__20_, SUMB_5__19_, SUMB_5__18_, SUMB_5__17_, SUMB_5__16_,
         SUMB_5__15_, SUMB_5__14_, SUMB_5__13_, SUMB_5__12_, SUMB_5__11_,
         SUMB_5__10_, SUMB_5__9_, SUMB_5__8_, SUMB_5__7_, SUMB_5__6_,
         SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_,
         SUMB_4__22_, SUMB_4__21_, SUMB_4__20_, SUMB_4__19_, SUMB_4__18_,
         SUMB_4__17_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_, SUMB_4__13_,
         SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_, SUMB_4__8_,
         SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_,
         SUMB_4__2_, SUMB_4__1_, SUMB_3__22_, SUMB_3__21_, SUMB_3__20_,
         SUMB_3__19_, SUMB_3__18_, SUMB_3__17_, SUMB_3__16_, SUMB_3__15_,
         SUMB_3__14_, SUMB_3__13_, SUMB_3__12_, SUMB_3__11_, SUMB_3__10_,
         SUMB_3__9_, SUMB_3__8_, SUMB_3__7_, SUMB_3__6_, SUMB_3__5_,
         SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_, SUMB_2__22_,
         SUMB_2__21_, SUMB_2__20_, SUMB_2__19_, SUMB_2__18_, SUMB_2__17_,
         SUMB_2__16_, SUMB_2__15_, SUMB_2__14_, SUMB_2__13_, SUMB_2__12_,
         SUMB_2__11_, SUMB_2__10_, SUMB_2__9_, SUMB_2__8_, SUMB_2__7_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__22_, SUMB_1__21_, SUMB_1__20_, SUMB_1__19_,
         SUMB_1__18_, SUMB_1__17_, SUMB_1__16_, SUMB_1__15_, SUMB_1__14_,
         SUMB_1__13_, SUMB_1__12_, SUMB_1__11_, SUMB_1__10_, SUMB_1__9_,
         SUMB_1__8_, SUMB_1__7_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_,
         SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, QA, QB, A1_45_, A1_44_, A1_43_,
         A1_42_, A1_41_, A1_40_, A1_39_, A1_38_, A1_37_, A1_36_, A1_35_,
         A1_34_, A1_33_, A1_32_, A1_31_, A1_30_, A1_29_, A1_28_, A1_27_,
         A1_26_, A1_25_, A1_24_, A1_23_, A1_22_, A1_21_, A1_20_, A1_19_,
         A1_18_, A1_17_, A1_16_, A1_15_, A1_14_, A1_13_, A1_12_, A1_11_,
         A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_,
         A1_0_, A2_45_, A2_44_, A2_43_, A2_42_, A2_41_, A2_40_, A2_39_, A2_38_,
         A2_37_, A2_36_, A2_35_, A2_34_, A2_33_, A2_32_, A2_31_, A2_30_,
         A2_29_, A2_28_, A2_27_, A2_26_, A2_25_, A2_24_, A2_23_, A2_22_, n1,
         n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21;

  FA_X1 S14_23_0 ( .A(A[23]), .B(B[23]), .CI(SUMB_23__0_), .CO(A2_22_), .S(
        A1_21_) );
  FA_X1 S4_0 ( .A(ab_23__0_), .B(CARRYB_22__0_), .CI(SUMB_22__1_), .CO(
        CARRYB_23__0_), .S(SUMB_23__0_) );
  FA_X1 S4_1 ( .A(ab_23__1_), .B(CARRYB_22__1_), .CI(SUMB_22__2_), .CO(
        CARRYB_23__1_), .S(SUMB_23__1_) );
  FA_X1 S4_2 ( .A(ab_23__2_), .B(CARRYB_22__2_), .CI(SUMB_22__3_), .CO(
        CARRYB_23__2_), .S(SUMB_23__2_) );
  FA_X1 S4_3 ( .A(ab_23__3_), .B(CARRYB_22__3_), .CI(SUMB_22__4_), .CO(
        CARRYB_23__3_), .S(SUMB_23__3_) );
  FA_X1 S4_4 ( .A(ab_23__4_), .B(CARRYB_22__4_), .CI(SUMB_22__5_), .CO(
        CARRYB_23__4_), .S(SUMB_23__4_) );
  FA_X1 S4_5 ( .A(ab_23__5_), .B(CARRYB_22__5_), .CI(SUMB_22__6_), .CO(
        CARRYB_23__5_), .S(SUMB_23__5_) );
  FA_X1 S4_6 ( .A(ab_23__6_), .B(CARRYB_22__6_), .CI(SUMB_22__7_), .CO(
        CARRYB_23__6_), .S(SUMB_23__6_) );
  FA_X1 S4_7 ( .A(ab_23__7_), .B(CARRYB_22__7_), .CI(SUMB_22__8_), .CO(
        CARRYB_23__7_), .S(SUMB_23__7_) );
  FA_X1 S4_8 ( .A(ab_23__8_), .B(CARRYB_22__8_), .CI(SUMB_22__9_), .CO(
        CARRYB_23__8_), .S(SUMB_23__8_) );
  FA_X1 S4_9 ( .A(ab_23__9_), .B(CARRYB_22__9_), .CI(SUMB_22__10_), .CO(
        CARRYB_23__9_), .S(SUMB_23__9_) );
  FA_X1 S4_10 ( .A(ab_23__10_), .B(CARRYB_22__10_), .CI(SUMB_22__11_), .CO(
        CARRYB_23__10_), .S(SUMB_23__10_) );
  FA_X1 S4_11 ( .A(ab_23__11_), .B(CARRYB_22__11_), .CI(SUMB_22__12_), .CO(
        CARRYB_23__11_), .S(SUMB_23__11_) );
  FA_X1 S4_12 ( .A(ab_23__12_), .B(CARRYB_22__12_), .CI(SUMB_22__13_), .CO(
        CARRYB_23__12_), .S(SUMB_23__12_) );
  FA_X1 S4_13 ( .A(ab_23__13_), .B(CARRYB_22__13_), .CI(SUMB_22__14_), .CO(
        CARRYB_23__13_), .S(SUMB_23__13_) );
  FA_X1 S4_14 ( .A(ab_23__14_), .B(CARRYB_22__14_), .CI(SUMB_22__15_), .CO(
        CARRYB_23__14_), .S(SUMB_23__14_) );
  FA_X1 S4_15 ( .A(ab_23__15_), .B(CARRYB_22__15_), .CI(SUMB_22__16_), .CO(
        CARRYB_23__15_), .S(SUMB_23__15_) );
  FA_X1 S4_16 ( .A(ab_23__16_), .B(CARRYB_22__16_), .CI(SUMB_22__17_), .CO(
        CARRYB_23__16_), .S(SUMB_23__16_) );
  FA_X1 S4_17 ( .A(ab_23__17_), .B(CARRYB_22__17_), .CI(SUMB_22__18_), .CO(
        CARRYB_23__17_), .S(SUMB_23__17_) );
  FA_X1 S4_18 ( .A(ab_23__18_), .B(CARRYB_22__18_), .CI(SUMB_22__19_), .CO(
        CARRYB_23__18_), .S(SUMB_23__18_) );
  FA_X1 S4_19 ( .A(ab_23__19_), .B(CARRYB_22__19_), .CI(SUMB_22__20_), .CO(
        CARRYB_23__19_), .S(SUMB_23__19_) );
  FA_X1 S4_20 ( .A(ab_23__20_), .B(CARRYB_22__20_), .CI(SUMB_22__21_), .CO(
        CARRYB_23__20_), .S(SUMB_23__20_) );
  FA_X1 S4_21 ( .A(ab_23__21_), .B(CARRYB_22__21_), .CI(SUMB_22__22_), .CO(
        CARRYB_23__21_), .S(SUMB_23__21_) );
  FA_X1 S5_22 ( .A(ab_23__22_), .B(CARRYB_22__22_), .CI(ab_22__23_), .CO(
        CARRYB_23__22_), .S(SUMB_23__22_) );
  FA_X1 S14_23 ( .A(n3), .B(n1), .CI(ab_23__23_), .CO(CARRYB_23__23_), .S(
        SUMB_23__23_) );
  FA_X1 S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), .CO(
        CARRYB_22__0_), .S(A1_20_) );
  FA_X1 S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), .CO(
        CARRYB_22__1_), .S(SUMB_22__1_) );
  FA_X1 S2_22_2 ( .A(ab_22__2_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), .CO(
        CARRYB_22__2_), .S(SUMB_22__2_) );
  FA_X1 S2_22_3 ( .A(ab_22__3_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), .CO(
        CARRYB_22__3_), .S(SUMB_22__3_) );
  FA_X1 S2_22_4 ( .A(ab_22__4_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), .CO(
        CARRYB_22__4_), .S(SUMB_22__4_) );
  FA_X1 S2_22_5 ( .A(ab_22__5_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), .CO(
        CARRYB_22__5_), .S(SUMB_22__5_) );
  FA_X1 S2_22_6 ( .A(ab_22__6_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), .CO(
        CARRYB_22__6_), .S(SUMB_22__6_) );
  FA_X1 S2_22_7 ( .A(ab_22__7_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), .CO(
        CARRYB_22__7_), .S(SUMB_22__7_) );
  FA_X1 S2_22_8 ( .A(ab_22__8_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), .CO(
        CARRYB_22__8_), .S(SUMB_22__8_) );
  FA_X1 S2_22_9 ( .A(ab_22__9_), .B(CARRYB_21__9_), .CI(SUMB_21__10_), .CO(
        CARRYB_22__9_), .S(SUMB_22__9_) );
  FA_X1 S2_22_10 ( .A(ab_22__10_), .B(CARRYB_21__10_), .CI(SUMB_21__11_), .CO(
        CARRYB_22__10_), .S(SUMB_22__10_) );
  FA_X1 S2_22_11 ( .A(ab_22__11_), .B(CARRYB_21__11_), .CI(SUMB_21__12_), .CO(
        CARRYB_22__11_), .S(SUMB_22__11_) );
  FA_X1 S2_22_12 ( .A(ab_22__12_), .B(CARRYB_21__12_), .CI(SUMB_21__13_), .CO(
        CARRYB_22__12_), .S(SUMB_22__12_) );
  FA_X1 S2_22_13 ( .A(ab_22__13_), .B(CARRYB_21__13_), .CI(SUMB_21__14_), .CO(
        CARRYB_22__13_), .S(SUMB_22__13_) );
  FA_X1 S2_22_14 ( .A(ab_22__14_), .B(CARRYB_21__14_), .CI(SUMB_21__15_), .CO(
        CARRYB_22__14_), .S(SUMB_22__14_) );
  FA_X1 S2_22_15 ( .A(ab_22__15_), .B(CARRYB_21__15_), .CI(SUMB_21__16_), .CO(
        CARRYB_22__15_), .S(SUMB_22__15_) );
  FA_X1 S2_22_16 ( .A(ab_22__16_), .B(CARRYB_21__16_), .CI(SUMB_21__17_), .CO(
        CARRYB_22__16_), .S(SUMB_22__16_) );
  FA_X1 S2_22_17 ( .A(ab_22__17_), .B(CARRYB_21__17_), .CI(SUMB_21__18_), .CO(
        CARRYB_22__17_), .S(SUMB_22__17_) );
  FA_X1 S2_22_18 ( .A(ab_22__18_), .B(CARRYB_21__18_), .CI(SUMB_21__19_), .CO(
        CARRYB_22__18_), .S(SUMB_22__18_) );
  FA_X1 S2_22_19 ( .A(ab_22__19_), .B(CARRYB_21__19_), .CI(SUMB_21__20_), .CO(
        CARRYB_22__19_), .S(SUMB_22__19_) );
  FA_X1 S2_22_20 ( .A(ab_22__20_), .B(CARRYB_21__20_), .CI(SUMB_21__21_), .CO(
        CARRYB_22__20_), .S(SUMB_22__20_) );
  FA_X1 S2_22_21 ( .A(ab_22__21_), .B(CARRYB_21__21_), .CI(SUMB_21__22_), .CO(
        CARRYB_22__21_), .S(SUMB_22__21_) );
  FA_X1 S3_22_22 ( .A(ab_22__22_), .B(CARRYB_21__22_), .CI(ab_21__23_), .CO(
        CARRYB_22__22_), .S(SUMB_22__22_) );
  FA_X1 S1_21_0 ( .A(ab_21__0_), .B(CARRYB_20__0_), .CI(SUMB_20__1_), .CO(
        CARRYB_21__0_), .S(A1_19_) );
  FA_X1 S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), .CO(
        CARRYB_21__1_), .S(SUMB_21__1_) );
  FA_X1 S2_21_2 ( .A(ab_21__2_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), .CO(
        CARRYB_21__2_), .S(SUMB_21__2_) );
  FA_X1 S2_21_3 ( .A(ab_21__3_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), .CO(
        CARRYB_21__3_), .S(SUMB_21__3_) );
  FA_X1 S2_21_4 ( .A(ab_21__4_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), .CO(
        CARRYB_21__4_), .S(SUMB_21__4_) );
  FA_X1 S2_21_5 ( .A(ab_21__5_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), .CO(
        CARRYB_21__5_), .S(SUMB_21__5_) );
  FA_X1 S2_21_6 ( .A(ab_21__6_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), .CO(
        CARRYB_21__6_), .S(SUMB_21__6_) );
  FA_X1 S2_21_7 ( .A(ab_21__7_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), .CO(
        CARRYB_21__7_), .S(SUMB_21__7_) );
  FA_X1 S2_21_8 ( .A(ab_21__8_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), .CO(
        CARRYB_21__8_), .S(SUMB_21__8_) );
  FA_X1 S2_21_9 ( .A(ab_21__9_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), .CO(
        CARRYB_21__9_), .S(SUMB_21__9_) );
  FA_X1 S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .CI(SUMB_20__11_), .CO(
        CARRYB_21__10_), .S(SUMB_21__10_) );
  FA_X1 S2_21_11 ( .A(ab_21__11_), .B(CARRYB_20__11_), .CI(SUMB_20__12_), .CO(
        CARRYB_21__11_), .S(SUMB_21__11_) );
  FA_X1 S2_21_12 ( .A(ab_21__12_), .B(CARRYB_20__12_), .CI(SUMB_20__13_), .CO(
        CARRYB_21__12_), .S(SUMB_21__12_) );
  FA_X1 S2_21_13 ( .A(ab_21__13_), .B(CARRYB_20__13_), .CI(SUMB_20__14_), .CO(
        CARRYB_21__13_), .S(SUMB_21__13_) );
  FA_X1 S2_21_14 ( .A(ab_21__14_), .B(CARRYB_20__14_), .CI(SUMB_20__15_), .CO(
        CARRYB_21__14_), .S(SUMB_21__14_) );
  FA_X1 S2_21_15 ( .A(ab_21__15_), .B(CARRYB_20__15_), .CI(SUMB_20__16_), .CO(
        CARRYB_21__15_), .S(SUMB_21__15_) );
  FA_X1 S2_21_16 ( .A(ab_21__16_), .B(CARRYB_20__16_), .CI(SUMB_20__17_), .CO(
        CARRYB_21__16_), .S(SUMB_21__16_) );
  FA_X1 S2_21_17 ( .A(ab_21__17_), .B(CARRYB_20__17_), .CI(SUMB_20__18_), .CO(
        CARRYB_21__17_), .S(SUMB_21__17_) );
  FA_X1 S2_21_18 ( .A(ab_21__18_), .B(CARRYB_20__18_), .CI(SUMB_20__19_), .CO(
        CARRYB_21__18_), .S(SUMB_21__18_) );
  FA_X1 S2_21_19 ( .A(ab_21__19_), .B(CARRYB_20__19_), .CI(SUMB_20__20_), .CO(
        CARRYB_21__19_), .S(SUMB_21__19_) );
  FA_X1 S2_21_20 ( .A(ab_21__20_), .B(CARRYB_20__20_), .CI(SUMB_20__21_), .CO(
        CARRYB_21__20_), .S(SUMB_21__20_) );
  FA_X1 S2_21_21 ( .A(ab_21__21_), .B(CARRYB_20__21_), .CI(SUMB_20__22_), .CO(
        CARRYB_21__21_), .S(SUMB_21__21_) );
  FA_X1 S3_21_22 ( .A(ab_21__22_), .B(CARRYB_20__22_), .CI(ab_20__23_), .CO(
        CARRYB_21__22_), .S(SUMB_21__22_) );
  FA_X1 S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), .CO(
        CARRYB_20__0_), .S(A1_18_) );
  FA_X1 S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), .CO(
        CARRYB_20__1_), .S(SUMB_20__1_) );
  FA_X1 S2_20_2 ( .A(ab_20__2_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), .CO(
        CARRYB_20__2_), .S(SUMB_20__2_) );
  FA_X1 S2_20_3 ( .A(ab_20__3_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), .CO(
        CARRYB_20__3_), .S(SUMB_20__3_) );
  FA_X1 S2_20_4 ( .A(ab_20__4_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), .CO(
        CARRYB_20__4_), .S(SUMB_20__4_) );
  FA_X1 S2_20_5 ( .A(ab_20__5_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), .CO(
        CARRYB_20__5_), .S(SUMB_20__5_) );
  FA_X1 S2_20_6 ( .A(ab_20__6_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), .CO(
        CARRYB_20__6_), .S(SUMB_20__6_) );
  FA_X1 S2_20_7 ( .A(ab_20__7_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), .CO(
        CARRYB_20__7_), .S(SUMB_20__7_) );
  FA_X1 S2_20_8 ( .A(ab_20__8_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), .CO(
        CARRYB_20__8_), .S(SUMB_20__8_) );
  FA_X1 S2_20_9 ( .A(ab_20__9_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), .CO(
        CARRYB_20__9_), .S(SUMB_20__9_) );
  FA_X1 S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), .CO(
        CARRYB_20__10_), .S(SUMB_20__10_) );
  FA_X1 S2_20_11 ( .A(ab_20__11_), .B(CARRYB_19__11_), .CI(SUMB_19__12_), .CO(
        CARRYB_20__11_), .S(SUMB_20__11_) );
  FA_X1 S2_20_12 ( .A(ab_20__12_), .B(CARRYB_19__12_), .CI(SUMB_19__13_), .CO(
        CARRYB_20__12_), .S(SUMB_20__12_) );
  FA_X1 S2_20_13 ( .A(ab_20__13_), .B(CARRYB_19__13_), .CI(SUMB_19__14_), .CO(
        CARRYB_20__13_), .S(SUMB_20__13_) );
  FA_X1 S2_20_14 ( .A(ab_20__14_), .B(CARRYB_19__14_), .CI(SUMB_19__15_), .CO(
        CARRYB_20__14_), .S(SUMB_20__14_) );
  FA_X1 S2_20_15 ( .A(ab_20__15_), .B(CARRYB_19__15_), .CI(SUMB_19__16_), .CO(
        CARRYB_20__15_), .S(SUMB_20__15_) );
  FA_X1 S2_20_16 ( .A(ab_20__16_), .B(CARRYB_19__16_), .CI(SUMB_19__17_), .CO(
        CARRYB_20__16_), .S(SUMB_20__16_) );
  FA_X1 S2_20_17 ( .A(ab_20__17_), .B(CARRYB_19__17_), .CI(SUMB_19__18_), .CO(
        CARRYB_20__17_), .S(SUMB_20__17_) );
  FA_X1 S2_20_18 ( .A(ab_20__18_), .B(CARRYB_19__18_), .CI(SUMB_19__19_), .CO(
        CARRYB_20__18_), .S(SUMB_20__18_) );
  FA_X1 S2_20_19 ( .A(ab_20__19_), .B(CARRYB_19__19_), .CI(SUMB_19__20_), .CO(
        CARRYB_20__19_), .S(SUMB_20__19_) );
  FA_X1 S2_20_20 ( .A(ab_20__20_), .B(CARRYB_19__20_), .CI(SUMB_19__21_), .CO(
        CARRYB_20__20_), .S(SUMB_20__20_) );
  FA_X1 S2_20_21 ( .A(ab_20__21_), .B(CARRYB_19__21_), .CI(SUMB_19__22_), .CO(
        CARRYB_20__21_), .S(SUMB_20__21_) );
  FA_X1 S3_20_22 ( .A(ab_20__22_), .B(CARRYB_19__22_), .CI(ab_19__23_), .CO(
        CARRYB_20__22_), .S(SUMB_20__22_) );
  FA_X1 S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), .CO(
        CARRYB_19__0_), .S(A1_17_) );
  FA_X1 S2_19_1 ( .A(ab_19__1_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), .CO(
        CARRYB_19__1_), .S(SUMB_19__1_) );
  FA_X1 S2_19_2 ( .A(ab_19__2_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), .CO(
        CARRYB_19__2_), .S(SUMB_19__2_) );
  FA_X1 S2_19_3 ( .A(ab_19__3_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), .CO(
        CARRYB_19__3_), .S(SUMB_19__3_) );
  FA_X1 S2_19_4 ( .A(ab_19__4_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), .CO(
        CARRYB_19__4_), .S(SUMB_19__4_) );
  FA_X1 S2_19_5 ( .A(ab_19__5_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), .CO(
        CARRYB_19__5_), .S(SUMB_19__5_) );
  FA_X1 S2_19_6 ( .A(ab_19__6_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), .CO(
        CARRYB_19__6_), .S(SUMB_19__6_) );
  FA_X1 S2_19_7 ( .A(ab_19__7_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), .CO(
        CARRYB_19__7_), .S(SUMB_19__7_) );
  FA_X1 S2_19_8 ( .A(ab_19__8_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), .CO(
        CARRYB_19__8_), .S(SUMB_19__8_) );
  FA_X1 S2_19_9 ( .A(ab_19__9_), .B(CARRYB_18__9_), .CI(SUMB_18__10_), .CO(
        CARRYB_19__9_), .S(SUMB_19__9_) );
  FA_X1 S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), .CO(
        CARRYB_19__10_), .S(SUMB_19__10_) );
  FA_X1 S2_19_11 ( .A(ab_19__11_), .B(CARRYB_18__11_), .CI(SUMB_18__12_), .CO(
        CARRYB_19__11_), .S(SUMB_19__11_) );
  FA_X1 S2_19_12 ( .A(ab_19__12_), .B(CARRYB_18__12_), .CI(SUMB_18__13_), .CO(
        CARRYB_19__12_), .S(SUMB_19__12_) );
  FA_X1 S2_19_13 ( .A(ab_19__13_), .B(CARRYB_18__13_), .CI(SUMB_18__14_), .CO(
        CARRYB_19__13_), .S(SUMB_19__13_) );
  FA_X1 S2_19_14 ( .A(ab_19__14_), .B(CARRYB_18__14_), .CI(SUMB_18__15_), .CO(
        CARRYB_19__14_), .S(SUMB_19__14_) );
  FA_X1 S2_19_15 ( .A(ab_19__15_), .B(CARRYB_18__15_), .CI(SUMB_18__16_), .CO(
        CARRYB_19__15_), .S(SUMB_19__15_) );
  FA_X1 S2_19_16 ( .A(ab_19__16_), .B(CARRYB_18__16_), .CI(SUMB_18__17_), .CO(
        CARRYB_19__16_), .S(SUMB_19__16_) );
  FA_X1 S2_19_17 ( .A(ab_19__17_), .B(CARRYB_18__17_), .CI(SUMB_18__18_), .CO(
        CARRYB_19__17_), .S(SUMB_19__17_) );
  FA_X1 S2_19_18 ( .A(ab_19__18_), .B(CARRYB_18__18_), .CI(SUMB_18__19_), .CO(
        CARRYB_19__18_), .S(SUMB_19__18_) );
  FA_X1 S2_19_19 ( .A(ab_19__19_), .B(CARRYB_18__19_), .CI(SUMB_18__20_), .CO(
        CARRYB_19__19_), .S(SUMB_19__19_) );
  FA_X1 S2_19_20 ( .A(ab_19__20_), .B(CARRYB_18__20_), .CI(SUMB_18__21_), .CO(
        CARRYB_19__20_), .S(SUMB_19__20_) );
  FA_X1 S2_19_21 ( .A(ab_19__21_), .B(CARRYB_18__21_), .CI(SUMB_18__22_), .CO(
        CARRYB_19__21_), .S(SUMB_19__21_) );
  FA_X1 S3_19_22 ( .A(ab_19__22_), .B(CARRYB_18__22_), .CI(ab_18__23_), .CO(
        CARRYB_19__22_), .S(SUMB_19__22_) );
  FA_X1 S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), .CO(
        CARRYB_18__0_), .S(A1_16_) );
  FA_X1 S2_18_1 ( .A(ab_18__1_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), .CO(
        CARRYB_18__1_), .S(SUMB_18__1_) );
  FA_X1 S2_18_2 ( .A(ab_18__2_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), .CO(
        CARRYB_18__2_), .S(SUMB_18__2_) );
  FA_X1 S2_18_3 ( .A(ab_18__3_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), .CO(
        CARRYB_18__3_), .S(SUMB_18__3_) );
  FA_X1 S2_18_4 ( .A(ab_18__4_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), .CO(
        CARRYB_18__4_), .S(SUMB_18__4_) );
  FA_X1 S2_18_5 ( .A(ab_18__5_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), .CO(
        CARRYB_18__5_), .S(SUMB_18__5_) );
  FA_X1 S2_18_6 ( .A(ab_18__6_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), .CO(
        CARRYB_18__6_), .S(SUMB_18__6_) );
  FA_X1 S2_18_7 ( .A(ab_18__7_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), .CO(
        CARRYB_18__7_), .S(SUMB_18__7_) );
  FA_X1 S2_18_8 ( .A(ab_18__8_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), .CO(
        CARRYB_18__8_), .S(SUMB_18__8_) );
  FA_X1 S2_18_9 ( .A(ab_18__9_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), .CO(
        CARRYB_18__9_), .S(SUMB_18__9_) );
  FA_X1 S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), .CO(
        CARRYB_18__10_), .S(SUMB_18__10_) );
  FA_X1 S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), .CO(
        CARRYB_18__11_), .S(SUMB_18__11_) );
  FA_X1 S2_18_12 ( .A(ab_18__12_), .B(CARRYB_17__12_), .CI(SUMB_17__13_), .CO(
        CARRYB_18__12_), .S(SUMB_18__12_) );
  FA_X1 S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .CI(SUMB_17__14_), .CO(
        CARRYB_18__13_), .S(SUMB_18__13_) );
  FA_X1 S2_18_14 ( .A(ab_18__14_), .B(CARRYB_17__14_), .CI(SUMB_17__15_), .CO(
        CARRYB_18__14_), .S(SUMB_18__14_) );
  FA_X1 S2_18_15 ( .A(ab_18__15_), .B(CARRYB_17__15_), .CI(SUMB_17__16_), .CO(
        CARRYB_18__15_), .S(SUMB_18__15_) );
  FA_X1 S2_18_16 ( .A(ab_18__16_), .B(CARRYB_17__16_), .CI(SUMB_17__17_), .CO(
        CARRYB_18__16_), .S(SUMB_18__16_) );
  FA_X1 S2_18_17 ( .A(ab_18__17_), .B(CARRYB_17__17_), .CI(SUMB_17__18_), .CO(
        CARRYB_18__17_), .S(SUMB_18__17_) );
  FA_X1 S2_18_18 ( .A(ab_18__18_), .B(CARRYB_17__18_), .CI(SUMB_17__19_), .CO(
        CARRYB_18__18_), .S(SUMB_18__18_) );
  FA_X1 S2_18_19 ( .A(ab_18__19_), .B(CARRYB_17__19_), .CI(SUMB_17__20_), .CO(
        CARRYB_18__19_), .S(SUMB_18__19_) );
  FA_X1 S2_18_20 ( .A(ab_18__20_), .B(CARRYB_17__20_), .CI(SUMB_17__21_), .CO(
        CARRYB_18__20_), .S(SUMB_18__20_) );
  FA_X1 S2_18_21 ( .A(ab_18__21_), .B(CARRYB_17__21_), .CI(SUMB_17__22_), .CO(
        CARRYB_18__21_), .S(SUMB_18__21_) );
  FA_X1 S3_18_22 ( .A(ab_18__22_), .B(CARRYB_17__22_), .CI(ab_17__23_), .CO(
        CARRYB_18__22_), .S(SUMB_18__22_) );
  FA_X1 S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), .CO(
        CARRYB_17__0_), .S(A1_15_) );
  FA_X1 S2_17_1 ( .A(ab_17__1_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), .CO(
        CARRYB_17__1_), .S(SUMB_17__1_) );
  FA_X1 S2_17_2 ( .A(ab_17__2_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), .CO(
        CARRYB_17__2_), .S(SUMB_17__2_) );
  FA_X1 S2_17_3 ( .A(ab_17__3_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), .CO(
        CARRYB_17__3_), .S(SUMB_17__3_) );
  FA_X1 S2_17_4 ( .A(ab_17__4_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), .CO(
        CARRYB_17__4_), .S(SUMB_17__4_) );
  FA_X1 S2_17_5 ( .A(ab_17__5_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), .CO(
        CARRYB_17__5_), .S(SUMB_17__5_) );
  FA_X1 S2_17_6 ( .A(ab_17__6_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), .CO(
        CARRYB_17__6_), .S(SUMB_17__6_) );
  FA_X1 S2_17_7 ( .A(ab_17__7_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), .CO(
        CARRYB_17__7_), .S(SUMB_17__7_) );
  FA_X1 S2_17_8 ( .A(ab_17__8_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), .CO(
        CARRYB_17__8_), .S(SUMB_17__8_) );
  FA_X1 S2_17_9 ( .A(ab_17__9_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), .CO(
        CARRYB_17__9_), .S(SUMB_17__9_) );
  FA_X1 S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), .CO(
        CARRYB_17__10_), .S(SUMB_17__10_) );
  FA_X1 S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), .CO(
        CARRYB_17__11_), .S(SUMB_17__11_) );
  FA_X1 S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), .CO(
        CARRYB_17__12_), .S(SUMB_17__12_) );
  FA_X1 S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), .CO(
        CARRYB_17__13_), .S(SUMB_17__13_) );
  FA_X1 S2_17_14 ( .A(ab_17__14_), .B(CARRYB_16__14_), .CI(SUMB_16__15_), .CO(
        CARRYB_17__14_), .S(SUMB_17__14_) );
  FA_X1 S2_17_15 ( .A(ab_17__15_), .B(CARRYB_16__15_), .CI(SUMB_16__16_), .CO(
        CARRYB_17__15_), .S(SUMB_17__15_) );
  FA_X1 S2_17_16 ( .A(ab_17__16_), .B(CARRYB_16__16_), .CI(SUMB_16__17_), .CO(
        CARRYB_17__16_), .S(SUMB_17__16_) );
  FA_X1 S2_17_17 ( .A(ab_17__17_), .B(CARRYB_16__17_), .CI(SUMB_16__18_), .CO(
        CARRYB_17__17_), .S(SUMB_17__17_) );
  FA_X1 S2_17_18 ( .A(ab_17__18_), .B(CARRYB_16__18_), .CI(SUMB_16__19_), .CO(
        CARRYB_17__18_), .S(SUMB_17__18_) );
  FA_X1 S2_17_19 ( .A(ab_17__19_), .B(CARRYB_16__19_), .CI(SUMB_16__20_), .CO(
        CARRYB_17__19_), .S(SUMB_17__19_) );
  FA_X1 S2_17_20 ( .A(ab_17__20_), .B(CARRYB_16__20_), .CI(SUMB_16__21_), .CO(
        CARRYB_17__20_), .S(SUMB_17__20_) );
  FA_X1 S2_17_21 ( .A(ab_17__21_), .B(CARRYB_16__21_), .CI(SUMB_16__22_), .CO(
        CARRYB_17__21_), .S(SUMB_17__21_) );
  FA_X1 S3_17_22 ( .A(ab_17__22_), .B(CARRYB_16__22_), .CI(ab_16__23_), .CO(
        CARRYB_17__22_), .S(SUMB_17__22_) );
  FA_X1 S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(A1_14_) );
  FA_X1 S2_16_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  FA_X1 S2_16_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  FA_X1 S2_16_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  FA_X1 S2_16_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  FA_X1 S2_16_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  FA_X1 S2_16_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  FA_X1 S2_16_7 ( .A(ab_16__7_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), .CO(
        CARRYB_16__7_), .S(SUMB_16__7_) );
  FA_X1 S2_16_8 ( .A(ab_16__8_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), .CO(
        CARRYB_16__8_), .S(SUMB_16__8_) );
  FA_X1 S2_16_9 ( .A(ab_16__9_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), .CO(
        CARRYB_16__9_), .S(SUMB_16__9_) );
  FA_X1 S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), .CO(
        CARRYB_16__10_), .S(SUMB_16__10_) );
  FA_X1 S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), .CO(
        CARRYB_16__11_), .S(SUMB_16__11_) );
  FA_X1 S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), .CO(
        CARRYB_16__12_), .S(SUMB_16__12_) );
  FA_X1 S2_16_13 ( .A(ab_16__13_), .B(CARRYB_15__13_), .CI(SUMB_15__14_), .CO(
        CARRYB_16__13_), .S(SUMB_16__13_) );
  FA_X1 S2_16_14 ( .A(ab_16__14_), .B(CARRYB_15__14_), .CI(SUMB_15__15_), .CO(
        CARRYB_16__14_), .S(SUMB_16__14_) );
  FA_X1 S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .CI(SUMB_15__16_), .CO(
        CARRYB_16__15_), .S(SUMB_16__15_) );
  FA_X1 S2_16_16 ( .A(ab_16__16_), .B(CARRYB_15__16_), .CI(SUMB_15__17_), .CO(
        CARRYB_16__16_), .S(SUMB_16__16_) );
  FA_X1 S2_16_17 ( .A(ab_16__17_), .B(CARRYB_15__17_), .CI(SUMB_15__18_), .CO(
        CARRYB_16__17_), .S(SUMB_16__17_) );
  FA_X1 S2_16_18 ( .A(ab_16__18_), .B(CARRYB_15__18_), .CI(SUMB_15__19_), .CO(
        CARRYB_16__18_), .S(SUMB_16__18_) );
  FA_X1 S2_16_19 ( .A(ab_16__19_), .B(CARRYB_15__19_), .CI(SUMB_15__20_), .CO(
        CARRYB_16__19_), .S(SUMB_16__19_) );
  FA_X1 S2_16_20 ( .A(ab_16__20_), .B(CARRYB_15__20_), .CI(SUMB_15__21_), .CO(
        CARRYB_16__20_), .S(SUMB_16__20_) );
  FA_X1 S2_16_21 ( .A(ab_16__21_), .B(CARRYB_15__21_), .CI(SUMB_15__22_), .CO(
        CARRYB_16__21_), .S(SUMB_16__21_) );
  FA_X1 S3_16_22 ( .A(ab_16__22_), .B(CARRYB_15__22_), .CI(ab_15__23_), .CO(
        CARRYB_16__22_), .S(SUMB_16__22_) );
  FA_X1 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  FA_X1 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  FA_X1 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  FA_X1 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  FA_X1 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  FA_X1 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  FA_X1 S2_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  FA_X1 S2_15_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), .CO(
        CARRYB_15__7_), .S(SUMB_15__7_) );
  FA_X1 S2_15_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), .CO(
        CARRYB_15__8_), .S(SUMB_15__8_) );
  FA_X1 S2_15_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), .CO(
        CARRYB_15__9_), .S(SUMB_15__9_) );
  FA_X1 S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), .CO(
        CARRYB_15__10_), .S(SUMB_15__10_) );
  FA_X1 S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), .CO(
        CARRYB_15__11_), .S(SUMB_15__11_) );
  FA_X1 S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), .CO(
        CARRYB_15__12_), .S(SUMB_15__12_) );
  FA_X1 S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), .CO(
        CARRYB_15__13_), .S(SUMB_15__13_) );
  FA_X1 S2_15_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), .CO(
        CARRYB_15__14_), .S(SUMB_15__14_) );
  FA_X1 S2_15_15 ( .A(ab_15__15_), .B(CARRYB_14__15_), .CI(SUMB_14__16_), .CO(
        CARRYB_15__15_), .S(SUMB_15__15_) );
  FA_X1 S2_15_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .CI(SUMB_14__17_), .CO(
        CARRYB_15__16_), .S(SUMB_15__16_) );
  FA_X1 S2_15_17 ( .A(ab_15__17_), .B(CARRYB_14__17_), .CI(SUMB_14__18_), .CO(
        CARRYB_15__17_), .S(SUMB_15__17_) );
  FA_X1 S2_15_18 ( .A(ab_15__18_), .B(CARRYB_14__18_), .CI(SUMB_14__19_), .CO(
        CARRYB_15__18_), .S(SUMB_15__18_) );
  FA_X1 S2_15_19 ( .A(ab_15__19_), .B(CARRYB_14__19_), .CI(SUMB_14__20_), .CO(
        CARRYB_15__19_), .S(SUMB_15__19_) );
  FA_X1 S2_15_20 ( .A(ab_15__20_), .B(CARRYB_14__20_), .CI(SUMB_14__21_), .CO(
        CARRYB_15__20_), .S(SUMB_15__20_) );
  FA_X1 S2_15_21 ( .A(ab_15__21_), .B(CARRYB_14__21_), .CI(SUMB_14__22_), .CO(
        CARRYB_15__21_), .S(SUMB_15__21_) );
  FA_X1 S3_15_22 ( .A(ab_15__22_), .B(CARRYB_14__22_), .CI(ab_14__23_), .CO(
        CARRYB_15__22_), .S(SUMB_15__22_) );
  FA_X1 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  FA_X1 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  FA_X1 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  FA_X1 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  FA_X1 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  FA_X1 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  FA_X1 S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  FA_X1 S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), .CO(
        CARRYB_14__7_), .S(SUMB_14__7_) );
  FA_X1 S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), .CO(
        CARRYB_14__8_), .S(SUMB_14__8_) );
  FA_X1 S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), .CO(
        CARRYB_14__9_), .S(SUMB_14__9_) );
  FA_X1 S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), .CO(
        CARRYB_14__10_), .S(SUMB_14__10_) );
  FA_X1 S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), .CO(
        CARRYB_14__11_), .S(SUMB_14__11_) );
  FA_X1 S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), .CO(
        CARRYB_14__12_), .S(SUMB_14__12_) );
  FA_X1 S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), .CO(
        CARRYB_14__13_), .S(SUMB_14__13_) );
  FA_X1 S2_14_14 ( .A(ab_14__14_), .B(CARRYB_13__14_), .CI(SUMB_13__15_), .CO(
        CARRYB_14__14_), .S(SUMB_14__14_) );
  FA_X1 S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), .CO(
        CARRYB_14__15_), .S(SUMB_14__15_) );
  FA_X1 S2_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), .CO(
        CARRYB_14__16_), .S(SUMB_14__16_) );
  FA_X1 S2_14_17 ( .A(ab_14__17_), .B(CARRYB_13__17_), .CI(SUMB_13__18_), .CO(
        CARRYB_14__17_), .S(SUMB_14__17_) );
  FA_X1 S2_14_18 ( .A(ab_14__18_), .B(CARRYB_13__18_), .CI(SUMB_13__19_), .CO(
        CARRYB_14__18_), .S(SUMB_14__18_) );
  FA_X1 S2_14_19 ( .A(ab_14__19_), .B(CARRYB_13__19_), .CI(SUMB_13__20_), .CO(
        CARRYB_14__19_), .S(SUMB_14__19_) );
  FA_X1 S2_14_20 ( .A(ab_14__20_), .B(CARRYB_13__20_), .CI(SUMB_13__21_), .CO(
        CARRYB_14__20_), .S(SUMB_14__20_) );
  FA_X1 S2_14_21 ( .A(ab_14__21_), .B(CARRYB_13__21_), .CI(SUMB_13__22_), .CO(
        CARRYB_14__21_), .S(SUMB_14__21_) );
  FA_X1 S3_14_22 ( .A(ab_14__22_), .B(CARRYB_13__22_), .CI(ab_13__23_), .CO(
        CARRYB_14__22_), .S(SUMB_14__22_) );
  FA_X1 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  FA_X1 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  FA_X1 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  FA_X1 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  FA_X1 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  FA_X1 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  FA_X1 S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  FA_X1 S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), .CO(
        CARRYB_13__7_), .S(SUMB_13__7_) );
  FA_X1 S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), .CO(
        CARRYB_13__8_), .S(SUMB_13__8_) );
  FA_X1 S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), .CO(
        CARRYB_13__9_), .S(SUMB_13__9_) );
  FA_X1 S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), .CO(
        CARRYB_13__10_), .S(SUMB_13__10_) );
  FA_X1 S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), .CO(
        CARRYB_13__11_), .S(SUMB_13__11_) );
  FA_X1 S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), .CO(
        CARRYB_13__12_), .S(SUMB_13__12_) );
  FA_X1 S2_13_13 ( .A(ab_13__13_), .B(CARRYB_12__13_), .CI(SUMB_12__14_), .CO(
        CARRYB_13__13_), .S(SUMB_13__13_) );
  FA_X1 S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), .CO(
        CARRYB_13__14_), .S(SUMB_13__14_) );
  FA_X1 S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), .CO(
        CARRYB_13__15_), .S(SUMB_13__15_) );
  FA_X1 S2_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), .CO(
        CARRYB_13__16_), .S(SUMB_13__16_) );
  FA_X1 S2_13_17 ( .A(ab_13__17_), .B(CARRYB_12__17_), .CI(SUMB_12__18_), .CO(
        CARRYB_13__17_), .S(SUMB_13__17_) );
  FA_X1 S2_13_18 ( .A(ab_13__18_), .B(CARRYB_12__18_), .CI(SUMB_12__19_), .CO(
        CARRYB_13__18_), .S(SUMB_13__18_) );
  FA_X1 S2_13_19 ( .A(ab_13__19_), .B(CARRYB_12__19_), .CI(SUMB_12__20_), .CO(
        CARRYB_13__19_), .S(SUMB_13__19_) );
  FA_X1 S2_13_20 ( .A(ab_13__20_), .B(CARRYB_12__20_), .CI(SUMB_12__21_), .CO(
        CARRYB_13__20_), .S(SUMB_13__20_) );
  FA_X1 S2_13_21 ( .A(ab_13__21_), .B(CARRYB_12__21_), .CI(SUMB_12__22_), .CO(
        CARRYB_13__21_), .S(SUMB_13__21_) );
  FA_X1 S3_13_22 ( .A(ab_13__22_), .B(CARRYB_12__22_), .CI(ab_12__23_), .CO(
        CARRYB_13__22_), .S(SUMB_13__22_) );
  FA_X1 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  FA_X1 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  FA_X1 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  FA_X1 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  FA_X1 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  FA_X1 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  FA_X1 S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  FA_X1 S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), .CO(
        CARRYB_12__7_), .S(SUMB_12__7_) );
  FA_X1 S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), .CO(
        CARRYB_12__8_), .S(SUMB_12__8_) );
  FA_X1 S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), .CO(
        CARRYB_12__9_), .S(SUMB_12__9_) );
  FA_X1 S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), .CO(
        CARRYB_12__10_), .S(SUMB_12__10_) );
  FA_X1 S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), .CO(
        CARRYB_12__11_), .S(SUMB_12__11_) );
  FA_X1 S2_12_12 ( .A(ab_12__12_), .B(CARRYB_11__12_), .CI(SUMB_11__13_), .CO(
        CARRYB_12__12_), .S(SUMB_12__12_) );
  FA_X1 S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), .CO(
        CARRYB_12__13_), .S(SUMB_12__13_) );
  FA_X1 S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), .CO(
        CARRYB_12__14_), .S(SUMB_12__14_) );
  FA_X1 S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), .CO(
        CARRYB_12__15_), .S(SUMB_12__15_) );
  FA_X1 S2_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), .CO(
        CARRYB_12__16_), .S(SUMB_12__16_) );
  FA_X1 S2_12_17 ( .A(ab_12__17_), .B(CARRYB_11__17_), .CI(SUMB_11__18_), .CO(
        CARRYB_12__17_), .S(SUMB_12__17_) );
  FA_X1 S2_12_18 ( .A(ab_12__18_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), .CO(
        CARRYB_12__18_), .S(SUMB_12__18_) );
  FA_X1 S2_12_19 ( .A(ab_12__19_), .B(CARRYB_11__19_), .CI(SUMB_11__20_), .CO(
        CARRYB_12__19_), .S(SUMB_12__19_) );
  FA_X1 S2_12_20 ( .A(ab_12__20_), .B(CARRYB_11__20_), .CI(SUMB_11__21_), .CO(
        CARRYB_12__20_), .S(SUMB_12__20_) );
  FA_X1 S2_12_21 ( .A(ab_12__21_), .B(CARRYB_11__21_), .CI(SUMB_11__22_), .CO(
        CARRYB_12__21_), .S(SUMB_12__21_) );
  FA_X1 S3_12_22 ( .A(ab_12__22_), .B(CARRYB_11__22_), .CI(ab_11__23_), .CO(
        CARRYB_12__22_), .S(SUMB_12__22_) );
  FA_X1 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  FA_X1 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  FA_X1 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  FA_X1 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  FA_X1 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  FA_X1 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  FA_X1 S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  FA_X1 S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), .CO(
        CARRYB_11__7_), .S(SUMB_11__7_) );
  FA_X1 S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), .CO(
        CARRYB_11__8_), .S(SUMB_11__8_) );
  FA_X1 S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), .CO(
        CARRYB_11__9_), .S(SUMB_11__9_) );
  FA_X1 S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), .CO(
        CARRYB_11__10_), .S(SUMB_11__10_) );
  FA_X1 S2_11_11 ( .A(ab_11__11_), .B(CARRYB_10__11_), .CI(SUMB_10__12_), .CO(
        CARRYB_11__11_), .S(SUMB_11__11_) );
  FA_X1 S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), .CO(
        CARRYB_11__12_), .S(SUMB_11__12_) );
  FA_X1 S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), .CO(
        CARRYB_11__13_), .S(SUMB_11__13_) );
  FA_X1 S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), .CO(
        CARRYB_11__14_), .S(SUMB_11__14_) );
  FA_X1 S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), .CO(
        CARRYB_11__15_), .S(SUMB_11__15_) );
  FA_X1 S2_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(SUMB_10__17_), .CO(
        CARRYB_11__16_), .S(SUMB_11__16_) );
  FA_X1 S2_11_17 ( .A(ab_11__17_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), .CO(
        CARRYB_11__17_), .S(SUMB_11__17_) );
  FA_X1 S2_11_18 ( .A(ab_11__18_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), .CO(
        CARRYB_11__18_), .S(SUMB_11__18_) );
  FA_X1 S2_11_19 ( .A(ab_11__19_), .B(CARRYB_10__19_), .CI(SUMB_10__20_), .CO(
        CARRYB_11__19_), .S(SUMB_11__19_) );
  FA_X1 S2_11_20 ( .A(ab_11__20_), .B(CARRYB_10__20_), .CI(SUMB_10__21_), .CO(
        CARRYB_11__20_), .S(SUMB_11__20_) );
  FA_X1 S2_11_21 ( .A(ab_11__21_), .B(CARRYB_10__21_), .CI(SUMB_10__22_), .CO(
        CARRYB_11__21_), .S(SUMB_11__21_) );
  FA_X1 S3_11_22 ( .A(ab_11__22_), .B(CARRYB_10__22_), .CI(ab_10__23_), .CO(
        CARRYB_11__22_), .S(SUMB_11__22_) );
  FA_X1 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  FA_X1 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  FA_X1 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  FA_X1 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  FA_X1 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  FA_X1 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  FA_X1 S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  FA_X1 S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  FA_X1 S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  FA_X1 S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  FA_X1 S2_10_10 ( .A(ab_10__10_), .B(CARRYB_9__10_), .CI(SUMB_9__11_), .CO(
        CARRYB_10__10_), .S(SUMB_10__10_) );
  FA_X1 S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), .CO(
        CARRYB_10__11_), .S(SUMB_10__11_) );
  FA_X1 S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), .CO(
        CARRYB_10__12_), .S(SUMB_10__12_) );
  FA_X1 S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), .CO(
        CARRYB_10__13_), .S(SUMB_10__13_) );
  FA_X1 S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), .CO(
        CARRYB_10__14_), .S(SUMB_10__14_) );
  FA_X1 S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), .CO(
        CARRYB_10__15_), .S(SUMB_10__15_) );
  FA_X1 S2_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), .CO(
        CARRYB_10__16_), .S(SUMB_10__16_) );
  FA_X1 S2_10_17 ( .A(ab_10__17_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), .CO(
        CARRYB_10__17_), .S(SUMB_10__17_) );
  FA_X1 S2_10_18 ( .A(ab_10__18_), .B(CARRYB_9__18_), .CI(SUMB_9__19_), .CO(
        CARRYB_10__18_), .S(SUMB_10__18_) );
  FA_X1 S2_10_19 ( .A(ab_10__19_), .B(CARRYB_9__19_), .CI(SUMB_9__20_), .CO(
        CARRYB_10__19_), .S(SUMB_10__19_) );
  FA_X1 S2_10_20 ( .A(ab_10__20_), .B(CARRYB_9__20_), .CI(SUMB_9__21_), .CO(
        CARRYB_10__20_), .S(SUMB_10__20_) );
  FA_X1 S2_10_21 ( .A(ab_10__21_), .B(CARRYB_9__21_), .CI(SUMB_9__22_), .CO(
        CARRYB_10__21_), .S(SUMB_10__21_) );
  FA_X1 S3_10_22 ( .A(ab_10__22_), .B(CARRYB_9__22_), .CI(ab_9__23_), .CO(
        CARRYB_10__22_), .S(SUMB_10__22_) );
  FA_X1 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  FA_X1 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  FA_X1 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  FA_X1 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  FA_X1 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  FA_X1 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  FA_X1 S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  FA_X1 S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  FA_X1 S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  FA_X1 S2_9_9 ( .A(ab_9__9_), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  FA_X1 S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), .CO(
        CARRYB_9__10_), .S(SUMB_9__10_) );
  FA_X1 S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), .CO(
        CARRYB_9__11_), .S(SUMB_9__11_) );
  FA_X1 S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), .CO(
        CARRYB_9__12_), .S(SUMB_9__12_) );
  FA_X1 S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), .CO(
        CARRYB_9__13_), .S(SUMB_9__13_) );
  FA_X1 S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), .CO(
        CARRYB_9__14_), .S(SUMB_9__14_) );
  FA_X1 S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), .CO(
        CARRYB_9__15_), .S(SUMB_9__15_) );
  FA_X1 S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), .CO(
        CARRYB_9__16_), .S(SUMB_9__16_) );
  FA_X1 S2_9_17 ( .A(ab_9__17_), .B(CARRYB_8__17_), .CI(SUMB_8__18_), .CO(
        CARRYB_9__17_), .S(SUMB_9__17_) );
  FA_X1 S2_9_18 ( .A(ab_9__18_), .B(CARRYB_8__18_), .CI(SUMB_8__19_), .CO(
        CARRYB_9__18_), .S(SUMB_9__18_) );
  FA_X1 S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), .CO(
        CARRYB_9__19_), .S(SUMB_9__19_) );
  FA_X1 S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(SUMB_8__21_), .CO(
        CARRYB_9__20_), .S(SUMB_9__20_) );
  FA_X1 S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), .CO(
        CARRYB_9__21_), .S(SUMB_9__21_) );
  FA_X1 S3_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .CI(ab_8__23_), .CO(
        CARRYB_9__22_), .S(SUMB_9__22_) );
  FA_X1 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  FA_X1 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  FA_X1 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  FA_X1 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  FA_X1 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  FA_X1 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  FA_X1 S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  FA_X1 S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  FA_X1 S2_8_8 ( .A(ab_8__8_), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  FA_X1 S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  FA_X1 S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), .CO(
        CARRYB_8__10_), .S(SUMB_8__10_) );
  FA_X1 S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), .CO(
        CARRYB_8__11_), .S(SUMB_8__11_) );
  FA_X1 S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), .CO(
        CARRYB_8__12_), .S(SUMB_8__12_) );
  FA_X1 S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), .CO(
        CARRYB_8__13_), .S(SUMB_8__13_) );
  FA_X1 S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), .CO(
        CARRYB_8__14_), .S(SUMB_8__14_) );
  FA_X1 S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), .CO(
        CARRYB_8__15_), .S(SUMB_8__15_) );
  FA_X1 S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), .CO(
        CARRYB_8__16_), .S(SUMB_8__16_) );
  FA_X1 S2_8_17 ( .A(ab_8__17_), .B(CARRYB_7__17_), .CI(SUMB_7__18_), .CO(
        CARRYB_8__17_), .S(SUMB_8__17_) );
  FA_X1 S2_8_18 ( .A(ab_8__18_), .B(CARRYB_7__18_), .CI(SUMB_7__19_), .CO(
        CARRYB_8__18_), .S(SUMB_8__18_) );
  FA_X1 S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), .CO(
        CARRYB_8__19_), .S(SUMB_8__19_) );
  FA_X1 S2_8_20 ( .A(ab_8__20_), .B(CARRYB_7__20_), .CI(SUMB_7__21_), .CO(
        CARRYB_8__20_), .S(SUMB_8__20_) );
  FA_X1 S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), .CO(
        CARRYB_8__21_), .S(SUMB_8__21_) );
  FA_X1 S3_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(ab_7__23_), .CO(
        CARRYB_8__22_), .S(SUMB_8__22_) );
  FA_X1 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(A1_5_) );
  FA_X1 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S2_7_7 ( .A(ab_7__7_), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  FA_X1 S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  FA_X1 S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  FA_X1 S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), .CO(
        CARRYB_7__10_), .S(SUMB_7__10_) );
  FA_X1 S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), .CO(
        CARRYB_7__11_), .S(SUMB_7__11_) );
  FA_X1 S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), .CO(
        CARRYB_7__12_), .S(SUMB_7__12_) );
  FA_X1 S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), .CO(
        CARRYB_7__13_), .S(SUMB_7__13_) );
  FA_X1 S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), .CO(
        CARRYB_7__14_), .S(SUMB_7__14_) );
  FA_X1 S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), .CO(
        CARRYB_7__15_), .S(SUMB_7__15_) );
  FA_X1 S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), .CO(
        CARRYB_7__16_), .S(SUMB_7__16_) );
  FA_X1 S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), .CO(
        CARRYB_7__17_), .S(SUMB_7__17_) );
  FA_X1 S2_7_18 ( .A(ab_7__18_), .B(CARRYB_6__18_), .CI(SUMB_6__19_), .CO(
        CARRYB_7__18_), .S(SUMB_7__18_) );
  FA_X1 S2_7_19 ( .A(ab_7__19_), .B(CARRYB_6__19_), .CI(SUMB_6__20_), .CO(
        CARRYB_7__19_), .S(SUMB_7__19_) );
  FA_X1 S2_7_20 ( .A(ab_7__20_), .B(CARRYB_6__20_), .CI(SUMB_6__21_), .CO(
        CARRYB_7__20_), .S(SUMB_7__20_) );
  FA_X1 S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), .CO(
        CARRYB_7__21_), .S(SUMB_7__21_) );
  FA_X1 S3_7_22 ( .A(ab_7__22_), .B(CARRYB_6__22_), .CI(ab_6__23_), .CO(
        CARRYB_7__22_), .S(SUMB_7__22_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S2_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  FA_X1 S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  FA_X1 S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  FA_X1 S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), .CO(
        CARRYB_6__10_), .S(SUMB_6__10_) );
  FA_X1 S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), .CO(
        CARRYB_6__11_), .S(SUMB_6__11_) );
  FA_X1 S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), .CO(
        CARRYB_6__12_), .S(SUMB_6__12_) );
  FA_X1 S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), .CO(
        CARRYB_6__13_), .S(SUMB_6__13_) );
  FA_X1 S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), .CO(
        CARRYB_6__14_), .S(SUMB_6__14_) );
  FA_X1 S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), .CO(
        CARRYB_6__15_), .S(SUMB_6__15_) );
  FA_X1 S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), .CO(
        CARRYB_6__16_), .S(SUMB_6__16_) );
  FA_X1 S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), .CO(
        CARRYB_6__17_), .S(SUMB_6__17_) );
  FA_X1 S2_6_18 ( .A(ab_6__18_), .B(CARRYB_5__18_), .CI(SUMB_5__19_), .CO(
        CARRYB_6__18_), .S(SUMB_6__18_) );
  FA_X1 S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), .CO(
        CARRYB_6__19_), .S(SUMB_6__19_) );
  FA_X1 S2_6_20 ( .A(ab_6__20_), .B(CARRYB_5__20_), .CI(SUMB_5__21_), .CO(
        CARRYB_6__20_), .S(SUMB_6__20_) );
  FA_X1 S2_6_21 ( .A(ab_6__21_), .B(CARRYB_5__21_), .CI(SUMB_5__22_), .CO(
        CARRYB_6__21_), .S(SUMB_6__21_) );
  FA_X1 S3_6_22 ( .A(ab_6__22_), .B(CARRYB_5__22_), .CI(ab_5__23_), .CO(
        CARRYB_6__22_), .S(SUMB_6__22_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  FA_X1 S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  FA_X1 S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  FA_X1 S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), .CO(
        CARRYB_5__10_), .S(SUMB_5__10_) );
  FA_X1 S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), .CO(
        CARRYB_5__11_), .S(SUMB_5__11_) );
  FA_X1 S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), .CO(
        CARRYB_5__12_), .S(SUMB_5__12_) );
  FA_X1 S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), .CO(
        CARRYB_5__13_), .S(SUMB_5__13_) );
  FA_X1 S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), .CO(
        CARRYB_5__14_), .S(SUMB_5__14_) );
  FA_X1 S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), .CO(
        CARRYB_5__15_), .S(SUMB_5__15_) );
  FA_X1 S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), .CO(
        CARRYB_5__16_), .S(SUMB_5__16_) );
  FA_X1 S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), .CO(
        CARRYB_5__17_), .S(SUMB_5__17_) );
  FA_X1 S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), .CO(
        CARRYB_5__18_), .S(SUMB_5__18_) );
  FA_X1 S2_5_19 ( .A(ab_5__19_), .B(CARRYB_4__19_), .CI(SUMB_4__20_), .CO(
        CARRYB_5__19_), .S(SUMB_5__19_) );
  FA_X1 S2_5_20 ( .A(ab_5__20_), .B(CARRYB_4__20_), .CI(SUMB_4__21_), .CO(
        CARRYB_5__20_), .S(SUMB_5__20_) );
  FA_X1 S2_5_21 ( .A(ab_5__21_), .B(CARRYB_4__21_), .CI(SUMB_4__22_), .CO(
        CARRYB_5__21_), .S(SUMB_5__21_) );
  FA_X1 S3_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(ab_4__23_), .CO(
        CARRYB_5__22_), .S(SUMB_5__22_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  FA_X1 S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  FA_X1 S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  FA_X1 S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), .CO(
        CARRYB_4__10_), .S(SUMB_4__10_) );
  FA_X1 S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), .CO(
        CARRYB_4__11_), .S(SUMB_4__11_) );
  FA_X1 S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), .CO(
        CARRYB_4__12_), .S(SUMB_4__12_) );
  FA_X1 S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), .CO(
        CARRYB_4__13_), .S(SUMB_4__13_) );
  FA_X1 S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), .CO(
        CARRYB_4__14_), .S(SUMB_4__14_) );
  FA_X1 S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), .CO(
        CARRYB_4__15_), .S(SUMB_4__15_) );
  FA_X1 S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), .CO(
        CARRYB_4__16_), .S(SUMB_4__16_) );
  FA_X1 S2_4_17 ( .A(ab_4__17_), .B(CARRYB_3__17_), .CI(SUMB_3__18_), .CO(
        CARRYB_4__17_), .S(SUMB_4__17_) );
  FA_X1 S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), .CO(
        CARRYB_4__18_), .S(SUMB_4__18_) );
  FA_X1 S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), .CO(
        CARRYB_4__19_), .S(SUMB_4__19_) );
  FA_X1 S2_4_20 ( .A(ab_4__20_), .B(CARRYB_3__20_), .CI(SUMB_3__21_), .CO(
        CARRYB_4__20_), .S(SUMB_4__20_) );
  FA_X1 S2_4_21 ( .A(ab_4__21_), .B(CARRYB_3__21_), .CI(SUMB_3__22_), .CO(
        CARRYB_4__21_), .S(SUMB_4__21_) );
  FA_X1 S3_4_22 ( .A(ab_4__22_), .B(CARRYB_3__22_), .CI(ab_3__23_), .CO(
        CARRYB_4__22_), .S(SUMB_4__22_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  FA_X1 S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  FA_X1 S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  FA_X1 S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), .CO(
        CARRYB_3__10_), .S(SUMB_3__10_) );
  FA_X1 S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), .CO(
        CARRYB_3__11_), .S(SUMB_3__11_) );
  FA_X1 S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), .CO(
        CARRYB_3__12_), .S(SUMB_3__12_) );
  FA_X1 S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), .CO(
        CARRYB_3__13_), .S(SUMB_3__13_) );
  FA_X1 S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), .CO(
        CARRYB_3__14_), .S(SUMB_3__14_) );
  FA_X1 S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), .CO(
        CARRYB_3__15_), .S(SUMB_3__15_) );
  FA_X1 S2_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(SUMB_2__17_), .CO(
        CARRYB_3__16_), .S(SUMB_3__16_) );
  FA_X1 S2_3_17 ( .A(ab_3__17_), .B(CARRYB_2__17_), .CI(SUMB_2__18_), .CO(
        CARRYB_3__17_), .S(SUMB_3__17_) );
  FA_X1 S2_3_18 ( .A(ab_3__18_), .B(CARRYB_2__18_), .CI(SUMB_2__19_), .CO(
        CARRYB_3__18_), .S(SUMB_3__18_) );
  FA_X1 S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), .CO(
        CARRYB_3__19_), .S(SUMB_3__19_) );
  FA_X1 S2_3_20 ( .A(ab_3__20_), .B(CARRYB_2__20_), .CI(SUMB_2__21_), .CO(
        CARRYB_3__20_), .S(SUMB_3__20_) );
  FA_X1 S2_3_21 ( .A(ab_3__21_), .B(CARRYB_2__21_), .CI(SUMB_2__22_), .CO(
        CARRYB_3__21_), .S(SUMB_3__21_) );
  FA_X1 S3_3_22 ( .A(ab_3__22_), .B(CARRYB_2__22_), .CI(ab_2__23_), .CO(
        CARRYB_3__22_), .S(SUMB_3__22_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S2_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(SUMB_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  FA_X1 S2_2_7 ( .A(ab_2__7_), .B(CARRYB_1__7_), .CI(SUMB_1__8_), .CO(
        CARRYB_2__7_), .S(SUMB_2__7_) );
  FA_X1 S2_2_8 ( .A(ab_2__8_), .B(CARRYB_1__8_), .CI(SUMB_1__9_), .CO(
        CARRYB_2__8_), .S(SUMB_2__8_) );
  FA_X1 S2_2_9 ( .A(ab_2__9_), .B(CARRYB_1__9_), .CI(SUMB_1__10_), .CO(
        CARRYB_2__9_), .S(SUMB_2__9_) );
  FA_X1 S2_2_10 ( .A(ab_2__10_), .B(CARRYB_1__10_), .CI(SUMB_1__11_), .CO(
        CARRYB_2__10_), .S(SUMB_2__10_) );
  FA_X1 S2_2_11 ( .A(ab_2__11_), .B(CARRYB_1__11_), .CI(SUMB_1__12_), .CO(
        CARRYB_2__11_), .S(SUMB_2__11_) );
  FA_X1 S2_2_12 ( .A(ab_2__12_), .B(CARRYB_1__12_), .CI(SUMB_1__13_), .CO(
        CARRYB_2__12_), .S(SUMB_2__12_) );
  FA_X1 S2_2_13 ( .A(ab_2__13_), .B(CARRYB_1__13_), .CI(SUMB_1__14_), .CO(
        CARRYB_2__13_), .S(SUMB_2__13_) );
  FA_X1 S2_2_14 ( .A(ab_2__14_), .B(CARRYB_1__14_), .CI(SUMB_1__15_), .CO(
        CARRYB_2__14_), .S(SUMB_2__14_) );
  FA_X1 S2_2_15 ( .A(ab_2__15_), .B(CARRYB_1__15_), .CI(SUMB_1__16_), .CO(
        CARRYB_2__15_), .S(SUMB_2__15_) );
  FA_X1 S2_2_16 ( .A(ab_2__16_), .B(CARRYB_1__16_), .CI(SUMB_1__17_), .CO(
        CARRYB_2__16_), .S(SUMB_2__16_) );
  FA_X1 S2_2_17 ( .A(ab_2__17_), .B(CARRYB_1__17_), .CI(SUMB_1__18_), .CO(
        CARRYB_2__17_), .S(SUMB_2__17_) );
  FA_X1 S2_2_18 ( .A(ab_2__18_), .B(CARRYB_1__18_), .CI(SUMB_1__19_), .CO(
        CARRYB_2__18_), .S(SUMB_2__18_) );
  FA_X1 S2_2_19 ( .A(ab_2__19_), .B(CARRYB_1__19_), .CI(SUMB_1__20_), .CO(
        CARRYB_2__19_), .S(SUMB_2__19_) );
  FA_X1 S2_2_20 ( .A(ab_2__20_), .B(CARRYB_1__20_), .CI(SUMB_1__21_), .CO(
        CARRYB_2__20_), .S(SUMB_2__20_) );
  FA_X1 S2_2_21 ( .A(ab_2__21_), .B(CARRYB_1__21_), .CI(SUMB_1__22_), .CO(
        CARRYB_2__21_), .S(SUMB_2__21_) );
  FA_X1 S3_2_22 ( .A(ab_2__22_), .B(CARRYB_1__22_), .CI(ab_1__23_), .CO(
        CARRYB_2__22_), .S(SUMB_2__22_) );
  iir_filter_DW01_add_4 FS_1 ( .A({A1_45_, A1_44_, A1_43_, A1_42_, A1_41_, 
        A1_40_, A1_39_, A1_38_, A1_37_, A1_36_, A1_35_, A1_34_, A1_33_, A1_32_, 
        A1_31_, A1_30_, A1_29_, A1_28_, A1_27_, A1_26_, A1_25_, A1_24_, A1_23_, 
        A1_22_, A1_21_, A1_20_, A1_19_, A1_18_, A1_17_, A1_16_, A1_15_, A1_14_, 
        A1_13_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, A1_5_, 
        A1_4_, A1_3_, A1_2_, A1_1_, A1_0_}), .B({A2_45_, A2_44_, A2_43_, 
        A2_42_, A2_41_, A2_40_, A2_39_, A2_38_, A2_37_, A2_36_, A2_35_, A2_34_, 
        A2_33_, A2_32_, A2_31_, A2_30_, A2_29_, A2_28_, A2_27_, A2_26_, A2_25_, 
        A2_24_, A2_23_, A2_22_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({PRODUCT[47], SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, PRODUCT[44:22], SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21}) );
  BUF_X1 U2 ( .A(QB), .Z(n1) );
  BUF_X1 U3 ( .A(QB), .Z(n2) );
  BUF_X1 U4 ( .A(QA), .Z(n3) );
  BUF_X1 U5 ( .A(QA), .Z(n4) );
  INV_X1 U6 ( .A(A[2]), .ZN(n36) );
  INV_X1 U7 ( .A(A[3]), .ZN(n35) );
  INV_X1 U8 ( .A(A[4]), .ZN(n34) );
  INV_X1 U9 ( .A(A[5]), .ZN(n33) );
  INV_X1 U10 ( .A(A[6]), .ZN(n32) );
  INV_X1 U11 ( .A(B[1]), .ZN(n18) );
  INV_X1 U12 ( .A(A[1]), .ZN(n40) );
  INV_X1 U13 ( .A(B[0]), .ZN(n29) );
  INV_X1 U14 ( .A(A[0]), .ZN(n51) );
  INV_X1 U15 ( .A(B[22]), .ZN(n15) );
  INV_X1 U16 ( .A(B[21]), .ZN(n16) );
  INV_X1 U17 ( .A(B[20]), .ZN(n17) );
  INV_X1 U18 ( .A(B[19]), .ZN(n19) );
  INV_X1 U19 ( .A(B[18]), .ZN(n20) );
  INV_X1 U20 ( .A(B[17]), .ZN(n21) );
  INV_X1 U21 ( .A(B[16]), .ZN(n22) );
  INV_X1 U22 ( .A(B[15]), .ZN(n23) );
  INV_X1 U23 ( .A(B[14]), .ZN(n24) );
  INV_X1 U24 ( .A(B[13]), .ZN(n25) );
  INV_X1 U25 ( .A(B[12]), .ZN(n26) );
  INV_X1 U26 ( .A(B[11]), .ZN(n27) );
  INV_X1 U27 ( .A(B[10]), .ZN(n28) );
  INV_X1 U28 ( .A(B[9]), .ZN(n7) );
  INV_X1 U29 ( .A(B[8]), .ZN(n8) );
  INV_X1 U30 ( .A(B[7]), .ZN(n9) );
  INV_X1 U31 ( .A(B[6]), .ZN(n10) );
  INV_X1 U32 ( .A(B[5]), .ZN(n11) );
  INV_X1 U33 ( .A(B[4]), .ZN(n12) );
  INV_X1 U34 ( .A(B[3]), .ZN(n13) );
  INV_X1 U35 ( .A(B[2]), .ZN(n14) );
  INV_X1 U36 ( .A(A[7]), .ZN(n31) );
  INV_X1 U37 ( .A(A[8]), .ZN(n30) );
  INV_X1 U38 ( .A(A[10]), .ZN(n50) );
  INV_X1 U39 ( .A(A[11]), .ZN(n49) );
  INV_X1 U40 ( .A(A[12]), .ZN(n48) );
  INV_X1 U41 ( .A(A[13]), .ZN(n47) );
  INV_X1 U42 ( .A(A[14]), .ZN(n46) );
  INV_X1 U43 ( .A(A[9]), .ZN(n6) );
  INV_X1 U44 ( .A(A[22]), .ZN(n37) );
  INV_X1 U45 ( .A(A[15]), .ZN(n45) );
  INV_X1 U46 ( .A(A[16]), .ZN(n44) );
  INV_X1 U47 ( .A(A[17]), .ZN(n43) );
  INV_X1 U48 ( .A(A[18]), .ZN(n42) );
  INV_X1 U49 ( .A(A[19]), .ZN(n41) );
  INV_X1 U50 ( .A(A[20]), .ZN(n39) );
  INV_X1 U51 ( .A(A[21]), .ZN(n38) );
  AND2_X1 U52 ( .A1(SUMB_23__23_), .A2(CARRYB_23__22_), .ZN(A2_45_) );
  XOR2_X1 U53 ( .A(CARRYB_23__22_), .B(SUMB_23__23_), .Z(A1_44_) );
  AND2_X1 U54 ( .A1(SUMB_23__22_), .A2(CARRYB_23__21_), .ZN(A2_44_) );
  XOR2_X1 U55 ( .A(CARRYB_23__21_), .B(SUMB_23__22_), .Z(A1_43_) );
  AND2_X1 U56 ( .A1(SUMB_23__21_), .A2(CARRYB_23__20_), .ZN(A2_43_) );
  XOR2_X1 U57 ( .A(CARRYB_23__20_), .B(SUMB_23__21_), .Z(A1_42_) );
  AND2_X1 U58 ( .A1(SUMB_23__20_), .A2(CARRYB_23__19_), .ZN(A2_42_) );
  XOR2_X1 U59 ( .A(CARRYB_23__19_), .B(SUMB_23__20_), .Z(A1_41_) );
  AND2_X1 U60 ( .A1(SUMB_23__19_), .A2(CARRYB_23__18_), .ZN(A2_41_) );
  XOR2_X1 U61 ( .A(CARRYB_23__18_), .B(SUMB_23__19_), .Z(A1_40_) );
  AND2_X1 U62 ( .A1(SUMB_23__18_), .A2(CARRYB_23__17_), .ZN(A2_40_) );
  XOR2_X1 U63 ( .A(CARRYB_23__17_), .B(SUMB_23__18_), .Z(A1_39_) );
  AND2_X1 U64 ( .A1(SUMB_23__17_), .A2(CARRYB_23__16_), .ZN(A2_39_) );
  XOR2_X1 U65 ( .A(CARRYB_23__16_), .B(SUMB_23__17_), .Z(A1_38_) );
  AND2_X1 U66 ( .A1(SUMB_23__16_), .A2(CARRYB_23__15_), .ZN(A2_38_) );
  XOR2_X1 U67 ( .A(CARRYB_23__15_), .B(SUMB_23__16_), .Z(A1_37_) );
  AND2_X1 U68 ( .A1(SUMB_23__15_), .A2(CARRYB_23__14_), .ZN(A2_37_) );
  XOR2_X1 U69 ( .A(CARRYB_23__14_), .B(SUMB_23__15_), .Z(A1_36_) );
  AND2_X1 U70 ( .A1(SUMB_23__14_), .A2(CARRYB_23__13_), .ZN(A2_36_) );
  XOR2_X1 U71 ( .A(CARRYB_23__13_), .B(SUMB_23__14_), .Z(A1_35_) );
  AND2_X1 U72 ( .A1(SUMB_23__13_), .A2(CARRYB_23__12_), .ZN(A2_35_) );
  XOR2_X1 U73 ( .A(CARRYB_23__12_), .B(SUMB_23__13_), .Z(A1_34_) );
  AND2_X1 U74 ( .A1(SUMB_23__12_), .A2(CARRYB_23__11_), .ZN(A2_34_) );
  XOR2_X1 U75 ( .A(CARRYB_23__11_), .B(SUMB_23__12_), .Z(A1_33_) );
  AND2_X1 U76 ( .A1(SUMB_23__11_), .A2(CARRYB_23__10_), .ZN(A2_33_) );
  XOR2_X1 U77 ( .A(CARRYB_23__10_), .B(SUMB_23__11_), .Z(A1_32_) );
  AND2_X1 U78 ( .A1(SUMB_23__10_), .A2(CARRYB_23__9_), .ZN(A2_32_) );
  XOR2_X1 U79 ( .A(CARRYB_23__9_), .B(SUMB_23__10_), .Z(A1_31_) );
  AND2_X1 U80 ( .A1(SUMB_23__9_), .A2(CARRYB_23__8_), .ZN(A2_31_) );
  XOR2_X1 U81 ( .A(CARRYB_23__8_), .B(SUMB_23__9_), .Z(A1_30_) );
  AND2_X1 U82 ( .A1(SUMB_23__8_), .A2(CARRYB_23__7_), .ZN(A2_30_) );
  XOR2_X1 U83 ( .A(CARRYB_23__7_), .B(SUMB_23__8_), .Z(A1_29_) );
  AND2_X1 U84 ( .A1(SUMB_23__7_), .A2(CARRYB_23__6_), .ZN(A2_29_) );
  XOR2_X1 U85 ( .A(CARRYB_23__6_), .B(SUMB_23__7_), .Z(A1_28_) );
  AND2_X1 U86 ( .A1(SUMB_23__6_), .A2(CARRYB_23__5_), .ZN(A2_28_) );
  XOR2_X1 U87 ( .A(CARRYB_23__5_), .B(SUMB_23__6_), .Z(A1_27_) );
  AND2_X1 U88 ( .A1(SUMB_23__5_), .A2(CARRYB_23__4_), .ZN(A2_27_) );
  XOR2_X1 U89 ( .A(CARRYB_23__4_), .B(SUMB_23__5_), .Z(A1_26_) );
  AND2_X1 U90 ( .A1(SUMB_23__4_), .A2(CARRYB_23__3_), .ZN(A2_26_) );
  XOR2_X1 U91 ( .A(CARRYB_23__3_), .B(SUMB_23__4_), .Z(A1_25_) );
  AND2_X1 U92 ( .A1(SUMB_23__3_), .A2(CARRYB_23__2_), .ZN(A2_25_) );
  XOR2_X1 U93 ( .A(CARRYB_23__2_), .B(SUMB_23__3_), .Z(A1_24_) );
  AND2_X1 U94 ( .A1(SUMB_23__2_), .A2(CARRYB_23__1_), .ZN(A2_24_) );
  XOR2_X1 U95 ( .A(CARRYB_23__1_), .B(SUMB_23__2_), .Z(A1_23_) );
  AND2_X1 U96 ( .A1(SUMB_23__1_), .A2(CARRYB_23__0_), .ZN(A2_23_) );
  XOR2_X1 U97 ( .A(CARRYB_23__0_), .B(SUMB_23__1_), .Z(A1_22_) );
  AND2_X1 U98 ( .A1(ab_1__22_), .A2(ab_0__23_), .ZN(CARRYB_1__22_) );
  XOR2_X1 U99 ( .A(ab_1__22_), .B(ab_0__23_), .Z(SUMB_1__22_) );
  AND2_X1 U100 ( .A1(ab_1__21_), .A2(ab_0__22_), .ZN(CARRYB_1__21_) );
  XOR2_X1 U101 ( .A(ab_1__21_), .B(ab_0__22_), .Z(SUMB_1__21_) );
  AND2_X1 U102 ( .A1(ab_1__20_), .A2(ab_0__21_), .ZN(CARRYB_1__20_) );
  XOR2_X1 U103 ( .A(ab_1__20_), .B(ab_0__21_), .Z(SUMB_1__20_) );
  AND2_X1 U104 ( .A1(ab_1__19_), .A2(ab_0__20_), .ZN(CARRYB_1__19_) );
  XOR2_X1 U105 ( .A(ab_1__19_), .B(ab_0__20_), .Z(SUMB_1__19_) );
  AND2_X1 U106 ( .A1(ab_1__18_), .A2(ab_0__19_), .ZN(CARRYB_1__18_) );
  XOR2_X1 U107 ( .A(ab_1__18_), .B(ab_0__19_), .Z(SUMB_1__18_) );
  AND2_X1 U108 ( .A1(ab_1__17_), .A2(ab_0__18_), .ZN(CARRYB_1__17_) );
  XOR2_X1 U109 ( .A(ab_1__17_), .B(ab_0__18_), .Z(SUMB_1__17_) );
  AND2_X1 U110 ( .A1(ab_1__16_), .A2(ab_0__17_), .ZN(CARRYB_1__16_) );
  XOR2_X1 U111 ( .A(ab_1__16_), .B(ab_0__17_), .Z(SUMB_1__16_) );
  AND2_X1 U112 ( .A1(ab_1__15_), .A2(ab_0__16_), .ZN(CARRYB_1__15_) );
  XOR2_X1 U113 ( .A(ab_1__15_), .B(ab_0__16_), .Z(SUMB_1__15_) );
  AND2_X1 U114 ( .A1(ab_1__14_), .A2(ab_0__15_), .ZN(CARRYB_1__14_) );
  XOR2_X1 U115 ( .A(ab_1__14_), .B(ab_0__15_), .Z(SUMB_1__14_) );
  AND2_X1 U116 ( .A1(ab_1__13_), .A2(ab_0__14_), .ZN(CARRYB_1__13_) );
  XOR2_X1 U117 ( .A(ab_1__13_), .B(ab_0__14_), .Z(SUMB_1__13_) );
  AND2_X1 U118 ( .A1(ab_1__12_), .A2(ab_0__13_), .ZN(CARRYB_1__12_) );
  XOR2_X1 U119 ( .A(ab_1__12_), .B(ab_0__13_), .Z(SUMB_1__12_) );
  AND2_X1 U120 ( .A1(ab_1__11_), .A2(ab_0__12_), .ZN(CARRYB_1__11_) );
  XOR2_X1 U121 ( .A(ab_1__11_), .B(ab_0__12_), .Z(SUMB_1__11_) );
  AND2_X1 U122 ( .A1(ab_1__10_), .A2(ab_0__11_), .ZN(CARRYB_1__10_) );
  XOR2_X1 U123 ( .A(ab_1__10_), .B(ab_0__11_), .Z(SUMB_1__10_) );
  AND2_X1 U124 ( .A1(ab_1__9_), .A2(ab_0__10_), .ZN(CARRYB_1__9_) );
  XOR2_X1 U125 ( .A(ab_1__9_), .B(ab_0__10_), .Z(SUMB_1__9_) );
  AND2_X1 U126 ( .A1(ab_1__8_), .A2(ab_0__9_), .ZN(CARRYB_1__8_) );
  XOR2_X1 U127 ( .A(ab_1__8_), .B(ab_0__9_), .Z(SUMB_1__8_) );
  AND2_X1 U128 ( .A1(ab_1__7_), .A2(ab_0__8_), .ZN(CARRYB_1__7_) );
  XOR2_X1 U129 ( .A(ab_1__7_), .B(ab_0__8_), .Z(SUMB_1__7_) );
  AND2_X1 U130 ( .A1(ab_1__6_), .A2(ab_0__7_), .ZN(CARRYB_1__6_) );
  XOR2_X1 U131 ( .A(ab_1__6_), .B(ab_0__7_), .Z(SUMB_1__6_) );
  AND2_X1 U132 ( .A1(ab_1__5_), .A2(ab_0__6_), .ZN(CARRYB_1__5_) );
  XOR2_X1 U133 ( .A(ab_1__5_), .B(ab_0__6_), .Z(SUMB_1__5_) );
  AND2_X1 U134 ( .A1(ab_1__4_), .A2(ab_0__5_), .ZN(CARRYB_1__4_) );
  XOR2_X1 U135 ( .A(ab_1__4_), .B(ab_0__5_), .Z(SUMB_1__4_) );
  AND2_X1 U136 ( .A1(ab_1__3_), .A2(ab_0__4_), .ZN(CARRYB_1__3_) );
  XOR2_X1 U137 ( .A(ab_1__3_), .B(ab_0__4_), .Z(SUMB_1__3_) );
  AND2_X1 U138 ( .A1(ab_1__2_), .A2(ab_0__3_), .ZN(CARRYB_1__2_) );
  XOR2_X1 U139 ( .A(ab_1__2_), .B(ab_0__3_), .Z(SUMB_1__2_) );
  AND2_X1 U140 ( .A1(ab_1__1_), .A2(ab_0__2_), .ZN(CARRYB_1__1_) );
  XOR2_X1 U141 ( .A(ab_1__1_), .B(ab_0__2_), .Z(SUMB_1__1_) );
  NOR2_X1 U142 ( .A1(n6), .A2(n7), .ZN(ab_9__9_) );
  NOR2_X1 U143 ( .A1(n6), .A2(n8), .ZN(ab_9__8_) );
  NOR2_X1 U144 ( .A1(n6), .A2(n9), .ZN(ab_9__7_) );
  NOR2_X1 U145 ( .A1(n6), .A2(n10), .ZN(ab_9__6_) );
  NOR2_X1 U146 ( .A1(n6), .A2(n11), .ZN(ab_9__5_) );
  NOR2_X1 U147 ( .A1(n6), .A2(n12), .ZN(ab_9__4_) );
  NOR2_X1 U148 ( .A1(n6), .A2(n13), .ZN(ab_9__3_) );
  NOR2_X1 U149 ( .A1(n6), .A2(n14), .ZN(ab_9__2_) );
  NOR2_X1 U150 ( .A1(A[9]), .A2(n1), .ZN(ab_9__23_) );
  NOR2_X1 U151 ( .A1(n6), .A2(n15), .ZN(ab_9__22_) );
  NOR2_X1 U152 ( .A1(n6), .A2(n16), .ZN(ab_9__21_) );
  NOR2_X1 U153 ( .A1(n6), .A2(n17), .ZN(ab_9__20_) );
  NOR2_X1 U154 ( .A1(n6), .A2(n18), .ZN(ab_9__1_) );
  NOR2_X1 U155 ( .A1(n6), .A2(n19), .ZN(ab_9__19_) );
  NOR2_X1 U156 ( .A1(n6), .A2(n20), .ZN(ab_9__18_) );
  NOR2_X1 U157 ( .A1(n6), .A2(n21), .ZN(ab_9__17_) );
  NOR2_X1 U158 ( .A1(n6), .A2(n22), .ZN(ab_9__16_) );
  NOR2_X1 U159 ( .A1(n6), .A2(n23), .ZN(ab_9__15_) );
  NOR2_X1 U160 ( .A1(n6), .A2(n24), .ZN(ab_9__14_) );
  NOR2_X1 U161 ( .A1(n6), .A2(n25), .ZN(ab_9__13_) );
  NOR2_X1 U162 ( .A1(n6), .A2(n26), .ZN(ab_9__12_) );
  NOR2_X1 U163 ( .A1(n6), .A2(n27), .ZN(ab_9__11_) );
  NOR2_X1 U164 ( .A1(n6), .A2(n28), .ZN(ab_9__10_) );
  NOR2_X1 U165 ( .A1(n6), .A2(n29), .ZN(ab_9__0_) );
  NOR2_X1 U166 ( .A1(n7), .A2(n30), .ZN(ab_8__9_) );
  NOR2_X1 U167 ( .A1(n8), .A2(n30), .ZN(ab_8__8_) );
  NOR2_X1 U168 ( .A1(n9), .A2(n30), .ZN(ab_8__7_) );
  NOR2_X1 U169 ( .A1(n10), .A2(n30), .ZN(ab_8__6_) );
  NOR2_X1 U170 ( .A1(n11), .A2(n30), .ZN(ab_8__5_) );
  NOR2_X1 U171 ( .A1(n12), .A2(n30), .ZN(ab_8__4_) );
  NOR2_X1 U172 ( .A1(n13), .A2(n30), .ZN(ab_8__3_) );
  NOR2_X1 U173 ( .A1(n14), .A2(n30), .ZN(ab_8__2_) );
  NOR2_X1 U174 ( .A1(A[8]), .A2(n1), .ZN(ab_8__23_) );
  NOR2_X1 U175 ( .A1(n15), .A2(n30), .ZN(ab_8__22_) );
  NOR2_X1 U176 ( .A1(n16), .A2(n30), .ZN(ab_8__21_) );
  NOR2_X1 U177 ( .A1(n17), .A2(n30), .ZN(ab_8__20_) );
  NOR2_X1 U178 ( .A1(n18), .A2(n30), .ZN(ab_8__1_) );
  NOR2_X1 U179 ( .A1(n19), .A2(n30), .ZN(ab_8__19_) );
  NOR2_X1 U180 ( .A1(n20), .A2(n30), .ZN(ab_8__18_) );
  NOR2_X1 U181 ( .A1(n21), .A2(n30), .ZN(ab_8__17_) );
  NOR2_X1 U182 ( .A1(n22), .A2(n30), .ZN(ab_8__16_) );
  NOR2_X1 U183 ( .A1(n23), .A2(n30), .ZN(ab_8__15_) );
  NOR2_X1 U184 ( .A1(n24), .A2(n30), .ZN(ab_8__14_) );
  NOR2_X1 U185 ( .A1(n25), .A2(n30), .ZN(ab_8__13_) );
  NOR2_X1 U186 ( .A1(n26), .A2(n30), .ZN(ab_8__12_) );
  NOR2_X1 U187 ( .A1(n27), .A2(n30), .ZN(ab_8__11_) );
  NOR2_X1 U188 ( .A1(n28), .A2(n30), .ZN(ab_8__10_) );
  NOR2_X1 U189 ( .A1(n29), .A2(n30), .ZN(ab_8__0_) );
  NOR2_X1 U190 ( .A1(n7), .A2(n31), .ZN(ab_7__9_) );
  NOR2_X1 U191 ( .A1(n8), .A2(n31), .ZN(ab_7__8_) );
  NOR2_X1 U192 ( .A1(n9), .A2(n31), .ZN(ab_7__7_) );
  NOR2_X1 U193 ( .A1(n10), .A2(n31), .ZN(ab_7__6_) );
  NOR2_X1 U194 ( .A1(n11), .A2(n31), .ZN(ab_7__5_) );
  NOR2_X1 U195 ( .A1(n12), .A2(n31), .ZN(ab_7__4_) );
  NOR2_X1 U196 ( .A1(n13), .A2(n31), .ZN(ab_7__3_) );
  NOR2_X1 U197 ( .A1(n14), .A2(n31), .ZN(ab_7__2_) );
  NOR2_X1 U198 ( .A1(A[7]), .A2(n1), .ZN(ab_7__23_) );
  NOR2_X1 U199 ( .A1(n15), .A2(n31), .ZN(ab_7__22_) );
  NOR2_X1 U200 ( .A1(n16), .A2(n31), .ZN(ab_7__21_) );
  NOR2_X1 U201 ( .A1(n17), .A2(n31), .ZN(ab_7__20_) );
  NOR2_X1 U202 ( .A1(n18), .A2(n31), .ZN(ab_7__1_) );
  NOR2_X1 U203 ( .A1(n19), .A2(n31), .ZN(ab_7__19_) );
  NOR2_X1 U204 ( .A1(n20), .A2(n31), .ZN(ab_7__18_) );
  NOR2_X1 U205 ( .A1(n21), .A2(n31), .ZN(ab_7__17_) );
  NOR2_X1 U206 ( .A1(n22), .A2(n31), .ZN(ab_7__16_) );
  NOR2_X1 U207 ( .A1(n23), .A2(n31), .ZN(ab_7__15_) );
  NOR2_X1 U208 ( .A1(n24), .A2(n31), .ZN(ab_7__14_) );
  NOR2_X1 U209 ( .A1(n25), .A2(n31), .ZN(ab_7__13_) );
  NOR2_X1 U210 ( .A1(n26), .A2(n31), .ZN(ab_7__12_) );
  NOR2_X1 U211 ( .A1(n27), .A2(n31), .ZN(ab_7__11_) );
  NOR2_X1 U212 ( .A1(n28), .A2(n31), .ZN(ab_7__10_) );
  NOR2_X1 U213 ( .A1(n29), .A2(n31), .ZN(ab_7__0_) );
  NOR2_X1 U214 ( .A1(n7), .A2(n32), .ZN(ab_6__9_) );
  NOR2_X1 U215 ( .A1(n8), .A2(n32), .ZN(ab_6__8_) );
  NOR2_X1 U216 ( .A1(n9), .A2(n32), .ZN(ab_6__7_) );
  NOR2_X1 U217 ( .A1(n10), .A2(n32), .ZN(ab_6__6_) );
  NOR2_X1 U218 ( .A1(n11), .A2(n32), .ZN(ab_6__5_) );
  NOR2_X1 U219 ( .A1(n12), .A2(n32), .ZN(ab_6__4_) );
  NOR2_X1 U220 ( .A1(n13), .A2(n32), .ZN(ab_6__3_) );
  NOR2_X1 U221 ( .A1(n14), .A2(n32), .ZN(ab_6__2_) );
  NOR2_X1 U222 ( .A1(A[6]), .A2(n1), .ZN(ab_6__23_) );
  NOR2_X1 U223 ( .A1(n15), .A2(n32), .ZN(ab_6__22_) );
  NOR2_X1 U224 ( .A1(n16), .A2(n32), .ZN(ab_6__21_) );
  NOR2_X1 U225 ( .A1(n17), .A2(n32), .ZN(ab_6__20_) );
  NOR2_X1 U226 ( .A1(n18), .A2(n32), .ZN(ab_6__1_) );
  NOR2_X1 U227 ( .A1(n19), .A2(n32), .ZN(ab_6__19_) );
  NOR2_X1 U228 ( .A1(n20), .A2(n32), .ZN(ab_6__18_) );
  NOR2_X1 U229 ( .A1(n21), .A2(n32), .ZN(ab_6__17_) );
  NOR2_X1 U230 ( .A1(n22), .A2(n32), .ZN(ab_6__16_) );
  NOR2_X1 U231 ( .A1(n23), .A2(n32), .ZN(ab_6__15_) );
  NOR2_X1 U232 ( .A1(n24), .A2(n32), .ZN(ab_6__14_) );
  NOR2_X1 U233 ( .A1(n25), .A2(n32), .ZN(ab_6__13_) );
  NOR2_X1 U234 ( .A1(n26), .A2(n32), .ZN(ab_6__12_) );
  NOR2_X1 U235 ( .A1(n27), .A2(n32), .ZN(ab_6__11_) );
  NOR2_X1 U236 ( .A1(n28), .A2(n32), .ZN(ab_6__10_) );
  NOR2_X1 U237 ( .A1(n29), .A2(n32), .ZN(ab_6__0_) );
  NOR2_X1 U238 ( .A1(n7), .A2(n33), .ZN(ab_5__9_) );
  NOR2_X1 U239 ( .A1(n8), .A2(n33), .ZN(ab_5__8_) );
  NOR2_X1 U240 ( .A1(n9), .A2(n33), .ZN(ab_5__7_) );
  NOR2_X1 U241 ( .A1(n10), .A2(n33), .ZN(ab_5__6_) );
  NOR2_X1 U242 ( .A1(n11), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U243 ( .A1(n12), .A2(n33), .ZN(ab_5__4_) );
  NOR2_X1 U244 ( .A1(n13), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U245 ( .A1(n14), .A2(n33), .ZN(ab_5__2_) );
  NOR2_X1 U246 ( .A1(A[5]), .A2(n1), .ZN(ab_5__23_) );
  NOR2_X1 U247 ( .A1(n15), .A2(n33), .ZN(ab_5__22_) );
  NOR2_X1 U248 ( .A1(n16), .A2(n33), .ZN(ab_5__21_) );
  NOR2_X1 U249 ( .A1(n17), .A2(n33), .ZN(ab_5__20_) );
  NOR2_X1 U250 ( .A1(n18), .A2(n33), .ZN(ab_5__1_) );
  NOR2_X1 U251 ( .A1(n19), .A2(n33), .ZN(ab_5__19_) );
  NOR2_X1 U252 ( .A1(n20), .A2(n33), .ZN(ab_5__18_) );
  NOR2_X1 U253 ( .A1(n21), .A2(n33), .ZN(ab_5__17_) );
  NOR2_X1 U254 ( .A1(n22), .A2(n33), .ZN(ab_5__16_) );
  NOR2_X1 U255 ( .A1(n23), .A2(n33), .ZN(ab_5__15_) );
  NOR2_X1 U256 ( .A1(n24), .A2(n33), .ZN(ab_5__14_) );
  NOR2_X1 U257 ( .A1(n25), .A2(n33), .ZN(ab_5__13_) );
  NOR2_X1 U258 ( .A1(n26), .A2(n33), .ZN(ab_5__12_) );
  NOR2_X1 U259 ( .A1(n27), .A2(n33), .ZN(ab_5__11_) );
  NOR2_X1 U260 ( .A1(n28), .A2(n33), .ZN(ab_5__10_) );
  NOR2_X1 U261 ( .A1(n29), .A2(n33), .ZN(ab_5__0_) );
  NOR2_X1 U262 ( .A1(n7), .A2(n34), .ZN(ab_4__9_) );
  NOR2_X1 U263 ( .A1(n8), .A2(n34), .ZN(ab_4__8_) );
  NOR2_X1 U264 ( .A1(n9), .A2(n34), .ZN(ab_4__7_) );
  NOR2_X1 U265 ( .A1(n10), .A2(n34), .ZN(ab_4__6_) );
  NOR2_X1 U266 ( .A1(n11), .A2(n34), .ZN(ab_4__5_) );
  NOR2_X1 U267 ( .A1(n12), .A2(n34), .ZN(ab_4__4_) );
  NOR2_X1 U268 ( .A1(n13), .A2(n34), .ZN(ab_4__3_) );
  NOR2_X1 U269 ( .A1(n14), .A2(n34), .ZN(ab_4__2_) );
  NOR2_X1 U270 ( .A1(A[4]), .A2(n1), .ZN(ab_4__23_) );
  NOR2_X1 U271 ( .A1(n15), .A2(n34), .ZN(ab_4__22_) );
  NOR2_X1 U272 ( .A1(n16), .A2(n34), .ZN(ab_4__21_) );
  NOR2_X1 U273 ( .A1(n17), .A2(n34), .ZN(ab_4__20_) );
  NOR2_X1 U274 ( .A1(n18), .A2(n34), .ZN(ab_4__1_) );
  NOR2_X1 U275 ( .A1(n19), .A2(n34), .ZN(ab_4__19_) );
  NOR2_X1 U276 ( .A1(n20), .A2(n34), .ZN(ab_4__18_) );
  NOR2_X1 U277 ( .A1(n21), .A2(n34), .ZN(ab_4__17_) );
  NOR2_X1 U278 ( .A1(n22), .A2(n34), .ZN(ab_4__16_) );
  NOR2_X1 U279 ( .A1(n23), .A2(n34), .ZN(ab_4__15_) );
  NOR2_X1 U280 ( .A1(n24), .A2(n34), .ZN(ab_4__14_) );
  NOR2_X1 U281 ( .A1(n25), .A2(n34), .ZN(ab_4__13_) );
  NOR2_X1 U282 ( .A1(n26), .A2(n34), .ZN(ab_4__12_) );
  NOR2_X1 U283 ( .A1(n27), .A2(n34), .ZN(ab_4__11_) );
  NOR2_X1 U284 ( .A1(n28), .A2(n34), .ZN(ab_4__10_) );
  NOR2_X1 U285 ( .A1(n29), .A2(n34), .ZN(ab_4__0_) );
  NOR2_X1 U286 ( .A1(n7), .A2(n35), .ZN(ab_3__9_) );
  NOR2_X1 U287 ( .A1(n8), .A2(n35), .ZN(ab_3__8_) );
  NOR2_X1 U288 ( .A1(n9), .A2(n35), .ZN(ab_3__7_) );
  NOR2_X1 U289 ( .A1(n10), .A2(n35), .ZN(ab_3__6_) );
  NOR2_X1 U290 ( .A1(n11), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U291 ( .A1(n12), .A2(n35), .ZN(ab_3__4_) );
  NOR2_X1 U292 ( .A1(n13), .A2(n35), .ZN(ab_3__3_) );
  NOR2_X1 U293 ( .A1(n14), .A2(n35), .ZN(ab_3__2_) );
  NOR2_X1 U294 ( .A1(A[3]), .A2(n1), .ZN(ab_3__23_) );
  NOR2_X1 U295 ( .A1(n15), .A2(n35), .ZN(ab_3__22_) );
  NOR2_X1 U296 ( .A1(n16), .A2(n35), .ZN(ab_3__21_) );
  NOR2_X1 U297 ( .A1(n17), .A2(n35), .ZN(ab_3__20_) );
  NOR2_X1 U298 ( .A1(n18), .A2(n35), .ZN(ab_3__1_) );
  NOR2_X1 U299 ( .A1(n19), .A2(n35), .ZN(ab_3__19_) );
  NOR2_X1 U300 ( .A1(n20), .A2(n35), .ZN(ab_3__18_) );
  NOR2_X1 U301 ( .A1(n21), .A2(n35), .ZN(ab_3__17_) );
  NOR2_X1 U302 ( .A1(n22), .A2(n35), .ZN(ab_3__16_) );
  NOR2_X1 U303 ( .A1(n23), .A2(n35), .ZN(ab_3__15_) );
  NOR2_X1 U304 ( .A1(n24), .A2(n35), .ZN(ab_3__14_) );
  NOR2_X1 U305 ( .A1(n25), .A2(n35), .ZN(ab_3__13_) );
  NOR2_X1 U306 ( .A1(n26), .A2(n35), .ZN(ab_3__12_) );
  NOR2_X1 U307 ( .A1(n27), .A2(n35), .ZN(ab_3__11_) );
  NOR2_X1 U308 ( .A1(n28), .A2(n35), .ZN(ab_3__10_) );
  NOR2_X1 U309 ( .A1(n29), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U310 ( .A1(n7), .A2(n36), .ZN(ab_2__9_) );
  NOR2_X1 U311 ( .A1(n8), .A2(n36), .ZN(ab_2__8_) );
  NOR2_X1 U312 ( .A1(n9), .A2(n36), .ZN(ab_2__7_) );
  NOR2_X1 U313 ( .A1(n10), .A2(n36), .ZN(ab_2__6_) );
  NOR2_X1 U314 ( .A1(n11), .A2(n36), .ZN(ab_2__5_) );
  NOR2_X1 U315 ( .A1(n12), .A2(n36), .ZN(ab_2__4_) );
  NOR2_X1 U316 ( .A1(n13), .A2(n36), .ZN(ab_2__3_) );
  NOR2_X1 U317 ( .A1(n14), .A2(n36), .ZN(ab_2__2_) );
  NOR2_X1 U318 ( .A1(A[2]), .A2(n1), .ZN(ab_2__23_) );
  NOR2_X1 U319 ( .A1(n15), .A2(n36), .ZN(ab_2__22_) );
  NOR2_X1 U320 ( .A1(n16), .A2(n36), .ZN(ab_2__21_) );
  NOR2_X1 U321 ( .A1(n17), .A2(n36), .ZN(ab_2__20_) );
  NOR2_X1 U322 ( .A1(n18), .A2(n36), .ZN(ab_2__1_) );
  NOR2_X1 U323 ( .A1(n19), .A2(n36), .ZN(ab_2__19_) );
  NOR2_X1 U324 ( .A1(n20), .A2(n36), .ZN(ab_2__18_) );
  NOR2_X1 U325 ( .A1(n21), .A2(n36), .ZN(ab_2__17_) );
  NOR2_X1 U326 ( .A1(n22), .A2(n36), .ZN(ab_2__16_) );
  NOR2_X1 U327 ( .A1(n23), .A2(n36), .ZN(ab_2__15_) );
  NOR2_X1 U328 ( .A1(n24), .A2(n36), .ZN(ab_2__14_) );
  NOR2_X1 U329 ( .A1(n25), .A2(n36), .ZN(ab_2__13_) );
  NOR2_X1 U330 ( .A1(n26), .A2(n36), .ZN(ab_2__12_) );
  NOR2_X1 U331 ( .A1(n27), .A2(n36), .ZN(ab_2__11_) );
  NOR2_X1 U332 ( .A1(n28), .A2(n36), .ZN(ab_2__10_) );
  NOR2_X1 U333 ( .A1(n29), .A2(n36), .ZN(ab_2__0_) );
  NOR2_X1 U334 ( .A1(B[9]), .A2(n4), .ZN(ab_23__9_) );
  NOR2_X1 U335 ( .A1(B[8]), .A2(n4), .ZN(ab_23__8_) );
  NOR2_X1 U336 ( .A1(B[7]), .A2(n4), .ZN(ab_23__7_) );
  NOR2_X1 U337 ( .A1(B[6]), .A2(n4), .ZN(ab_23__6_) );
  NOR2_X1 U338 ( .A1(B[5]), .A2(n3), .ZN(ab_23__5_) );
  NOR2_X1 U339 ( .A1(B[4]), .A2(n3), .ZN(ab_23__4_) );
  NOR2_X1 U340 ( .A1(B[3]), .A2(n3), .ZN(ab_23__3_) );
  NOR2_X1 U341 ( .A1(B[2]), .A2(n3), .ZN(ab_23__2_) );
  NOR2_X1 U342 ( .A1(n1), .A2(n3), .ZN(ab_23__23_) );
  NOR2_X1 U343 ( .A1(B[22]), .A2(n3), .ZN(ab_23__22_) );
  NOR2_X1 U344 ( .A1(B[21]), .A2(n3), .ZN(ab_23__21_) );
  NOR2_X1 U345 ( .A1(B[20]), .A2(n3), .ZN(ab_23__20_) );
  NOR2_X1 U346 ( .A1(B[1]), .A2(n3), .ZN(ab_23__1_) );
  NOR2_X1 U347 ( .A1(B[19]), .A2(n3), .ZN(ab_23__19_) );
  NOR2_X1 U348 ( .A1(B[18]), .A2(n3), .ZN(ab_23__18_) );
  NOR2_X1 U349 ( .A1(B[17]), .A2(n3), .ZN(ab_23__17_) );
  NOR2_X1 U350 ( .A1(B[16]), .A2(n3), .ZN(ab_23__16_) );
  NOR2_X1 U351 ( .A1(B[15]), .A2(n3), .ZN(ab_23__15_) );
  NOR2_X1 U352 ( .A1(B[14]), .A2(n3), .ZN(ab_23__14_) );
  NOR2_X1 U353 ( .A1(B[13]), .A2(n3), .ZN(ab_23__13_) );
  NOR2_X1 U354 ( .A1(B[12]), .A2(n3), .ZN(ab_23__12_) );
  NOR2_X1 U355 ( .A1(B[11]), .A2(n3), .ZN(ab_23__11_) );
  NOR2_X1 U356 ( .A1(B[10]), .A2(n3), .ZN(ab_23__10_) );
  NOR2_X1 U357 ( .A1(B[0]), .A2(n3), .ZN(ab_23__0_) );
  NOR2_X1 U358 ( .A1(n7), .A2(n37), .ZN(ab_22__9_) );
  NOR2_X1 U359 ( .A1(n8), .A2(n37), .ZN(ab_22__8_) );
  NOR2_X1 U360 ( .A1(n9), .A2(n37), .ZN(ab_22__7_) );
  NOR2_X1 U361 ( .A1(n10), .A2(n37), .ZN(ab_22__6_) );
  NOR2_X1 U362 ( .A1(n11), .A2(n37), .ZN(ab_22__5_) );
  NOR2_X1 U363 ( .A1(n12), .A2(n37), .ZN(ab_22__4_) );
  NOR2_X1 U364 ( .A1(n13), .A2(n37), .ZN(ab_22__3_) );
  NOR2_X1 U365 ( .A1(n14), .A2(n37), .ZN(ab_22__2_) );
  NOR2_X1 U366 ( .A1(A[22]), .A2(n1), .ZN(ab_22__23_) );
  NOR2_X1 U367 ( .A1(n15), .A2(n37), .ZN(ab_22__22_) );
  NOR2_X1 U368 ( .A1(n16), .A2(n37), .ZN(ab_22__21_) );
  NOR2_X1 U369 ( .A1(n17), .A2(n37), .ZN(ab_22__20_) );
  NOR2_X1 U370 ( .A1(n18), .A2(n37), .ZN(ab_22__1_) );
  NOR2_X1 U371 ( .A1(n19), .A2(n37), .ZN(ab_22__19_) );
  NOR2_X1 U372 ( .A1(n20), .A2(n37), .ZN(ab_22__18_) );
  NOR2_X1 U373 ( .A1(n21), .A2(n37), .ZN(ab_22__17_) );
  NOR2_X1 U374 ( .A1(n22), .A2(n37), .ZN(ab_22__16_) );
  NOR2_X1 U375 ( .A1(n23), .A2(n37), .ZN(ab_22__15_) );
  NOR2_X1 U376 ( .A1(n24), .A2(n37), .ZN(ab_22__14_) );
  NOR2_X1 U377 ( .A1(n25), .A2(n37), .ZN(ab_22__13_) );
  NOR2_X1 U378 ( .A1(n26), .A2(n37), .ZN(ab_22__12_) );
  NOR2_X1 U379 ( .A1(n27), .A2(n37), .ZN(ab_22__11_) );
  NOR2_X1 U380 ( .A1(n28), .A2(n37), .ZN(ab_22__10_) );
  NOR2_X1 U381 ( .A1(n29), .A2(n37), .ZN(ab_22__0_) );
  NOR2_X1 U382 ( .A1(n7), .A2(n38), .ZN(ab_21__9_) );
  NOR2_X1 U383 ( .A1(n8), .A2(n38), .ZN(ab_21__8_) );
  NOR2_X1 U384 ( .A1(n9), .A2(n38), .ZN(ab_21__7_) );
  NOR2_X1 U385 ( .A1(n10), .A2(n38), .ZN(ab_21__6_) );
  NOR2_X1 U386 ( .A1(n11), .A2(n38), .ZN(ab_21__5_) );
  NOR2_X1 U387 ( .A1(n12), .A2(n38), .ZN(ab_21__4_) );
  NOR2_X1 U388 ( .A1(n13), .A2(n38), .ZN(ab_21__3_) );
  NOR2_X1 U389 ( .A1(n14), .A2(n38), .ZN(ab_21__2_) );
  NOR2_X1 U390 ( .A1(A[21]), .A2(n1), .ZN(ab_21__23_) );
  NOR2_X1 U391 ( .A1(n15), .A2(n38), .ZN(ab_21__22_) );
  NOR2_X1 U392 ( .A1(n16), .A2(n38), .ZN(ab_21__21_) );
  NOR2_X1 U393 ( .A1(n17), .A2(n38), .ZN(ab_21__20_) );
  NOR2_X1 U394 ( .A1(n18), .A2(n38), .ZN(ab_21__1_) );
  NOR2_X1 U395 ( .A1(n19), .A2(n38), .ZN(ab_21__19_) );
  NOR2_X1 U396 ( .A1(n20), .A2(n38), .ZN(ab_21__18_) );
  NOR2_X1 U397 ( .A1(n21), .A2(n38), .ZN(ab_21__17_) );
  NOR2_X1 U398 ( .A1(n22), .A2(n38), .ZN(ab_21__16_) );
  NOR2_X1 U399 ( .A1(n23), .A2(n38), .ZN(ab_21__15_) );
  NOR2_X1 U400 ( .A1(n24), .A2(n38), .ZN(ab_21__14_) );
  NOR2_X1 U401 ( .A1(n25), .A2(n38), .ZN(ab_21__13_) );
  NOR2_X1 U402 ( .A1(n26), .A2(n38), .ZN(ab_21__12_) );
  NOR2_X1 U403 ( .A1(n27), .A2(n38), .ZN(ab_21__11_) );
  NOR2_X1 U404 ( .A1(n28), .A2(n38), .ZN(ab_21__10_) );
  NOR2_X1 U405 ( .A1(n29), .A2(n38), .ZN(ab_21__0_) );
  NOR2_X1 U406 ( .A1(n7), .A2(n39), .ZN(ab_20__9_) );
  NOR2_X1 U407 ( .A1(n8), .A2(n39), .ZN(ab_20__8_) );
  NOR2_X1 U408 ( .A1(n9), .A2(n39), .ZN(ab_20__7_) );
  NOR2_X1 U409 ( .A1(n10), .A2(n39), .ZN(ab_20__6_) );
  NOR2_X1 U410 ( .A1(n11), .A2(n39), .ZN(ab_20__5_) );
  NOR2_X1 U411 ( .A1(n12), .A2(n39), .ZN(ab_20__4_) );
  NOR2_X1 U412 ( .A1(n13), .A2(n39), .ZN(ab_20__3_) );
  NOR2_X1 U413 ( .A1(n14), .A2(n39), .ZN(ab_20__2_) );
  NOR2_X1 U414 ( .A1(A[20]), .A2(n1), .ZN(ab_20__23_) );
  NOR2_X1 U415 ( .A1(n15), .A2(n39), .ZN(ab_20__22_) );
  NOR2_X1 U416 ( .A1(n16), .A2(n39), .ZN(ab_20__21_) );
  NOR2_X1 U417 ( .A1(n17), .A2(n39), .ZN(ab_20__20_) );
  NOR2_X1 U418 ( .A1(n18), .A2(n39), .ZN(ab_20__1_) );
  NOR2_X1 U419 ( .A1(n19), .A2(n39), .ZN(ab_20__19_) );
  NOR2_X1 U420 ( .A1(n20), .A2(n39), .ZN(ab_20__18_) );
  NOR2_X1 U421 ( .A1(n21), .A2(n39), .ZN(ab_20__17_) );
  NOR2_X1 U422 ( .A1(n22), .A2(n39), .ZN(ab_20__16_) );
  NOR2_X1 U423 ( .A1(n23), .A2(n39), .ZN(ab_20__15_) );
  NOR2_X1 U424 ( .A1(n24), .A2(n39), .ZN(ab_20__14_) );
  NOR2_X1 U425 ( .A1(n25), .A2(n39), .ZN(ab_20__13_) );
  NOR2_X1 U426 ( .A1(n26), .A2(n39), .ZN(ab_20__12_) );
  NOR2_X1 U427 ( .A1(n27), .A2(n39), .ZN(ab_20__11_) );
  NOR2_X1 U428 ( .A1(n28), .A2(n39), .ZN(ab_20__10_) );
  NOR2_X1 U429 ( .A1(n29), .A2(n39), .ZN(ab_20__0_) );
  NOR2_X1 U430 ( .A1(n7), .A2(n40), .ZN(ab_1__9_) );
  NOR2_X1 U431 ( .A1(n8), .A2(n40), .ZN(ab_1__8_) );
  NOR2_X1 U432 ( .A1(n9), .A2(n40), .ZN(ab_1__7_) );
  NOR2_X1 U433 ( .A1(n10), .A2(n40), .ZN(ab_1__6_) );
  NOR2_X1 U434 ( .A1(n11), .A2(n40), .ZN(ab_1__5_) );
  NOR2_X1 U435 ( .A1(n12), .A2(n40), .ZN(ab_1__4_) );
  NOR2_X1 U436 ( .A1(n13), .A2(n40), .ZN(ab_1__3_) );
  NOR2_X1 U437 ( .A1(n14), .A2(n40), .ZN(ab_1__2_) );
  NOR2_X1 U438 ( .A1(A[1]), .A2(n1), .ZN(ab_1__23_) );
  NOR2_X1 U439 ( .A1(n15), .A2(n40), .ZN(ab_1__22_) );
  NOR2_X1 U440 ( .A1(n16), .A2(n40), .ZN(ab_1__21_) );
  NOR2_X1 U441 ( .A1(n17), .A2(n40), .ZN(ab_1__20_) );
  NOR2_X1 U442 ( .A1(n19), .A2(n40), .ZN(ab_1__19_) );
  NOR2_X1 U443 ( .A1(n20), .A2(n40), .ZN(ab_1__18_) );
  NOR2_X1 U444 ( .A1(n21), .A2(n40), .ZN(ab_1__17_) );
  NOR2_X1 U445 ( .A1(n22), .A2(n40), .ZN(ab_1__16_) );
  NOR2_X1 U446 ( .A1(n23), .A2(n40), .ZN(ab_1__15_) );
  NOR2_X1 U447 ( .A1(n24), .A2(n40), .ZN(ab_1__14_) );
  NOR2_X1 U448 ( .A1(n25), .A2(n40), .ZN(ab_1__13_) );
  NOR2_X1 U449 ( .A1(n26), .A2(n40), .ZN(ab_1__12_) );
  NOR2_X1 U450 ( .A1(n27), .A2(n40), .ZN(ab_1__11_) );
  NOR2_X1 U451 ( .A1(n28), .A2(n40), .ZN(ab_1__10_) );
  NOR2_X1 U452 ( .A1(n7), .A2(n41), .ZN(ab_19__9_) );
  NOR2_X1 U453 ( .A1(n8), .A2(n41), .ZN(ab_19__8_) );
  NOR2_X1 U454 ( .A1(n9), .A2(n41), .ZN(ab_19__7_) );
  NOR2_X1 U455 ( .A1(n10), .A2(n41), .ZN(ab_19__6_) );
  NOR2_X1 U456 ( .A1(n11), .A2(n41), .ZN(ab_19__5_) );
  NOR2_X1 U457 ( .A1(n12), .A2(n41), .ZN(ab_19__4_) );
  NOR2_X1 U458 ( .A1(n13), .A2(n41), .ZN(ab_19__3_) );
  NOR2_X1 U459 ( .A1(n14), .A2(n41), .ZN(ab_19__2_) );
  NOR2_X1 U460 ( .A1(A[19]), .A2(n1), .ZN(ab_19__23_) );
  NOR2_X1 U461 ( .A1(n15), .A2(n41), .ZN(ab_19__22_) );
  NOR2_X1 U462 ( .A1(n16), .A2(n41), .ZN(ab_19__21_) );
  NOR2_X1 U463 ( .A1(n17), .A2(n41), .ZN(ab_19__20_) );
  NOR2_X1 U464 ( .A1(n18), .A2(n41), .ZN(ab_19__1_) );
  NOR2_X1 U465 ( .A1(n19), .A2(n41), .ZN(ab_19__19_) );
  NOR2_X1 U466 ( .A1(n20), .A2(n41), .ZN(ab_19__18_) );
  NOR2_X1 U467 ( .A1(n21), .A2(n41), .ZN(ab_19__17_) );
  NOR2_X1 U468 ( .A1(n22), .A2(n41), .ZN(ab_19__16_) );
  NOR2_X1 U469 ( .A1(n23), .A2(n41), .ZN(ab_19__15_) );
  NOR2_X1 U470 ( .A1(n24), .A2(n41), .ZN(ab_19__14_) );
  NOR2_X1 U471 ( .A1(n25), .A2(n41), .ZN(ab_19__13_) );
  NOR2_X1 U472 ( .A1(n26), .A2(n41), .ZN(ab_19__12_) );
  NOR2_X1 U473 ( .A1(n27), .A2(n41), .ZN(ab_19__11_) );
  NOR2_X1 U474 ( .A1(n28), .A2(n41), .ZN(ab_19__10_) );
  NOR2_X1 U475 ( .A1(n29), .A2(n41), .ZN(ab_19__0_) );
  NOR2_X1 U476 ( .A1(n7), .A2(n42), .ZN(ab_18__9_) );
  NOR2_X1 U477 ( .A1(n8), .A2(n42), .ZN(ab_18__8_) );
  NOR2_X1 U478 ( .A1(n9), .A2(n42), .ZN(ab_18__7_) );
  NOR2_X1 U479 ( .A1(n10), .A2(n42), .ZN(ab_18__6_) );
  NOR2_X1 U480 ( .A1(n11), .A2(n42), .ZN(ab_18__5_) );
  NOR2_X1 U481 ( .A1(n12), .A2(n42), .ZN(ab_18__4_) );
  NOR2_X1 U482 ( .A1(n13), .A2(n42), .ZN(ab_18__3_) );
  NOR2_X1 U483 ( .A1(n14), .A2(n42), .ZN(ab_18__2_) );
  NOR2_X1 U484 ( .A1(A[18]), .A2(n1), .ZN(ab_18__23_) );
  NOR2_X1 U485 ( .A1(n15), .A2(n42), .ZN(ab_18__22_) );
  NOR2_X1 U486 ( .A1(n16), .A2(n42), .ZN(ab_18__21_) );
  NOR2_X1 U487 ( .A1(n17), .A2(n42), .ZN(ab_18__20_) );
  NOR2_X1 U488 ( .A1(n18), .A2(n42), .ZN(ab_18__1_) );
  NOR2_X1 U489 ( .A1(n19), .A2(n42), .ZN(ab_18__19_) );
  NOR2_X1 U490 ( .A1(n20), .A2(n42), .ZN(ab_18__18_) );
  NOR2_X1 U491 ( .A1(n21), .A2(n42), .ZN(ab_18__17_) );
  NOR2_X1 U492 ( .A1(n22), .A2(n42), .ZN(ab_18__16_) );
  NOR2_X1 U493 ( .A1(n23), .A2(n42), .ZN(ab_18__15_) );
  NOR2_X1 U494 ( .A1(n24), .A2(n42), .ZN(ab_18__14_) );
  NOR2_X1 U495 ( .A1(n25), .A2(n42), .ZN(ab_18__13_) );
  NOR2_X1 U496 ( .A1(n26), .A2(n42), .ZN(ab_18__12_) );
  NOR2_X1 U497 ( .A1(n27), .A2(n42), .ZN(ab_18__11_) );
  NOR2_X1 U498 ( .A1(n28), .A2(n42), .ZN(ab_18__10_) );
  NOR2_X1 U499 ( .A1(n29), .A2(n42), .ZN(ab_18__0_) );
  NOR2_X1 U500 ( .A1(n7), .A2(n43), .ZN(ab_17__9_) );
  NOR2_X1 U501 ( .A1(n8), .A2(n43), .ZN(ab_17__8_) );
  NOR2_X1 U502 ( .A1(n9), .A2(n43), .ZN(ab_17__7_) );
  NOR2_X1 U503 ( .A1(n10), .A2(n43), .ZN(ab_17__6_) );
  NOR2_X1 U504 ( .A1(n11), .A2(n43), .ZN(ab_17__5_) );
  NOR2_X1 U505 ( .A1(n12), .A2(n43), .ZN(ab_17__4_) );
  NOR2_X1 U506 ( .A1(n13), .A2(n43), .ZN(ab_17__3_) );
  NOR2_X1 U507 ( .A1(n14), .A2(n43), .ZN(ab_17__2_) );
  NOR2_X1 U508 ( .A1(A[17]), .A2(n1), .ZN(ab_17__23_) );
  NOR2_X1 U509 ( .A1(n15), .A2(n43), .ZN(ab_17__22_) );
  NOR2_X1 U510 ( .A1(n16), .A2(n43), .ZN(ab_17__21_) );
  NOR2_X1 U511 ( .A1(n17), .A2(n43), .ZN(ab_17__20_) );
  NOR2_X1 U512 ( .A1(n18), .A2(n43), .ZN(ab_17__1_) );
  NOR2_X1 U513 ( .A1(n19), .A2(n43), .ZN(ab_17__19_) );
  NOR2_X1 U514 ( .A1(n20), .A2(n43), .ZN(ab_17__18_) );
  NOR2_X1 U515 ( .A1(n21), .A2(n43), .ZN(ab_17__17_) );
  NOR2_X1 U516 ( .A1(n22), .A2(n43), .ZN(ab_17__16_) );
  NOR2_X1 U517 ( .A1(n23), .A2(n43), .ZN(ab_17__15_) );
  NOR2_X1 U518 ( .A1(n24), .A2(n43), .ZN(ab_17__14_) );
  NOR2_X1 U519 ( .A1(n25), .A2(n43), .ZN(ab_17__13_) );
  NOR2_X1 U520 ( .A1(n26), .A2(n43), .ZN(ab_17__12_) );
  NOR2_X1 U521 ( .A1(n27), .A2(n43), .ZN(ab_17__11_) );
  NOR2_X1 U522 ( .A1(n28), .A2(n43), .ZN(ab_17__10_) );
  NOR2_X1 U523 ( .A1(n29), .A2(n43), .ZN(ab_17__0_) );
  NOR2_X1 U524 ( .A1(n7), .A2(n44), .ZN(ab_16__9_) );
  NOR2_X1 U525 ( .A1(n8), .A2(n44), .ZN(ab_16__8_) );
  NOR2_X1 U526 ( .A1(n9), .A2(n44), .ZN(ab_16__7_) );
  NOR2_X1 U527 ( .A1(n10), .A2(n44), .ZN(ab_16__6_) );
  NOR2_X1 U528 ( .A1(n11), .A2(n44), .ZN(ab_16__5_) );
  NOR2_X1 U529 ( .A1(n12), .A2(n44), .ZN(ab_16__4_) );
  NOR2_X1 U530 ( .A1(n13), .A2(n44), .ZN(ab_16__3_) );
  NOR2_X1 U531 ( .A1(n14), .A2(n44), .ZN(ab_16__2_) );
  NOR2_X1 U532 ( .A1(A[16]), .A2(n1), .ZN(ab_16__23_) );
  NOR2_X1 U533 ( .A1(n15), .A2(n44), .ZN(ab_16__22_) );
  NOR2_X1 U534 ( .A1(n16), .A2(n44), .ZN(ab_16__21_) );
  NOR2_X1 U535 ( .A1(n17), .A2(n44), .ZN(ab_16__20_) );
  NOR2_X1 U536 ( .A1(n18), .A2(n44), .ZN(ab_16__1_) );
  NOR2_X1 U537 ( .A1(n19), .A2(n44), .ZN(ab_16__19_) );
  NOR2_X1 U538 ( .A1(n20), .A2(n44), .ZN(ab_16__18_) );
  NOR2_X1 U539 ( .A1(n21), .A2(n44), .ZN(ab_16__17_) );
  NOR2_X1 U540 ( .A1(n22), .A2(n44), .ZN(ab_16__16_) );
  NOR2_X1 U541 ( .A1(n23), .A2(n44), .ZN(ab_16__15_) );
  NOR2_X1 U542 ( .A1(n24), .A2(n44), .ZN(ab_16__14_) );
  NOR2_X1 U543 ( .A1(n25), .A2(n44), .ZN(ab_16__13_) );
  NOR2_X1 U544 ( .A1(n26), .A2(n44), .ZN(ab_16__12_) );
  NOR2_X1 U545 ( .A1(n27), .A2(n44), .ZN(ab_16__11_) );
  NOR2_X1 U546 ( .A1(n28), .A2(n44), .ZN(ab_16__10_) );
  NOR2_X1 U547 ( .A1(n29), .A2(n44), .ZN(ab_16__0_) );
  NOR2_X1 U548 ( .A1(n7), .A2(n45), .ZN(ab_15__9_) );
  NOR2_X1 U549 ( .A1(n8), .A2(n45), .ZN(ab_15__8_) );
  NOR2_X1 U550 ( .A1(n9), .A2(n45), .ZN(ab_15__7_) );
  NOR2_X1 U551 ( .A1(n10), .A2(n45), .ZN(ab_15__6_) );
  NOR2_X1 U552 ( .A1(n11), .A2(n45), .ZN(ab_15__5_) );
  NOR2_X1 U553 ( .A1(n12), .A2(n45), .ZN(ab_15__4_) );
  NOR2_X1 U554 ( .A1(n13), .A2(n45), .ZN(ab_15__3_) );
  NOR2_X1 U555 ( .A1(n14), .A2(n45), .ZN(ab_15__2_) );
  NOR2_X1 U556 ( .A1(A[15]), .A2(n1), .ZN(ab_15__23_) );
  NOR2_X1 U557 ( .A1(n15), .A2(n45), .ZN(ab_15__22_) );
  NOR2_X1 U558 ( .A1(n16), .A2(n45), .ZN(ab_15__21_) );
  NOR2_X1 U559 ( .A1(n17), .A2(n45), .ZN(ab_15__20_) );
  NOR2_X1 U560 ( .A1(n18), .A2(n45), .ZN(ab_15__1_) );
  NOR2_X1 U561 ( .A1(n19), .A2(n45), .ZN(ab_15__19_) );
  NOR2_X1 U562 ( .A1(n20), .A2(n45), .ZN(ab_15__18_) );
  NOR2_X1 U563 ( .A1(n21), .A2(n45), .ZN(ab_15__17_) );
  NOR2_X1 U564 ( .A1(n22), .A2(n45), .ZN(ab_15__16_) );
  NOR2_X1 U565 ( .A1(n23), .A2(n45), .ZN(ab_15__15_) );
  NOR2_X1 U566 ( .A1(n24), .A2(n45), .ZN(ab_15__14_) );
  NOR2_X1 U567 ( .A1(n25), .A2(n45), .ZN(ab_15__13_) );
  NOR2_X1 U568 ( .A1(n26), .A2(n45), .ZN(ab_15__12_) );
  NOR2_X1 U569 ( .A1(n27), .A2(n45), .ZN(ab_15__11_) );
  NOR2_X1 U570 ( .A1(n28), .A2(n45), .ZN(ab_15__10_) );
  NOR2_X1 U571 ( .A1(n29), .A2(n45), .ZN(ab_15__0_) );
  NOR2_X1 U572 ( .A1(n7), .A2(n46), .ZN(ab_14__9_) );
  NOR2_X1 U573 ( .A1(n8), .A2(n46), .ZN(ab_14__8_) );
  NOR2_X1 U574 ( .A1(n9), .A2(n46), .ZN(ab_14__7_) );
  NOR2_X1 U575 ( .A1(n10), .A2(n46), .ZN(ab_14__6_) );
  NOR2_X1 U576 ( .A1(n11), .A2(n46), .ZN(ab_14__5_) );
  NOR2_X1 U577 ( .A1(n12), .A2(n46), .ZN(ab_14__4_) );
  NOR2_X1 U578 ( .A1(n13), .A2(n46), .ZN(ab_14__3_) );
  NOR2_X1 U579 ( .A1(n14), .A2(n46), .ZN(ab_14__2_) );
  NOR2_X1 U580 ( .A1(A[14]), .A2(n2), .ZN(ab_14__23_) );
  NOR2_X1 U581 ( .A1(n15), .A2(n46), .ZN(ab_14__22_) );
  NOR2_X1 U582 ( .A1(n16), .A2(n46), .ZN(ab_14__21_) );
  NOR2_X1 U583 ( .A1(n17), .A2(n46), .ZN(ab_14__20_) );
  NOR2_X1 U584 ( .A1(n18), .A2(n46), .ZN(ab_14__1_) );
  NOR2_X1 U585 ( .A1(n19), .A2(n46), .ZN(ab_14__19_) );
  NOR2_X1 U586 ( .A1(n20), .A2(n46), .ZN(ab_14__18_) );
  NOR2_X1 U587 ( .A1(n21), .A2(n46), .ZN(ab_14__17_) );
  NOR2_X1 U588 ( .A1(n22), .A2(n46), .ZN(ab_14__16_) );
  NOR2_X1 U589 ( .A1(n23), .A2(n46), .ZN(ab_14__15_) );
  NOR2_X1 U590 ( .A1(n24), .A2(n46), .ZN(ab_14__14_) );
  NOR2_X1 U591 ( .A1(n25), .A2(n46), .ZN(ab_14__13_) );
  NOR2_X1 U592 ( .A1(n26), .A2(n46), .ZN(ab_14__12_) );
  NOR2_X1 U593 ( .A1(n27), .A2(n46), .ZN(ab_14__11_) );
  NOR2_X1 U594 ( .A1(n28), .A2(n46), .ZN(ab_14__10_) );
  NOR2_X1 U595 ( .A1(n29), .A2(n46), .ZN(ab_14__0_) );
  NOR2_X1 U596 ( .A1(n7), .A2(n47), .ZN(ab_13__9_) );
  NOR2_X1 U597 ( .A1(n8), .A2(n47), .ZN(ab_13__8_) );
  NOR2_X1 U598 ( .A1(n9), .A2(n47), .ZN(ab_13__7_) );
  NOR2_X1 U599 ( .A1(n10), .A2(n47), .ZN(ab_13__6_) );
  NOR2_X1 U600 ( .A1(n11), .A2(n47), .ZN(ab_13__5_) );
  NOR2_X1 U601 ( .A1(n12), .A2(n47), .ZN(ab_13__4_) );
  NOR2_X1 U602 ( .A1(n13), .A2(n47), .ZN(ab_13__3_) );
  NOR2_X1 U603 ( .A1(n14), .A2(n47), .ZN(ab_13__2_) );
  NOR2_X1 U604 ( .A1(A[13]), .A2(n2), .ZN(ab_13__23_) );
  NOR2_X1 U605 ( .A1(n15), .A2(n47), .ZN(ab_13__22_) );
  NOR2_X1 U606 ( .A1(n16), .A2(n47), .ZN(ab_13__21_) );
  NOR2_X1 U607 ( .A1(n17), .A2(n47), .ZN(ab_13__20_) );
  NOR2_X1 U608 ( .A1(n18), .A2(n47), .ZN(ab_13__1_) );
  NOR2_X1 U609 ( .A1(n19), .A2(n47), .ZN(ab_13__19_) );
  NOR2_X1 U610 ( .A1(n20), .A2(n47), .ZN(ab_13__18_) );
  NOR2_X1 U611 ( .A1(n21), .A2(n47), .ZN(ab_13__17_) );
  NOR2_X1 U612 ( .A1(n22), .A2(n47), .ZN(ab_13__16_) );
  NOR2_X1 U613 ( .A1(n23), .A2(n47), .ZN(ab_13__15_) );
  NOR2_X1 U614 ( .A1(n24), .A2(n47), .ZN(ab_13__14_) );
  NOR2_X1 U615 ( .A1(n25), .A2(n47), .ZN(ab_13__13_) );
  NOR2_X1 U616 ( .A1(n26), .A2(n47), .ZN(ab_13__12_) );
  NOR2_X1 U617 ( .A1(n27), .A2(n47), .ZN(ab_13__11_) );
  NOR2_X1 U618 ( .A1(n28), .A2(n47), .ZN(ab_13__10_) );
  NOR2_X1 U619 ( .A1(n29), .A2(n47), .ZN(ab_13__0_) );
  NOR2_X1 U620 ( .A1(n7), .A2(n48), .ZN(ab_12__9_) );
  NOR2_X1 U621 ( .A1(n8), .A2(n48), .ZN(ab_12__8_) );
  NOR2_X1 U622 ( .A1(n9), .A2(n48), .ZN(ab_12__7_) );
  NOR2_X1 U623 ( .A1(n10), .A2(n48), .ZN(ab_12__6_) );
  NOR2_X1 U624 ( .A1(n11), .A2(n48), .ZN(ab_12__5_) );
  NOR2_X1 U625 ( .A1(n12), .A2(n48), .ZN(ab_12__4_) );
  NOR2_X1 U626 ( .A1(n13), .A2(n48), .ZN(ab_12__3_) );
  NOR2_X1 U627 ( .A1(n14), .A2(n48), .ZN(ab_12__2_) );
  NOR2_X1 U628 ( .A1(A[12]), .A2(n2), .ZN(ab_12__23_) );
  NOR2_X1 U629 ( .A1(n15), .A2(n48), .ZN(ab_12__22_) );
  NOR2_X1 U630 ( .A1(n16), .A2(n48), .ZN(ab_12__21_) );
  NOR2_X1 U631 ( .A1(n17), .A2(n48), .ZN(ab_12__20_) );
  NOR2_X1 U632 ( .A1(n18), .A2(n48), .ZN(ab_12__1_) );
  NOR2_X1 U633 ( .A1(n19), .A2(n48), .ZN(ab_12__19_) );
  NOR2_X1 U634 ( .A1(n20), .A2(n48), .ZN(ab_12__18_) );
  NOR2_X1 U635 ( .A1(n21), .A2(n48), .ZN(ab_12__17_) );
  NOR2_X1 U636 ( .A1(n22), .A2(n48), .ZN(ab_12__16_) );
  NOR2_X1 U637 ( .A1(n23), .A2(n48), .ZN(ab_12__15_) );
  NOR2_X1 U638 ( .A1(n24), .A2(n48), .ZN(ab_12__14_) );
  NOR2_X1 U639 ( .A1(n25), .A2(n48), .ZN(ab_12__13_) );
  NOR2_X1 U640 ( .A1(n26), .A2(n48), .ZN(ab_12__12_) );
  NOR2_X1 U641 ( .A1(n27), .A2(n48), .ZN(ab_12__11_) );
  NOR2_X1 U642 ( .A1(n28), .A2(n48), .ZN(ab_12__10_) );
  NOR2_X1 U643 ( .A1(n29), .A2(n48), .ZN(ab_12__0_) );
  NOR2_X1 U644 ( .A1(n7), .A2(n49), .ZN(ab_11__9_) );
  NOR2_X1 U645 ( .A1(n8), .A2(n49), .ZN(ab_11__8_) );
  NOR2_X1 U646 ( .A1(n9), .A2(n49), .ZN(ab_11__7_) );
  NOR2_X1 U647 ( .A1(n10), .A2(n49), .ZN(ab_11__6_) );
  NOR2_X1 U648 ( .A1(n11), .A2(n49), .ZN(ab_11__5_) );
  NOR2_X1 U649 ( .A1(n12), .A2(n49), .ZN(ab_11__4_) );
  NOR2_X1 U650 ( .A1(n13), .A2(n49), .ZN(ab_11__3_) );
  NOR2_X1 U651 ( .A1(n14), .A2(n49), .ZN(ab_11__2_) );
  NOR2_X1 U652 ( .A1(A[11]), .A2(n2), .ZN(ab_11__23_) );
  NOR2_X1 U653 ( .A1(n15), .A2(n49), .ZN(ab_11__22_) );
  NOR2_X1 U654 ( .A1(n16), .A2(n49), .ZN(ab_11__21_) );
  NOR2_X1 U655 ( .A1(n17), .A2(n49), .ZN(ab_11__20_) );
  NOR2_X1 U656 ( .A1(n18), .A2(n49), .ZN(ab_11__1_) );
  NOR2_X1 U657 ( .A1(n19), .A2(n49), .ZN(ab_11__19_) );
  NOR2_X1 U658 ( .A1(n20), .A2(n49), .ZN(ab_11__18_) );
  NOR2_X1 U659 ( .A1(n21), .A2(n49), .ZN(ab_11__17_) );
  NOR2_X1 U660 ( .A1(n22), .A2(n49), .ZN(ab_11__16_) );
  NOR2_X1 U661 ( .A1(n23), .A2(n49), .ZN(ab_11__15_) );
  NOR2_X1 U662 ( .A1(n24), .A2(n49), .ZN(ab_11__14_) );
  NOR2_X1 U663 ( .A1(n25), .A2(n49), .ZN(ab_11__13_) );
  NOR2_X1 U664 ( .A1(n26), .A2(n49), .ZN(ab_11__12_) );
  NOR2_X1 U665 ( .A1(n27), .A2(n49), .ZN(ab_11__11_) );
  NOR2_X1 U666 ( .A1(n28), .A2(n49), .ZN(ab_11__10_) );
  NOR2_X1 U667 ( .A1(n29), .A2(n49), .ZN(ab_11__0_) );
  NOR2_X1 U668 ( .A1(n7), .A2(n50), .ZN(ab_10__9_) );
  NOR2_X1 U669 ( .A1(n8), .A2(n50), .ZN(ab_10__8_) );
  NOR2_X1 U670 ( .A1(n9), .A2(n50), .ZN(ab_10__7_) );
  NOR2_X1 U671 ( .A1(n10), .A2(n50), .ZN(ab_10__6_) );
  NOR2_X1 U672 ( .A1(n11), .A2(n50), .ZN(ab_10__5_) );
  NOR2_X1 U673 ( .A1(n12), .A2(n50), .ZN(ab_10__4_) );
  NOR2_X1 U674 ( .A1(n13), .A2(n50), .ZN(ab_10__3_) );
  NOR2_X1 U675 ( .A1(n14), .A2(n50), .ZN(ab_10__2_) );
  NOR2_X1 U676 ( .A1(A[10]), .A2(n2), .ZN(ab_10__23_) );
  NOR2_X1 U677 ( .A1(n15), .A2(n50), .ZN(ab_10__22_) );
  NOR2_X1 U678 ( .A1(n16), .A2(n50), .ZN(ab_10__21_) );
  NOR2_X1 U679 ( .A1(n17), .A2(n50), .ZN(ab_10__20_) );
  NOR2_X1 U680 ( .A1(n18), .A2(n50), .ZN(ab_10__1_) );
  NOR2_X1 U681 ( .A1(n19), .A2(n50), .ZN(ab_10__19_) );
  NOR2_X1 U682 ( .A1(n20), .A2(n50), .ZN(ab_10__18_) );
  NOR2_X1 U683 ( .A1(n21), .A2(n50), .ZN(ab_10__17_) );
  NOR2_X1 U684 ( .A1(n22), .A2(n50), .ZN(ab_10__16_) );
  NOR2_X1 U685 ( .A1(n23), .A2(n50), .ZN(ab_10__15_) );
  NOR2_X1 U686 ( .A1(n24), .A2(n50), .ZN(ab_10__14_) );
  NOR2_X1 U687 ( .A1(n25), .A2(n50), .ZN(ab_10__13_) );
  NOR2_X1 U688 ( .A1(n26), .A2(n50), .ZN(ab_10__12_) );
  NOR2_X1 U689 ( .A1(n27), .A2(n50), .ZN(ab_10__11_) );
  NOR2_X1 U690 ( .A1(n28), .A2(n50), .ZN(ab_10__10_) );
  NOR2_X1 U691 ( .A1(n29), .A2(n50), .ZN(ab_10__0_) );
  NOR2_X1 U692 ( .A1(n7), .A2(n51), .ZN(ab_0__9_) );
  NOR2_X1 U693 ( .A1(n8), .A2(n51), .ZN(ab_0__8_) );
  NOR2_X1 U694 ( .A1(n9), .A2(n51), .ZN(ab_0__7_) );
  NOR2_X1 U695 ( .A1(n10), .A2(n51), .ZN(ab_0__6_) );
  NOR2_X1 U696 ( .A1(n11), .A2(n51), .ZN(ab_0__5_) );
  NOR2_X1 U697 ( .A1(n12), .A2(n51), .ZN(ab_0__4_) );
  NOR2_X1 U698 ( .A1(n13), .A2(n51), .ZN(ab_0__3_) );
  NOR2_X1 U699 ( .A1(n14), .A2(n51), .ZN(ab_0__2_) );
  NOR2_X1 U700 ( .A1(A[0]), .A2(n1), .ZN(ab_0__23_) );
  NOR2_X1 U701 ( .A1(n15), .A2(n51), .ZN(ab_0__22_) );
  NOR2_X1 U702 ( .A1(n16), .A2(n51), .ZN(ab_0__21_) );
  NOR2_X1 U703 ( .A1(n17), .A2(n51), .ZN(ab_0__20_) );
  NOR2_X1 U704 ( .A1(n19), .A2(n51), .ZN(ab_0__19_) );
  NOR2_X1 U705 ( .A1(n20), .A2(n51), .ZN(ab_0__18_) );
  NOR2_X1 U706 ( .A1(n21), .A2(n51), .ZN(ab_0__17_) );
  NOR2_X1 U707 ( .A1(n22), .A2(n51), .ZN(ab_0__16_) );
  NOR2_X1 U708 ( .A1(n23), .A2(n51), .ZN(ab_0__15_) );
  NOR2_X1 U709 ( .A1(n24), .A2(n51), .ZN(ab_0__14_) );
  NOR2_X1 U710 ( .A1(n25), .A2(n51), .ZN(ab_0__13_) );
  NOR2_X1 U711 ( .A1(n26), .A2(n51), .ZN(ab_0__12_) );
  NOR2_X1 U712 ( .A1(n27), .A2(n51), .ZN(ab_0__11_) );
  NOR2_X1 U713 ( .A1(n28), .A2(n51), .ZN(ab_0__10_) );
  INV_X1 U714 ( .A(B[23]), .ZN(QB) );
  INV_X1 U715 ( .A(A[23]), .ZN(QA) );
  AND3_X1 U716 ( .A1(ab_1__1_), .A2(B[0]), .A3(A[0]), .ZN(CARRYB_1__0_) );
  NOR2_X1 U717 ( .A1(n40), .A2(n18), .ZN(ab_1__1_) );
  INV_X1 U719 ( .A(CARRYB_23__23_), .ZN(A1_45_) );
endmodule


module iir_filter_DW01_add_3 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   carry_23_, carry_22_, carry_21_, carry_20_, carry_19_, carry_18_,
         carry_17_, carry_16_, carry_15_, carry_14_, carry_13_, carry_12_,
         carry_11_, carry_10_, carry_9_, carry_8_, carry_7_, carry_6_,
         carry_5_, carry_4_, carry_3_, carry_2_, carry_1_;

  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry_23_), .S(SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry_22_), .CO(carry_23_), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry_21_), .CO(carry_22_), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry_20_), .CO(carry_21_), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry_19_), .CO(carry_20_), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry_18_), .CO(carry_19_), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry_17_), .CO(carry_18_), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry_16_), .CO(carry_17_), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry_15_), .CO(carry_16_), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry_14_), .CO(carry_15_), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry_13_), .CO(carry_14_), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry_12_), .CO(carry_13_), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry_11_), .CO(carry_12_), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry_10_), .CO(carry_11_), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry_9_), .CO(carry_10_), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry_8_), .CO(carry_9_), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry_7_), .CO(carry_8_), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry_6_), .CO(carry_7_), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry_5_), .CO(carry_6_), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry_4_), .CO(carry_5_), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry_3_), .CO(carry_4_), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry_2_), .CO(carry_3_), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry_1_), .CO(carry_2_), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(A[0]), .A2(B[0]), .ZN(carry_1_) );
  XOR2_X1 U2 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module iir_filter_DW01_add_2 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   carry_23_, carry_22_, carry_21_, carry_20_, carry_19_, carry_18_,
         carry_17_, carry_16_, carry_15_, carry_14_, carry_13_, carry_12_,
         carry_11_, carry_10_, carry_9_, carry_8_, carry_7_, carry_6_,
         carry_5_, carry_4_, carry_3_, carry_2_, carry_1_;

  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry_23_), .S(SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry_22_), .CO(carry_23_), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry_21_), .CO(carry_22_), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry_20_), .CO(carry_21_), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry_19_), .CO(carry_20_), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry_18_), .CO(carry_19_), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry_17_), .CO(carry_18_), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry_16_), .CO(carry_17_), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry_15_), .CO(carry_16_), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry_14_), .CO(carry_15_), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry_13_), .CO(carry_14_), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry_12_), .CO(carry_13_), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry_11_), .CO(carry_12_), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry_10_), .CO(carry_11_), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry_9_), .CO(carry_10_), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry_8_), .CO(carry_9_), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry_7_), .CO(carry_8_), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry_6_), .CO(carry_7_), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry_5_), .CO(carry_6_), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry_4_), .CO(carry_5_), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry_3_), .CO(carry_4_), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry_2_), .CO(carry_3_), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry_1_), .CO(carry_2_), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(A[0]), .A2(B[0]), .ZN(carry_1_) );
  XOR2_X1 U2 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module iir_filter_DW01_add_1 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   carry_23_, carry_22_, carry_21_, carry_20_, carry_19_, carry_18_,
         carry_17_, carry_16_, carry_15_, carry_14_, carry_13_, carry_12_,
         carry_11_, carry_10_, carry_9_, carry_8_, carry_7_, carry_6_,
         carry_5_, carry_4_, carry_3_, carry_2_, carry_1_;

  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry_23_), .S(SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry_22_), .CO(carry_23_), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry_21_), .CO(carry_22_), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry_20_), .CO(carry_21_), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry_19_), .CO(carry_20_), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry_18_), .CO(carry_19_), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry_17_), .CO(carry_18_), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry_16_), .CO(carry_17_), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry_15_), .CO(carry_16_), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry_14_), .CO(carry_15_), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry_13_), .CO(carry_14_), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry_12_), .CO(carry_13_), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry_11_), .CO(carry_12_), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry_10_), .CO(carry_11_), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry_9_), .CO(carry_10_), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry_8_), .CO(carry_9_), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry_7_), .CO(carry_8_), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry_6_), .CO(carry_7_), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry_5_), .CO(carry_6_), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry_4_), .CO(carry_5_), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry_3_), .CO(carry_4_), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry_2_), .CO(carry_3_), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry_1_), .CO(carry_2_), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(A[0]), .A2(B[0]), .ZN(carry_1_) );
  XOR2_X1 U2 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module iir_filter_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] DIFF;
  input CI;
  output CO;
  wire   B_0_, carry_23_, carry_22_, carry_21_, carry_20_, carry_19_,
         carry_18_, carry_17_, carry_16_, carry_15_, carry_14_, carry_13_,
         carry_12_, carry_11_, carry_10_, carry_9_, carry_8_, carry_7_,
         carry_6_, carry_5_, carry_4_, carry_3_, carry_2_, carry_1_, B_not_23_,
         B_not_22_, B_not_21_, B_not_20_, B_not_19_, B_not_18_, B_not_17_,
         B_not_16_, B_not_15_, B_not_14_, B_not_13_, B_not_12_, B_not_11_,
         B_not_10_, B_not_9_, B_not_8_, B_not_7_, B_not_6_, B_not_5_, B_not_4_,
         B_not_3_, B_not_2_, B_not_1_;
  assign DIFF[0] = B_0_;
  assign B_0_ = B[0];

  FA_X1 U2_23 ( .A(A[23]), .B(B_not_23_), .CI(carry_23_), .S(DIFF[23]) );
  FA_X1 U2_22 ( .A(A[22]), .B(B_not_22_), .CI(carry_22_), .CO(carry_23_), .S(
        DIFF[22]) );
  FA_X1 U2_21 ( .A(A[21]), .B(B_not_21_), .CI(carry_21_), .CO(carry_22_), .S(
        DIFF[21]) );
  FA_X1 U2_20 ( .A(A[20]), .B(B_not_20_), .CI(carry_20_), .CO(carry_21_), .S(
        DIFF[20]) );
  FA_X1 U2_19 ( .A(A[19]), .B(B_not_19_), .CI(carry_19_), .CO(carry_20_), .S(
        DIFF[19]) );
  FA_X1 U2_18 ( .A(A[18]), .B(B_not_18_), .CI(carry_18_), .CO(carry_19_), .S(
        DIFF[18]) );
  FA_X1 U2_17 ( .A(A[17]), .B(B_not_17_), .CI(carry_17_), .CO(carry_18_), .S(
        DIFF[17]) );
  FA_X1 U2_16 ( .A(A[16]), .B(B_not_16_), .CI(carry_16_), .CO(carry_17_), .S(
        DIFF[16]) );
  FA_X1 U2_15 ( .A(A[15]), .B(B_not_15_), .CI(carry_15_), .CO(carry_16_), .S(
        DIFF[15]) );
  FA_X1 U2_14 ( .A(A[14]), .B(B_not_14_), .CI(carry_14_), .CO(carry_15_), .S(
        DIFF[14]) );
  FA_X1 U2_13 ( .A(A[13]), .B(B_not_13_), .CI(carry_13_), .CO(carry_14_), .S(
        DIFF[13]) );
  FA_X1 U2_12 ( .A(A[12]), .B(B_not_12_), .CI(carry_12_), .CO(carry_13_), .S(
        DIFF[12]) );
  FA_X1 U2_11 ( .A(A[11]), .B(B_not_11_), .CI(carry_11_), .CO(carry_12_), .S(
        DIFF[11]) );
  AND2_X1 U1 ( .A1(carry_10_), .A2(B_not_10_), .ZN(carry_11_) );
  XOR2_X1 U2 ( .A(B_not_10_), .B(carry_10_), .Z(DIFF[10]) );
  AND2_X1 U3 ( .A1(carry_9_), .A2(B_not_9_), .ZN(carry_10_) );
  XOR2_X1 U4 ( .A(B_not_9_), .B(carry_9_), .Z(DIFF[9]) );
  AND2_X1 U5 ( .A1(carry_8_), .A2(B_not_8_), .ZN(carry_9_) );
  XOR2_X1 U6 ( .A(B_not_8_), .B(carry_8_), .Z(DIFF[8]) );
  AND2_X1 U7 ( .A1(carry_7_), .A2(B_not_7_), .ZN(carry_8_) );
  XOR2_X1 U8 ( .A(B_not_7_), .B(carry_7_), .Z(DIFF[7]) );
  AND2_X1 U9 ( .A1(carry_6_), .A2(B_not_6_), .ZN(carry_7_) );
  XOR2_X1 U10 ( .A(B_not_6_), .B(carry_6_), .Z(DIFF[6]) );
  AND2_X1 U11 ( .A1(carry_5_), .A2(B_not_5_), .ZN(carry_6_) );
  XOR2_X1 U12 ( .A(B_not_5_), .B(carry_5_), .Z(DIFF[5]) );
  AND2_X1 U13 ( .A1(carry_4_), .A2(B_not_4_), .ZN(carry_5_) );
  XOR2_X1 U14 ( .A(B_not_4_), .B(carry_4_), .Z(DIFF[4]) );
  AND2_X1 U15 ( .A1(carry_3_), .A2(B_not_3_), .ZN(carry_4_) );
  XOR2_X1 U16 ( .A(B_not_3_), .B(carry_3_), .Z(DIFF[3]) );
  AND2_X1 U17 ( .A1(carry_2_), .A2(B_not_2_), .ZN(carry_3_) );
  XOR2_X1 U18 ( .A(B_not_2_), .B(carry_2_), .Z(DIFF[2]) );
  AND2_X1 U19 ( .A1(carry_1_), .A2(B_not_1_), .ZN(carry_2_) );
  XOR2_X1 U20 ( .A(B_not_1_), .B(carry_1_), .Z(DIFF[1]) );
  INV_X1 U21 ( .A(B_0_), .ZN(carry_1_) );
  INV_X1 U22 ( .A(B[9]), .ZN(B_not_9_) );
  INV_X1 U23 ( .A(B[8]), .ZN(B_not_8_) );
  INV_X1 U24 ( .A(B[7]), .ZN(B_not_7_) );
  INV_X1 U25 ( .A(B[6]), .ZN(B_not_6_) );
  INV_X1 U26 ( .A(B[5]), .ZN(B_not_5_) );
  INV_X1 U27 ( .A(B[4]), .ZN(B_not_4_) );
  INV_X1 U28 ( .A(B[3]), .ZN(B_not_3_) );
  INV_X1 U29 ( .A(B[2]), .ZN(B_not_2_) );
  INV_X1 U30 ( .A(B[23]), .ZN(B_not_23_) );
  INV_X1 U31 ( .A(B[22]), .ZN(B_not_22_) );
  INV_X1 U32 ( .A(B[21]), .ZN(B_not_21_) );
  INV_X1 U33 ( .A(B[20]), .ZN(B_not_20_) );
  INV_X1 U34 ( .A(B[1]), .ZN(B_not_1_) );
  INV_X1 U35 ( .A(B[19]), .ZN(B_not_19_) );
  INV_X1 U36 ( .A(B[18]), .ZN(B_not_18_) );
  INV_X1 U37 ( .A(B[17]), .ZN(B_not_17_) );
  INV_X1 U38 ( .A(B[16]), .ZN(B_not_16_) );
  INV_X1 U39 ( .A(B[15]), .ZN(B_not_15_) );
  INV_X1 U40 ( .A(B[14]), .ZN(B_not_14_) );
  INV_X1 U41 ( .A(B[13]), .ZN(B_not_13_) );
  INV_X1 U42 ( .A(B[12]), .ZN(B_not_12_) );
  INV_X1 U43 ( .A(B[11]), .ZN(B_not_11_) );
  INV_X1 U44 ( .A(B[10]), .ZN(B_not_10_) );
endmodule


module iir_filter_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   carry_23_, carry_22_, carry_21_, carry_20_, carry_19_, carry_18_,
         carry_17_, carry_16_, carry_15_, carry_14_, carry_13_, carry_12_,
         carry_11_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37;

  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry_23_), .S(SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry_22_), .CO(carry_23_), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry_21_), .CO(carry_22_), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry_20_), .CO(carry_21_), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry_19_), .CO(carry_20_), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry_18_), .CO(carry_19_), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry_17_), .CO(carry_18_), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry_16_), .CO(carry_17_), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry_15_), .CO(carry_16_), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry_14_), .CO(carry_15_), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry_13_), .CO(carry_14_), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry_12_), .CO(carry_13_), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry_11_), .CO(carry_12_), .S(
        SUM[11]) );
  OAI21_X1 U1 ( .B1(n1), .B2(n2), .A(n3), .ZN(carry_11_) );
  OAI21_X1 U2 ( .B1(A[10]), .B2(n4), .A(B[10]), .ZN(n3) );
  INV_X1 U3 ( .A(n1), .ZN(n4) );
  INV_X1 U4 ( .A(A[10]), .ZN(n2) );
  AOI21_X1 U5 ( .B1(n5), .B2(A[9]), .A(n6), .ZN(n1) );
  INV_X1 U6 ( .A(n7), .ZN(n6) );
  OAI21_X1 U7 ( .B1(A[9]), .B2(n5), .A(B[9]), .ZN(n7) );
  OAI21_X1 U8 ( .B1(n8), .B2(n9), .A(n10), .ZN(n5) );
  OAI21_X1 U9 ( .B1(A[8]), .B2(n11), .A(B[8]), .ZN(n10) );
  INV_X1 U10 ( .A(n8), .ZN(n11) );
  INV_X1 U11 ( .A(A[8]), .ZN(n9) );
  AOI21_X1 U12 ( .B1(n12), .B2(A[7]), .A(n13), .ZN(n8) );
  INV_X1 U13 ( .A(n14), .ZN(n13) );
  OAI21_X1 U14 ( .B1(A[7]), .B2(n12), .A(B[7]), .ZN(n14) );
  OAI21_X1 U15 ( .B1(n15), .B2(n16), .A(n17), .ZN(n12) );
  OAI21_X1 U16 ( .B1(A[6]), .B2(n18), .A(B[6]), .ZN(n17) );
  INV_X1 U17 ( .A(A[6]), .ZN(n16) );
  INV_X1 U18 ( .A(n18), .ZN(n15) );
  OAI21_X1 U19 ( .B1(n19), .B2(n20), .A(n21), .ZN(n18) );
  OAI21_X1 U20 ( .B1(A[5]), .B2(n22), .A(B[5]), .ZN(n21) );
  INV_X1 U21 ( .A(A[5]), .ZN(n20) );
  INV_X1 U22 ( .A(n22), .ZN(n19) );
  OAI21_X1 U23 ( .B1(n23), .B2(n24), .A(n25), .ZN(n22) );
  OAI21_X1 U24 ( .B1(A[4]), .B2(n26), .A(B[4]), .ZN(n25) );
  INV_X1 U25 ( .A(A[4]), .ZN(n24) );
  INV_X1 U26 ( .A(n26), .ZN(n23) );
  OAI21_X1 U27 ( .B1(n27), .B2(n28), .A(n29), .ZN(n26) );
  OAI21_X1 U28 ( .B1(A[3]), .B2(n30), .A(B[3]), .ZN(n29) );
  INV_X1 U29 ( .A(A[3]), .ZN(n28) );
  INV_X1 U30 ( .A(n30), .ZN(n27) );
  OAI21_X1 U31 ( .B1(n31), .B2(n32), .A(n33), .ZN(n30) );
  OAI21_X1 U32 ( .B1(A[2]), .B2(n34), .A(B[2]), .ZN(n33) );
  INV_X1 U33 ( .A(A[2]), .ZN(n32) );
  INV_X1 U34 ( .A(n34), .ZN(n31) );
  OAI21_X1 U35 ( .B1(n35), .B2(n36), .A(n37), .ZN(n34) );
  OAI211_X1 U36 ( .C1(A[1]), .C2(B[1]), .A(A[0]), .B(B[0]), .ZN(n37) );
  INV_X1 U37 ( .A(B[1]), .ZN(n36) );
  INV_X1 U38 ( .A(A[1]), .ZN(n35) );
endmodule


module iir_filter ( clk, rst_n, vIn, dIn, coeffs_fb, coeffs_ff, dOut, vOut );
  input [11:0] dIn;
  input [47:0] coeffs_fb;
  input [95:0] coeffs_ff;
  output [11:0] dOut;
  input clk, rst_n, vIn;
  output vOut;
  wire   delayed_controls_0__1_, delayed_controls_1__0_,
         delayed_controls_1__1_, delayed_controls_2__0_, DP_N4, DP_N2, DP_y_0_,
         DP_y_1_, DP_y_2_, DP_y_3_, DP_y_4_, DP_y_5_, DP_y_6_, DP_y_7_,
         DP_y_8_, DP_y_9_, DP_y_10_, DP_y_11_, DP_y_23, DP_sw1_0_, DP_sw1_1_,
         DP_sw1_2_, DP_sw1_3_, DP_sw1_4_, DP_sw1_5_, DP_sw1_6_, DP_sw1_7_,
         DP_sw1_8_, DP_sw1_9_, DP_sw1_10_, DP_sw1_11_, DP_sw1_12_, DP_sw1_13_,
         DP_sw1_14_, DP_sw1_15_, DP_sw1_16_, DP_sw1_17_, DP_sw1_18_,
         DP_sw1_19_, DP_sw1_20_, DP_sw1_21_, DP_sw1_22_, DP_sw1_23_, DP_sw0_0_,
         DP_sw0_1_, DP_sw0_2_, DP_sw0_3_, DP_sw0_4_, DP_sw0_5_, DP_sw0_6_,
         DP_sw0_7_, DP_sw0_8_, DP_sw0_9_, DP_sw0_10_, DP_sw0_11_, DP_sw0_12_,
         DP_sw0_13_, DP_sw0_14_, DP_sw0_15_, DP_sw0_16_, DP_sw0_17_,
         DP_sw0_18_, DP_sw0_19_, DP_sw0_20_, DP_sw0_21_, DP_sw0_22_,
         DP_sw0_23_, DP_w_0_, DP_w_1_, DP_w_2_, DP_w_3_, DP_w_4_, DP_w_5_,
         DP_w_6_, DP_w_7_, DP_w_8_, DP_w_9_, DP_w_10_, DP_w_11_, DP_w_12_,
         DP_w_13_, DP_w_14_, DP_w_15_, DP_w_16_, DP_w_17_, DP_w_18_, DP_w_19_,
         DP_w_20_, DP_w_21_, DP_w_22_, DP_w_23_, CU_nextState_0_, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n72, n73, n74, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n560, n562, n564, n566, n568,
         n570, n572, n574, n576, n578, n580, n582, n584, n586, n588, n590,
         n592, n594, n596, n598, n600, n602, n604, n606, n706, n707, n711,
         n712, n716, n717, n721, n722, n726, n727, n731, n732, n736, n737,
         n741, n742, n746, n747, n751, n752, n756, n757, n761, n762, n766,
         n767, n771, n772, n776, n777, n781, n782, n786, n787, n791, n792,
         n796, n797, n801, n802, n806, n807, n811, n812, n816, n817, n820,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140;
  wire   [0:23] DP_ff;
  wire   [0:23] DP_ff_part;
  wire   [0:23] DP_fb;
  wire   [0:23] DP_pipe13;
  wire   [0:23] DP_pipe0_coeff_pipe03;
  wire   [0:23] DP_pipe12;
  wire   [0:23] DP_pipe0_coeff_pipe02;
  wire   [0:23] DP_pipe11;
  wire   [0:23] DP_pipe0_coeff_pipe01;
  wire   [0:23] DP_pipe10;
  wire   [0:23] DP_pipe0_coeff_pipe00;
  wire   [0:23] DP_pipe03;
  wire   [0:23] DP_pipe02;
  wire   [0:23] DP_pipe01;
  wire   [0:23] DP_pipe00;
  wire   [0:23] DP_ret1;
  wire   [0:23] DP_sw1_coeff_ret1;
  wire   [0:23] DP_ret0;
  wire   [0:23] DP_sw0_coeff_ret0;
  wire   [0:23] DP_sw2;
  wire   [95:0] DP_coeffs_ff_int;
  wire   [47:0] DP_coeffs_fb_int;
  wire   [0:11] DP_x;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154;

  DFFR_X1 DP_reg_in_Q_reg_0_ ( .D(n1002), .CK(clk), .RN(n1091), .Q(DP_x[0]), 
        .QN(n301) );
  DFFR_X1 DP_reg_in_Q_reg_1_ ( .D(n1001), .CK(clk), .RN(n1091), .Q(DP_x[1]), 
        .QN(n300) );
  DFFR_X1 DP_reg_in_Q_reg_2_ ( .D(n1000), .CK(clk), .RN(n1091), .Q(DP_x[2]), 
        .QN(n299) );
  DFFR_X1 DP_reg_in_Q_reg_3_ ( .D(n999), .CK(clk), .RN(n1091), .Q(DP_x[3]), 
        .QN(n298) );
  DFFR_X1 DP_reg_in_Q_reg_4_ ( .D(n998), .CK(clk), .RN(n1091), .Q(DP_x[4]), 
        .QN(n297) );
  DFFR_X1 DP_reg_in_Q_reg_5_ ( .D(n997), .CK(clk), .RN(n1091), .Q(DP_x[5]), 
        .QN(n296) );
  DFFR_X1 DP_reg_in_Q_reg_6_ ( .D(n996), .CK(clk), .RN(n1091), .Q(DP_x[6]), 
        .QN(n295) );
  DFFR_X1 DP_reg_in_Q_reg_7_ ( .D(n995), .CK(clk), .RN(n1091), .Q(DP_x[7]), 
        .QN(n294) );
  DFFR_X1 DP_reg_in_Q_reg_8_ ( .D(n994), .CK(clk), .RN(n1091), .Q(DP_x[8]), 
        .QN(n293) );
  DFFR_X1 DP_reg_in_Q_reg_9_ ( .D(n993), .CK(clk), .RN(n1091), .Q(DP_x[9]), 
        .QN(n292) );
  DFFR_X1 DP_reg_in_Q_reg_10_ ( .D(n992), .CK(clk), .RN(n1091), .Q(DP_x[10]), 
        .QN(n291) );
  DFFR_X1 DP_reg_in_Q_reg_11_ ( .D(n991), .CK(clk), .RN(n1091), .Q(DP_x[11]), 
        .QN(n290) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_0_ ( .D(n990), .CK(clk), .RN(n1092), .Q(
        DP_coeffs_fb_int[23]), .QN(n289) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_1_ ( .D(n989), .CK(clk), .RN(n1092), .Q(
        DP_coeffs_fb_int[22]), .QN(n288) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_2_ ( .D(n988), .CK(clk), .RN(n1092), .Q(
        DP_coeffs_fb_int[21]), .QN(n287) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_3_ ( .D(n987), .CK(clk), .RN(n1092), .Q(
        DP_coeffs_fb_int[20]), .QN(n286) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_4_ ( .D(n986), .CK(clk), .RN(n1092), .Q(
        DP_coeffs_fb_int[19]), .QN(n285) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_5_ ( .D(n985), .CK(clk), .RN(n1092), .Q(
        DP_coeffs_fb_int[18]), .QN(n284) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_6_ ( .D(n984), .CK(clk), .RN(n1092), .Q(
        DP_coeffs_fb_int[17]), .QN(n283) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_7_ ( .D(n983), .CK(clk), .RN(n1092), .Q(
        DP_coeffs_fb_int[16]), .QN(n282) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_8_ ( .D(n982), .CK(clk), .RN(n1092), .Q(
        DP_coeffs_fb_int[15]), .QN(n281) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_9_ ( .D(n981), .CK(clk), .RN(n1092), .Q(
        DP_coeffs_fb_int[14]), .QN(n280) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_10_ ( .D(n980), .CK(clk), .RN(n1092), .Q(
        DP_coeffs_fb_int[13]), .QN(n279) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_11_ ( .D(n979), .CK(clk), .RN(n1092), .Q(
        DP_coeffs_fb_int[12]), .QN(n278) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_12_ ( .D(n978), .CK(clk), .RN(n1093), .Q(
        DP_coeffs_fb_int[11]), .QN(n277) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_13_ ( .D(n977), .CK(clk), .RN(n1093), .Q(
        DP_coeffs_fb_int[10]), .QN(n519) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_14_ ( .D(n976), .CK(clk), .RN(n1093), .Q(
        DP_coeffs_fb_int[9]), .QN(n518) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_15_ ( .D(n975), .CK(clk), .RN(n1093), .Q(
        DP_coeffs_fb_int[8]), .QN(n517) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_16_ ( .D(n974), .CK(clk), .RN(n1093), .Q(
        DP_coeffs_fb_int[7]), .QN(n516) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_17_ ( .D(n973), .CK(clk), .RN(n1093), .Q(
        DP_coeffs_fb_int[6]), .QN(n515) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_18_ ( .D(n972), .CK(clk), .RN(n1093), .Q(
        DP_coeffs_fb_int[5]), .QN(n514) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_19_ ( .D(n971), .CK(clk), .RN(n1093), .Q(
        DP_coeffs_fb_int[4]), .QN(n513) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_20_ ( .D(n970), .CK(clk), .RN(n1093), .Q(
        DP_coeffs_fb_int[3]), .QN(n512) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_21_ ( .D(n969), .CK(clk), .RN(n1093), .Q(
        DP_coeffs_fb_int[2]), .QN(n511) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_22_ ( .D(n968), .CK(clk), .RN(n1093), .Q(
        DP_coeffs_fb_int[1]), .QN(n510) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_23_ ( .D(n967), .CK(clk), .RN(n1093), .Q(
        DP_coeffs_fb_int[0]), .QN(n509) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_0_ ( .D(n966), .CK(clk), .RN(n1094), .Q(
        DP_coeffs_fb_int[47]), .QN(n508) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_1_ ( .D(n965), .CK(clk), .RN(n1094), .Q(
        DP_coeffs_fb_int[46]), .QN(n507) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_2_ ( .D(n964), .CK(clk), .RN(n1094), .Q(
        DP_coeffs_fb_int[45]), .QN(n506) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_3_ ( .D(n963), .CK(clk), .RN(n1094), .Q(
        DP_coeffs_fb_int[44]), .QN(n505) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_4_ ( .D(n962), .CK(clk), .RN(n1094), .Q(
        DP_coeffs_fb_int[43]), .QN(n504) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_5_ ( .D(n961), .CK(clk), .RN(n1094), .Q(
        DP_coeffs_fb_int[42]), .QN(n503) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_6_ ( .D(n960), .CK(clk), .RN(n1094), .Q(
        DP_coeffs_fb_int[41]), .QN(n502) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_7_ ( .D(n959), .CK(clk), .RN(n1094), .Q(
        DP_coeffs_fb_int[40]), .QN(n501) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_8_ ( .D(n958), .CK(clk), .RN(n1094), .Q(
        DP_coeffs_fb_int[39]), .QN(n500) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_9_ ( .D(n957), .CK(clk), .RN(n1094), .Q(
        DP_coeffs_fb_int[38]), .QN(n499) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_10_ ( .D(n956), .CK(clk), .RN(n1094), .Q(
        DP_coeffs_fb_int[37]), .QN(n498) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_11_ ( .D(n955), .CK(clk), .RN(n1094), .Q(
        DP_coeffs_fb_int[36]), .QN(n497) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_12_ ( .D(n954), .CK(clk), .RN(n1095), .Q(
        DP_coeffs_fb_int[35]), .QN(n496) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_13_ ( .D(n953), .CK(clk), .RN(n1095), .Q(
        DP_coeffs_fb_int[34]), .QN(n495) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_14_ ( .D(n952), .CK(clk), .RN(n1095), .Q(
        DP_coeffs_fb_int[33]), .QN(n494) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_15_ ( .D(n951), .CK(clk), .RN(n1095), .Q(
        DP_coeffs_fb_int[32]), .QN(n493) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_16_ ( .D(n950), .CK(clk), .RN(n1095), .Q(
        DP_coeffs_fb_int[31]), .QN(n492) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_17_ ( .D(n949), .CK(clk), .RN(n1095), .Q(
        DP_coeffs_fb_int[30]), .QN(n491) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_18_ ( .D(n948), .CK(clk), .RN(n1095), .Q(
        DP_coeffs_fb_int[29]), .QN(n490) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_19_ ( .D(n947), .CK(clk), .RN(n1095), .Q(
        DP_coeffs_fb_int[28]), .QN(n489) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_20_ ( .D(n946), .CK(clk), .RN(n1095), .Q(
        DP_coeffs_fb_int[27]), .QN(n488) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_21_ ( .D(n945), .CK(clk), .RN(n1095), .Q(
        DP_coeffs_fb_int[26]), .QN(n487) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_22_ ( .D(n944), .CK(clk), .RN(n1095), .Q(
        DP_coeffs_fb_int[25]), .QN(n486) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_23_ ( .D(n943), .CK(clk), .RN(n1095), .Q(
        DP_coeffs_fb_int[24]), .QN(n485) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_0_ ( .D(n942), .CK(clk), .RN(n1096), .Q(
        DP_coeffs_ff_int[23]), .QN(n484) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_1_ ( .D(n941), .CK(clk), .RN(n1096), .Q(
        DP_coeffs_ff_int[22]), .QN(n483) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_2_ ( .D(n940), .CK(clk), .RN(n1096), .Q(
        DP_coeffs_ff_int[21]), .QN(n482) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_3_ ( .D(n939), .CK(clk), .RN(n1096), .Q(
        DP_coeffs_ff_int[20]), .QN(n481) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_4_ ( .D(n938), .CK(clk), .RN(n1096), .Q(
        DP_coeffs_ff_int[19]), .QN(n480) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_5_ ( .D(n937), .CK(clk), .RN(n1096), .Q(
        DP_coeffs_ff_int[18]), .QN(n479) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_6_ ( .D(n936), .CK(clk), .RN(n1096), .Q(
        DP_coeffs_ff_int[17]), .QN(n478) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_7_ ( .D(n935), .CK(clk), .RN(n1096), .Q(
        DP_coeffs_ff_int[16]), .QN(n477) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_8_ ( .D(n934), .CK(clk), .RN(n1096), .Q(
        DP_coeffs_ff_int[15]), .QN(n476) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_9_ ( .D(n933), .CK(clk), .RN(n1096), .Q(
        DP_coeffs_ff_int[14]), .QN(n475) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_10_ ( .D(n932), .CK(clk), .RN(n1096), .Q(
        DP_coeffs_ff_int[13]), .QN(n474) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_11_ ( .D(n931), .CK(clk), .RN(n1096), .Q(
        DP_coeffs_ff_int[12]), .QN(n473) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_12_ ( .D(n930), .CK(clk), .RN(n1097), .Q(
        DP_coeffs_ff_int[11]), .QN(n472) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_13_ ( .D(n929), .CK(clk), .RN(n1097), .Q(
        DP_coeffs_ff_int[10]), .QN(n471) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_14_ ( .D(n928), .CK(clk), .RN(n1097), .Q(
        DP_coeffs_ff_int[9]), .QN(n470) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_15_ ( .D(n927), .CK(clk), .RN(n1097), .Q(
        DP_coeffs_ff_int[8]), .QN(n469) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_16_ ( .D(n926), .CK(clk), .RN(n1097), .Q(
        DP_coeffs_ff_int[7]), .QN(n468) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_17_ ( .D(n925), .CK(clk), .RN(n1097), .Q(
        DP_coeffs_ff_int[6]), .QN(n467) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_18_ ( .D(n924), .CK(clk), .RN(n1097), .Q(
        DP_coeffs_ff_int[5]), .QN(n466) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_19_ ( .D(n923), .CK(clk), .RN(n1097), .Q(
        DP_coeffs_ff_int[4]), .QN(n465) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_20_ ( .D(n922), .CK(clk), .RN(n1097), .Q(
        DP_coeffs_ff_int[3]), .QN(n464) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_21_ ( .D(n921), .CK(clk), .RN(n1097), .Q(
        DP_coeffs_ff_int[2]), .QN(n463) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_22_ ( .D(n920), .CK(clk), .RN(n1097), .Q(
        DP_coeffs_ff_int[1]), .QN(n462) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_23_ ( .D(n919), .CK(clk), .RN(n1097), .Q(
        DP_coeffs_ff_int[0]), .QN(n461) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_0_ ( .D(n918), .CK(clk), .RN(n1098), .Q(
        DP_coeffs_ff_int[47]), .QN(n460) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_1_ ( .D(n917), .CK(clk), .RN(n1098), .Q(
        DP_coeffs_ff_int[46]), .QN(n459) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_2_ ( .D(n916), .CK(clk), .RN(n1098), .Q(
        DP_coeffs_ff_int[45]), .QN(n458) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_3_ ( .D(n915), .CK(clk), .RN(n1098), .Q(
        DP_coeffs_ff_int[44]), .QN(n457) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_4_ ( .D(n914), .CK(clk), .RN(n1098), .Q(
        DP_coeffs_ff_int[43]), .QN(n456) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_5_ ( .D(n913), .CK(clk), .RN(n1098), .Q(
        DP_coeffs_ff_int[42]), .QN(n455) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_6_ ( .D(n912), .CK(clk), .RN(n1098), .Q(
        DP_coeffs_ff_int[41]), .QN(n454) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_7_ ( .D(n911), .CK(clk), .RN(n1098), .Q(
        DP_coeffs_ff_int[40]), .QN(n453) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_8_ ( .D(n910), .CK(clk), .RN(n1098), .Q(
        DP_coeffs_ff_int[39]), .QN(n452) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_9_ ( .D(n909), .CK(clk), .RN(n1098), .Q(
        DP_coeffs_ff_int[38]), .QN(n451) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_10_ ( .D(n908), .CK(clk), .RN(n1098), .Q(
        DP_coeffs_ff_int[37]), .QN(n450) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_11_ ( .D(n907), .CK(clk), .RN(n1098), .Q(
        DP_coeffs_ff_int[36]), .QN(n449) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_12_ ( .D(n906), .CK(clk), .RN(n1099), .Q(
        DP_coeffs_ff_int[35]), .QN(n448) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_13_ ( .D(n905), .CK(clk), .RN(n1099), .Q(
        DP_coeffs_ff_int[34]), .QN(n447) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_14_ ( .D(n904), .CK(clk), .RN(n1099), .Q(
        DP_coeffs_ff_int[33]), .QN(n446) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_15_ ( .D(n903), .CK(clk), .RN(n1099), .Q(
        DP_coeffs_ff_int[32]), .QN(n445) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_16_ ( .D(n902), .CK(clk), .RN(n1099), .Q(
        DP_coeffs_ff_int[31]), .QN(n444) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_17_ ( .D(n901), .CK(clk), .RN(n1099), .Q(
        DP_coeffs_ff_int[30]), .QN(n443) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_18_ ( .D(n900), .CK(clk), .RN(n1099), .Q(
        DP_coeffs_ff_int[29]), .QN(n442) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_19_ ( .D(n899), .CK(clk), .RN(n1099), .Q(
        DP_coeffs_ff_int[28]), .QN(n441) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_20_ ( .D(n898), .CK(clk), .RN(n1099), .Q(
        DP_coeffs_ff_int[27]), .QN(n440) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_21_ ( .D(n897), .CK(clk), .RN(n1099), .Q(
        DP_coeffs_ff_int[26]), .QN(n439) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_22_ ( .D(n896), .CK(clk), .RN(n1099), .Q(
        DP_coeffs_ff_int[25]), .QN(n438) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_23_ ( .D(n895), .CK(clk), .RN(n1099), .Q(
        DP_coeffs_ff_int[24]), .QN(n437) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_0_ ( .D(n894), .CK(clk), .RN(n1100), .Q(
        DP_coeffs_ff_int[71]), .QN(n436) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_1_ ( .D(n893), .CK(clk), .RN(n1100), .Q(
        DP_coeffs_ff_int[70]), .QN(n435) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_2_ ( .D(n892), .CK(clk), .RN(n1100), .Q(
        DP_coeffs_ff_int[69]), .QN(n434) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_3_ ( .D(n891), .CK(clk), .RN(n1100), .Q(
        DP_coeffs_ff_int[68]), .QN(n433) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_4_ ( .D(n890), .CK(clk), .RN(n1100), .Q(
        DP_coeffs_ff_int[67]), .QN(n432) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_5_ ( .D(n889), .CK(clk), .RN(n1100), .Q(
        DP_coeffs_ff_int[66]), .QN(n431) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_6_ ( .D(n888), .CK(clk), .RN(n1100), .Q(
        DP_coeffs_ff_int[65]), .QN(n430) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_7_ ( .D(n887), .CK(clk), .RN(n1100), .Q(
        DP_coeffs_ff_int[64]), .QN(n429) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_8_ ( .D(n886), .CK(clk), .RN(n1100), .Q(
        DP_coeffs_ff_int[63]), .QN(n428) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_9_ ( .D(n885), .CK(clk), .RN(n1100), .Q(
        DP_coeffs_ff_int[62]), .QN(n427) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_10_ ( .D(n884), .CK(clk), .RN(n1100), .Q(
        DP_coeffs_ff_int[61]), .QN(n426) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_11_ ( .D(n883), .CK(clk), .RN(n1100), .Q(
        DP_coeffs_ff_int[60]), .QN(n425) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_12_ ( .D(n882), .CK(clk), .RN(n1101), .Q(
        DP_coeffs_ff_int[59]), .QN(n424) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_13_ ( .D(n881), .CK(clk), .RN(n1101), .Q(
        DP_coeffs_ff_int[58]), .QN(n423) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_14_ ( .D(n880), .CK(clk), .RN(n1101), .Q(
        DP_coeffs_ff_int[57]), .QN(n422) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_15_ ( .D(n879), .CK(clk), .RN(n1101), .Q(
        DP_coeffs_ff_int[56]), .QN(n421) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_16_ ( .D(n878), .CK(clk), .RN(n1101), .Q(
        DP_coeffs_ff_int[55]), .QN(n420) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_17_ ( .D(n877), .CK(clk), .RN(n1101), .Q(
        DP_coeffs_ff_int[54]), .QN(n419) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_18_ ( .D(n876), .CK(clk), .RN(n1101), .Q(
        DP_coeffs_ff_int[53]), .QN(n418) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_19_ ( .D(n875), .CK(clk), .RN(n1101), .Q(
        DP_coeffs_ff_int[52]), .QN(n417) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_20_ ( .D(n874), .CK(clk), .RN(n1101), .Q(
        DP_coeffs_ff_int[51]), .QN(n416) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_21_ ( .D(n873), .CK(clk), .RN(n1101), .Q(
        DP_coeffs_ff_int[50]), .QN(n415) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_22_ ( .D(n872), .CK(clk), .RN(n1101), .Q(
        DP_coeffs_ff_int[49]), .QN(n414) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_23_ ( .D(n871), .CK(clk), .RN(n1101), .Q(
        DP_coeffs_ff_int[48]), .QN(n413) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_0_ ( .D(n870), .CK(clk), .RN(n1102), .Q(
        DP_coeffs_ff_int[95]), .QN(n412) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_1_ ( .D(n869), .CK(clk), .RN(n1102), .Q(
        DP_coeffs_ff_int[94]), .QN(n411) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_2_ ( .D(n868), .CK(clk), .RN(n1102), .Q(
        DP_coeffs_ff_int[93]), .QN(n410) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_3_ ( .D(n867), .CK(clk), .RN(n1102), .Q(
        DP_coeffs_ff_int[92]), .QN(n409) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_4_ ( .D(n866), .CK(clk), .RN(n1102), .Q(
        DP_coeffs_ff_int[91]), .QN(n408) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_5_ ( .D(n865), .CK(clk), .RN(n1102), .Q(
        DP_coeffs_ff_int[90]), .QN(n407) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_6_ ( .D(n864), .CK(clk), .RN(n1102), .Q(
        DP_coeffs_ff_int[89]), .QN(n406) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_7_ ( .D(n863), .CK(clk), .RN(n1102), .Q(
        DP_coeffs_ff_int[88]), .QN(n405) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_8_ ( .D(n862), .CK(clk), .RN(n1102), .Q(
        DP_coeffs_ff_int[87]), .QN(n404) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_9_ ( .D(n861), .CK(clk), .RN(n1102), .Q(
        DP_coeffs_ff_int[86]), .QN(n403) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_10_ ( .D(n860), .CK(clk), .RN(n1102), .Q(
        DP_coeffs_ff_int[85]), .QN(n402) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_11_ ( .D(n859), .CK(clk), .RN(n1102), .Q(
        DP_coeffs_ff_int[84]), .QN(n401) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_12_ ( .D(n858), .CK(clk), .RN(n1103), .Q(
        DP_coeffs_ff_int[83]), .QN(n400) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_13_ ( .D(n857), .CK(clk), .RN(n1103), .Q(
        DP_coeffs_ff_int[82]), .QN(n399) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_14_ ( .D(n856), .CK(clk), .RN(n1103), .Q(
        DP_coeffs_ff_int[81]), .QN(n398) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_15_ ( .D(n855), .CK(clk), .RN(n1103), .Q(
        DP_coeffs_ff_int[80]), .QN(n397) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_16_ ( .D(n854), .CK(clk), .RN(n1103), .Q(
        DP_coeffs_ff_int[79]), .QN(n396) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_17_ ( .D(n853), .CK(clk), .RN(n1103), .Q(
        DP_coeffs_ff_int[78]), .QN(n395) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_18_ ( .D(n852), .CK(clk), .RN(n1103), .Q(
        DP_coeffs_ff_int[77]), .QN(n394) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_19_ ( .D(n851), .CK(clk), .RN(n1103), .Q(
        DP_coeffs_ff_int[76]), .QN(n393) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_20_ ( .D(n850), .CK(clk), .RN(n1103), .Q(
        DP_coeffs_ff_int[75]), .QN(n392) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_21_ ( .D(n849), .CK(clk), .RN(n1103), .Q(
        DP_coeffs_ff_int[74]), .QN(n391) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_22_ ( .D(n848), .CK(clk), .RN(n1103), .Q(
        DP_coeffs_ff_int[73]), .QN(n390) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_23_ ( .D(n847), .CK(clk), .RN(n1103), .Q(
        DP_coeffs_ff_int[72]), .QN(n389) );
  DFFR_X1 CU_presentState_reg_1_ ( .D(n1034), .CK(clk), .RN(n1104), .Q(
        delayed_controls_0__1_) );
  DFFR_X1 DP_reg_sw1_Q_reg_0_ ( .D(n846), .CK(clk), .RN(n1104), .Q(DP_sw1_0_), 
        .QN(n1003) );
  DFFR_X1 DP_reg_pipe02_Q_reg_0_ ( .D(DP_sw1_0_), .CK(clk), .RN(n1104), .Q(
        DP_pipe02[0]) );
  DFFR_X1 DP_reg_ret1_Q_reg_0_ ( .D(DP_sw1_coeff_ret1[0]), .CK(clk), .RN(n1104), .Q(DP_ret1[0]) );
  DFFR_X1 DP_reg_ret1_Q_reg_1_ ( .D(DP_sw1_coeff_ret1[1]), .CK(clk), .RN(n1104), .Q(DP_ret1[1]) );
  DFFR_X1 DP_reg_ret1_Q_reg_2_ ( .D(DP_sw1_coeff_ret1[2]), .CK(clk), .RN(n1104), .Q(DP_ret1[2]) );
  DFFR_X1 DP_reg_ret1_Q_reg_3_ ( .D(DP_sw1_coeff_ret1[3]), .CK(clk), .RN(n1104), .Q(DP_ret1[3]) );
  DFFR_X1 DP_reg_ret1_Q_reg_4_ ( .D(DP_sw1_coeff_ret1[4]), .CK(clk), .RN(n1104), .Q(DP_ret1[4]) );
  DFFR_X1 DP_reg_ret1_Q_reg_5_ ( .D(DP_sw1_coeff_ret1[5]), .CK(clk), .RN(n1104), .Q(DP_ret1[5]) );
  DFFR_X1 DP_reg_ret1_Q_reg_6_ ( .D(DP_sw1_coeff_ret1[6]), .CK(clk), .RN(n1104), .Q(DP_ret1[6]) );
  DFFR_X1 DP_reg_ret1_Q_reg_7_ ( .D(DP_sw1_coeff_ret1[7]), .CK(clk), .RN(n1104), .Q(DP_ret1[7]) );
  DFFR_X1 DP_reg_ret1_Q_reg_8_ ( .D(DP_sw1_coeff_ret1[8]), .CK(clk), .RN(n1104), .Q(DP_ret1[8]) );
  DFFR_X1 DP_reg_ret1_Q_reg_9_ ( .D(DP_sw1_coeff_ret1[9]), .CK(clk), .RN(n1105), .Q(DP_ret1[9]) );
  DFFR_X1 DP_reg_ret1_Q_reg_10_ ( .D(DP_sw1_coeff_ret1[10]), .CK(clk), .RN(
        n1105), .Q(DP_ret1[10]) );
  DFFR_X1 DP_reg_ret1_Q_reg_11_ ( .D(DP_sw1_coeff_ret1[11]), .CK(clk), .RN(
        n1105), .Q(DP_ret1[11]) );
  DFFR_X1 DP_reg_ret1_Q_reg_12_ ( .D(DP_sw1_coeff_ret1[12]), .CK(clk), .RN(
        n1105), .Q(DP_ret1[12]) );
  DFFR_X1 DP_reg_ret1_Q_reg_13_ ( .D(DP_sw1_coeff_ret1[13]), .CK(clk), .RN(
        n1105), .Q(DP_ret1[13]) );
  DFFR_X1 DP_reg_ret1_Q_reg_14_ ( .D(DP_sw1_coeff_ret1[14]), .CK(clk), .RN(
        n1105), .Q(DP_ret1[14]) );
  DFFR_X1 DP_reg_ret1_Q_reg_15_ ( .D(DP_sw1_coeff_ret1[15]), .CK(clk), .RN(
        n1105), .Q(DP_ret1[15]) );
  DFFR_X1 DP_reg_ret1_Q_reg_16_ ( .D(DP_sw1_coeff_ret1[16]), .CK(clk), .RN(
        n1105), .Q(DP_ret1[16]) );
  DFFR_X1 DP_reg_ret1_Q_reg_17_ ( .D(DP_sw1_coeff_ret1[17]), .CK(clk), .RN(
        n1105), .Q(DP_ret1[17]) );
  DFFR_X1 DP_reg_ret1_Q_reg_18_ ( .D(DP_sw1_coeff_ret1[18]), .CK(clk), .RN(
        n1105), .Q(DP_ret1[18]) );
  DFFR_X1 DP_reg_ret1_Q_reg_19_ ( .D(DP_sw1_coeff_ret1[19]), .CK(clk), .RN(
        n1105), .Q(DP_ret1[19]) );
  DFFR_X1 DP_reg_ret1_Q_reg_20_ ( .D(DP_sw1_coeff_ret1[20]), .CK(clk), .RN(
        n1105), .Q(DP_ret1[20]) );
  DFFR_X1 DP_reg_ret1_Q_reg_21_ ( .D(DP_sw1_coeff_ret1[21]), .CK(clk), .RN(
        n1106), .Q(DP_ret1[21]) );
  DFFR_X1 DP_reg_ret1_Q_reg_22_ ( .D(DP_sw1_coeff_ret1[22]), .CK(clk), .RN(
        n1106), .Q(DP_ret1[22]) );
  DFFR_X1 DP_reg_ret1_Q_reg_23_ ( .D(DP_sw1_coeff_ret1[23]), .CK(clk), .RN(
        n1106), .Q(DP_ret1[23]) );
  DFFR_X1 DP_reg_sw0_Q_reg_0_ ( .D(n820), .CK(clk), .RN(n1106), .Q(DP_sw0_0_), 
        .QN(n1005) );
  DFFR_X1 DP_reg_pipe01_Q_reg_0_ ( .D(DP_sw0_0_), .CK(clk), .RN(n1106), .Q(
        DP_pipe01[0]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_0_ ( .D(DP_w_0_), .CK(clk), .RN(n1106), .Q(
        DP_pipe00[0]) );
  DFFR_X1 DP_reg_sw0_Q_reg_1_ ( .D(n817), .CK(clk), .RN(n1106), .Q(DP_sw0_1_)
         );
  DFFR_X1 DP_reg_sw1_Q_reg_1_ ( .D(n816), .CK(clk), .RN(n1106), .Q(DP_sw1_1_), 
        .QN(n1006) );
  DFFR_X1 DP_reg_pipe02_Q_reg_1_ ( .D(DP_sw1_1_), .CK(clk), .RN(n1106), .Q(
        DP_pipe02[1]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_1_ ( .D(DP_sw0_1_), .CK(clk), .RN(n1106), .Q(
        DP_pipe01[1]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_1_ ( .D(DP_w_1_), .CK(clk), .RN(n1106), .Q(
        DP_pipe00[1]) );
  DFFR_X1 DP_reg_sw0_Q_reg_2_ ( .D(n812), .CK(clk), .RN(n1106), .Q(DP_sw0_2_)
         );
  DFFR_X1 DP_reg_sw1_Q_reg_2_ ( .D(n811), .CK(clk), .RN(n1107), .Q(DP_sw1_2_), 
        .QN(n1007) );
  DFFR_X1 DP_reg_pipe02_Q_reg_2_ ( .D(DP_sw1_2_), .CK(clk), .RN(n1107), .Q(
        DP_pipe02[2]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_2_ ( .D(DP_sw0_2_), .CK(clk), .RN(n1107), .Q(
        DP_pipe01[2]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_2_ ( .D(DP_w_2_), .CK(clk), .RN(n1107), .Q(
        DP_pipe00[2]) );
  DFFR_X1 DP_reg_sw0_Q_reg_3_ ( .D(n807), .CK(clk), .RN(n1107), .Q(DP_sw0_3_)
         );
  DFFR_X1 DP_reg_sw1_Q_reg_3_ ( .D(n806), .CK(clk), .RN(n1107), .Q(DP_sw1_3_), 
        .QN(n1008) );
  DFFR_X1 DP_reg_pipe02_Q_reg_3_ ( .D(DP_sw1_3_), .CK(clk), .RN(n1107), .Q(
        DP_pipe02[3]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_3_ ( .D(DP_sw0_3_), .CK(clk), .RN(n1107), .Q(
        DP_pipe01[3]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_3_ ( .D(DP_w_3_), .CK(clk), .RN(n1107), .Q(
        DP_pipe00[3]) );
  DFFR_X1 DP_reg_sw0_Q_reg_4_ ( .D(n802), .CK(clk), .RN(n1107), .Q(DP_sw0_4_)
         );
  DFFR_X1 DP_reg_sw1_Q_reg_4_ ( .D(n801), .CK(clk), .RN(n1107), .Q(DP_sw1_4_), 
        .QN(n1009) );
  DFFR_X1 DP_reg_pipe02_Q_reg_4_ ( .D(DP_sw1_4_), .CK(clk), .RN(n1107), .Q(
        DP_pipe02[4]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_4_ ( .D(DP_sw0_4_), .CK(clk), .RN(n1108), .Q(
        DP_pipe01[4]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_4_ ( .D(DP_w_4_), .CK(clk), .RN(n1108), .Q(
        DP_pipe00[4]) );
  DFFR_X1 DP_reg_sw0_Q_reg_5_ ( .D(n797), .CK(clk), .RN(n1108), .Q(DP_sw0_5_)
         );
  DFFR_X1 DP_reg_sw1_Q_reg_5_ ( .D(n796), .CK(clk), .RN(n1108), .Q(DP_sw1_5_), 
        .QN(n1010) );
  DFFR_X1 DP_reg_pipe02_Q_reg_5_ ( .D(DP_sw1_5_), .CK(clk), .RN(n1108), .Q(
        DP_pipe02[5]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_5_ ( .D(DP_sw0_5_), .CK(clk), .RN(n1108), .Q(
        DP_pipe01[5]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_5_ ( .D(DP_w_5_), .CK(clk), .RN(n1108), .Q(
        DP_pipe00[5]) );
  DFFR_X1 DP_reg_sw0_Q_reg_6_ ( .D(n792), .CK(clk), .RN(n1108), .Q(DP_sw0_6_)
         );
  DFFR_X1 DP_reg_sw1_Q_reg_6_ ( .D(n791), .CK(clk), .RN(n1108), .Q(DP_sw1_6_), 
        .QN(n1011) );
  DFFR_X1 DP_reg_pipe02_Q_reg_6_ ( .D(DP_sw1_6_), .CK(clk), .RN(n1108), .Q(
        DP_pipe02[6]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_6_ ( .D(DP_sw0_6_), .CK(clk), .RN(n1108), .Q(
        DP_pipe01[6]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_6_ ( .D(DP_w_6_), .CK(clk), .RN(n1108), .Q(
        DP_pipe00[6]) );
  DFFR_X1 DP_reg_sw0_Q_reg_7_ ( .D(n787), .CK(clk), .RN(n1109), .Q(DP_sw0_7_)
         );
  DFFR_X1 DP_reg_sw1_Q_reg_7_ ( .D(n786), .CK(clk), .RN(n1109), .Q(DP_sw1_7_), 
        .QN(n1012) );
  DFFR_X1 DP_reg_pipe02_Q_reg_7_ ( .D(DP_sw1_7_), .CK(clk), .RN(n1109), .Q(
        DP_pipe02[7]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_7_ ( .D(DP_sw0_7_), .CK(clk), .RN(n1109), .Q(
        DP_pipe01[7]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_7_ ( .D(DP_w_7_), .CK(clk), .RN(n1109), .Q(
        DP_pipe00[7]) );
  DFFR_X1 DP_reg_sw0_Q_reg_8_ ( .D(n782), .CK(clk), .RN(n1109), .Q(DP_sw0_8_)
         );
  DFFR_X1 DP_reg_sw1_Q_reg_8_ ( .D(n781), .CK(clk), .RN(n1109), .Q(DP_sw1_8_), 
        .QN(n1013) );
  DFFR_X1 DP_reg_pipe02_Q_reg_8_ ( .D(DP_sw1_8_), .CK(clk), .RN(n1109), .Q(
        DP_pipe02[8]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_8_ ( .D(DP_sw0_8_), .CK(clk), .RN(n1109), .Q(
        DP_pipe01[8]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_8_ ( .D(DP_w_8_), .CK(clk), .RN(n1109), .Q(
        DP_pipe00[8]) );
  DFFR_X1 DP_reg_sw0_Q_reg_9_ ( .D(n777), .CK(clk), .RN(n1109), .Q(DP_sw0_9_)
         );
  DFFR_X1 DP_reg_sw1_Q_reg_9_ ( .D(n776), .CK(clk), .RN(n1109), .Q(DP_sw1_9_), 
        .QN(n1014) );
  DFFR_X1 DP_reg_pipe02_Q_reg_9_ ( .D(DP_sw1_9_), .CK(clk), .RN(n1110), .Q(
        DP_pipe02[9]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_9_ ( .D(DP_sw0_9_), .CK(clk), .RN(n1110), .Q(
        DP_pipe01[9]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_9_ ( .D(DP_w_9_), .CK(clk), .RN(n1110), .Q(
        DP_pipe00[9]) );
  DFFR_X1 DP_reg_sw0_Q_reg_10_ ( .D(n772), .CK(clk), .RN(n1110), .Q(DP_sw0_10_) );
  DFFR_X1 DP_reg_sw1_Q_reg_10_ ( .D(n771), .CK(clk), .RN(n1110), .Q(DP_sw1_10_), .QN(n1015) );
  DFFR_X1 DP_reg_pipe02_Q_reg_10_ ( .D(DP_sw1_10_), .CK(clk), .RN(n1110), .Q(
        DP_pipe02[10]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_10_ ( .D(DP_sw0_10_), .CK(clk), .RN(n1110), .Q(
        DP_pipe01[10]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_10_ ( .D(DP_w_10_), .CK(clk), .RN(n1110), .Q(
        DP_pipe00[10]) );
  DFFR_X1 DP_reg_sw0_Q_reg_11_ ( .D(n767), .CK(clk), .RN(n1110), .Q(DP_sw0_11_) );
  DFFR_X1 DP_reg_sw1_Q_reg_11_ ( .D(n766), .CK(clk), .RN(n1110), .Q(DP_sw1_11_), .QN(n1016) );
  DFFR_X1 DP_reg_pipe02_Q_reg_11_ ( .D(DP_sw1_11_), .CK(clk), .RN(n1110), .Q(
        DP_pipe02[11]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_11_ ( .D(DP_sw0_11_), .CK(clk), .RN(n1110), .Q(
        DP_pipe01[11]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_11_ ( .D(DP_w_11_), .CK(clk), .RN(n1111), .Q(
        DP_pipe00[11]) );
  DFFR_X1 DP_reg_sw0_Q_reg_12_ ( .D(n762), .CK(clk), .RN(n1111), .Q(DP_sw0_12_) );
  DFFR_X1 DP_reg_sw1_Q_reg_12_ ( .D(n761), .CK(clk), .RN(n1111), .Q(DP_sw1_12_), .QN(n1017) );
  DFFR_X1 DP_reg_pipe02_Q_reg_12_ ( .D(DP_sw1_12_), .CK(clk), .RN(n1111), .Q(
        DP_pipe02[12]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_12_ ( .D(DP_sw0_12_), .CK(clk), .RN(n1111), .Q(
        DP_pipe01[12]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_12_ ( .D(DP_w_12_), .CK(clk), .RN(n1111), .Q(
        DP_pipe00[12]) );
  DFFR_X1 DP_reg_sw0_Q_reg_13_ ( .D(n757), .CK(clk), .RN(n1111), .Q(DP_sw0_13_) );
  DFFR_X1 DP_reg_sw1_Q_reg_13_ ( .D(n756), .CK(clk), .RN(n1111), .Q(DP_sw1_13_), .QN(n1018) );
  DFFR_X1 DP_reg_pipe02_Q_reg_13_ ( .D(DP_sw1_13_), .CK(clk), .RN(n1111), .Q(
        DP_pipe02[13]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_13_ ( .D(DP_sw0_13_), .CK(clk), .RN(n1111), .Q(
        DP_pipe01[13]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_13_ ( .D(DP_w_13_), .CK(clk), .RN(n1111), .Q(
        DP_pipe00[13]) );
  DFFR_X1 DP_reg_sw0_Q_reg_14_ ( .D(n752), .CK(clk), .RN(n1111), .Q(DP_sw0_14_) );
  DFFR_X1 DP_reg_sw1_Q_reg_14_ ( .D(n751), .CK(clk), .RN(n1112), .Q(DP_sw1_14_), .QN(n1019) );
  DFFR_X1 DP_reg_pipe02_Q_reg_14_ ( .D(DP_sw1_14_), .CK(clk), .RN(n1112), .Q(
        DP_pipe02[14]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_14_ ( .D(DP_sw0_14_), .CK(clk), .RN(n1112), .Q(
        DP_pipe01[14]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_14_ ( .D(DP_w_14_), .CK(clk), .RN(n1112), .Q(
        DP_pipe00[14]) );
  DFFR_X1 DP_reg_sw0_Q_reg_15_ ( .D(n747), .CK(clk), .RN(n1112), .Q(DP_sw0_15_) );
  DFFR_X1 DP_reg_sw1_Q_reg_15_ ( .D(n746), .CK(clk), .RN(n1112), .Q(DP_sw1_15_), .QN(n1020) );
  DFFR_X1 DP_reg_pipe02_Q_reg_15_ ( .D(DP_sw1_15_), .CK(clk), .RN(n1112), .Q(
        DP_pipe02[15]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_15_ ( .D(DP_sw0_15_), .CK(clk), .RN(n1112), .Q(
        DP_pipe01[15]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_15_ ( .D(DP_w_15_), .CK(clk), .RN(n1112), .Q(
        DP_pipe00[15]) );
  DFFR_X1 DP_reg_sw0_Q_reg_16_ ( .D(n742), .CK(clk), .RN(n1112), .Q(DP_sw0_16_) );
  DFFR_X1 DP_reg_sw1_Q_reg_16_ ( .D(n741), .CK(clk), .RN(n1112), .Q(DP_sw1_16_), .QN(n1021) );
  DFFR_X1 DP_reg_pipe02_Q_reg_16_ ( .D(DP_sw1_16_), .CK(clk), .RN(n1112), .Q(
        DP_pipe02[16]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_16_ ( .D(DP_sw0_16_), .CK(clk), .RN(n1113), .Q(
        DP_pipe01[16]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_16_ ( .D(DP_w_16_), .CK(clk), .RN(n1113), .Q(
        DP_pipe00[16]) );
  DFFR_X1 DP_reg_sw0_Q_reg_17_ ( .D(n737), .CK(clk), .RN(n1113), .Q(DP_sw0_17_) );
  DFFR_X1 DP_reg_sw1_Q_reg_17_ ( .D(n736), .CK(clk), .RN(n1113), .Q(DP_sw1_17_), .QN(n1022) );
  DFFR_X1 DP_reg_pipe02_Q_reg_17_ ( .D(DP_sw1_17_), .CK(clk), .RN(n1113), .Q(
        DP_pipe02[17]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_17_ ( .D(DP_sw0_17_), .CK(clk), .RN(n1113), .Q(
        DP_pipe01[17]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_17_ ( .D(DP_w_17_), .CK(clk), .RN(n1113), .Q(
        DP_pipe00[17]) );
  DFFR_X1 DP_reg_sw0_Q_reg_18_ ( .D(n732), .CK(clk), .RN(n1113), .Q(DP_sw0_18_) );
  DFFR_X1 DP_reg_sw1_Q_reg_18_ ( .D(n731), .CK(clk), .RN(n1113), .Q(DP_sw1_18_), .QN(n1023) );
  DFFR_X1 DP_reg_pipe02_Q_reg_18_ ( .D(DP_sw1_18_), .CK(clk), .RN(n1113), .Q(
        DP_pipe02[18]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_18_ ( .D(DP_sw0_18_), .CK(clk), .RN(n1113), .Q(
        DP_pipe01[18]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_18_ ( .D(DP_w_18_), .CK(clk), .RN(n1113), .Q(
        DP_pipe00[18]) );
  DFFR_X1 DP_reg_sw0_Q_reg_19_ ( .D(n727), .CK(clk), .RN(n1114), .Q(DP_sw0_19_) );
  DFFR_X1 DP_reg_sw1_Q_reg_19_ ( .D(n726), .CK(clk), .RN(n1114), .Q(DP_sw1_19_), .QN(n1024) );
  DFFR_X1 DP_reg_pipe02_Q_reg_19_ ( .D(DP_sw1_19_), .CK(clk), .RN(n1114), .Q(
        DP_pipe02[19]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_19_ ( .D(DP_sw0_19_), .CK(clk), .RN(n1114), .Q(
        DP_pipe01[19]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_19_ ( .D(DP_w_19_), .CK(clk), .RN(n1114), .Q(
        DP_pipe00[19]) );
  DFFR_X1 DP_reg_sw0_Q_reg_20_ ( .D(n722), .CK(clk), .RN(n1114), .Q(DP_sw0_20_) );
  DFFR_X1 DP_reg_sw1_Q_reg_20_ ( .D(n721), .CK(clk), .RN(n1114), .Q(DP_sw1_20_), .QN(n1025) );
  DFFR_X1 DP_reg_pipe02_Q_reg_20_ ( .D(DP_sw1_20_), .CK(clk), .RN(n1114), .Q(
        DP_pipe02[20]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_20_ ( .D(DP_sw0_20_), .CK(clk), .RN(n1114), .Q(
        DP_pipe01[20]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_20_ ( .D(DP_w_20_), .CK(clk), .RN(n1114), .Q(
        DP_pipe00[20]) );
  DFFR_X1 DP_reg_sw0_Q_reg_21_ ( .D(n717), .CK(clk), .RN(n1114), .Q(DP_sw0_21_) );
  DFFR_X1 DP_reg_sw1_Q_reg_21_ ( .D(n716), .CK(clk), .RN(n1114), .Q(DP_sw1_21_), .QN(n1026) );
  DFFR_X1 DP_reg_pipe02_Q_reg_21_ ( .D(DP_sw1_21_), .CK(clk), .RN(n1115), .Q(
        DP_pipe02[21]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_21_ ( .D(DP_sw0_21_), .CK(clk), .RN(n1115), .Q(
        DP_pipe01[21]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_21_ ( .D(DP_w_21_), .CK(clk), .RN(n1115), .Q(
        DP_pipe00[21]) );
  DFFR_X1 DP_reg_sw0_Q_reg_22_ ( .D(n712), .CK(clk), .RN(n1115), .Q(DP_sw0_22_) );
  DFFR_X1 DP_reg_sw1_Q_reg_22_ ( .D(n711), .CK(clk), .RN(n1115), .Q(DP_sw1_22_), .QN(n1027) );
  DFFR_X1 DP_reg_pipe02_Q_reg_22_ ( .D(DP_sw1_22_), .CK(clk), .RN(n1115), .Q(
        DP_pipe02[22]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_22_ ( .D(DP_sw0_22_), .CK(clk), .RN(n1115), .Q(
        DP_pipe01[22]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_22_ ( .D(DP_w_22_), .CK(clk), .RN(n1115), .Q(
        DP_pipe00[22]) );
  DFFR_X1 DP_reg_sw0_Q_reg_23_ ( .D(n707), .CK(clk), .RN(n1115), .Q(DP_sw0_23_) );
  DFFR_X1 DP_reg_sw1_Q_reg_23_ ( .D(n706), .CK(clk), .RN(n1115), .Q(DP_sw1_23_), .QN(n1004) );
  DFFR_X1 DP_reg_pipe02_Q_reg_23_ ( .D(DP_sw1_23_), .CK(clk), .RN(n1115), .Q(
        DP_pipe02[23]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_0_ ( .D(DP_pipe0_coeff_pipe02[0]), .CK(clk), 
        .RN(n1115), .Q(DP_pipe12[0]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_1_ ( .D(DP_pipe0_coeff_pipe02[1]), .CK(clk), 
        .RN(n1116), .Q(DP_pipe12[1]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_2_ ( .D(DP_pipe0_coeff_pipe02[2]), .CK(clk), 
        .RN(n1116), .Q(DP_pipe12[2]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_3_ ( .D(DP_pipe0_coeff_pipe02[3]), .CK(clk), 
        .RN(n1116), .Q(DP_pipe12[3]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_4_ ( .D(DP_pipe0_coeff_pipe02[4]), .CK(clk), 
        .RN(n1116), .Q(DP_pipe12[4]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_5_ ( .D(DP_pipe0_coeff_pipe02[5]), .CK(clk), 
        .RN(n1116), .Q(DP_pipe12[5]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_6_ ( .D(DP_pipe0_coeff_pipe02[6]), .CK(clk), 
        .RN(n1116), .Q(DP_pipe12[6]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_7_ ( .D(DP_pipe0_coeff_pipe02[7]), .CK(clk), 
        .RN(n1116), .Q(DP_pipe12[7]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_8_ ( .D(DP_pipe0_coeff_pipe02[8]), .CK(clk), 
        .RN(n1116), .Q(DP_pipe12[8]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_9_ ( .D(DP_pipe0_coeff_pipe02[9]), .CK(clk), 
        .RN(n1116), .Q(DP_pipe12[9]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_10_ ( .D(DP_pipe0_coeff_pipe02[10]), .CK(clk), 
        .RN(n1116), .Q(DP_pipe12[10]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_11_ ( .D(DP_pipe0_coeff_pipe02[11]), .CK(clk), 
        .RN(n1116), .Q(DP_pipe12[11]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_12_ ( .D(DP_pipe0_coeff_pipe02[12]), .CK(clk), 
        .RN(n1116), .Q(DP_pipe12[12]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_13_ ( .D(DP_pipe0_coeff_pipe02[13]), .CK(clk), 
        .RN(n1117), .Q(DP_pipe12[13]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_14_ ( .D(DP_pipe0_coeff_pipe02[14]), .CK(clk), 
        .RN(n1117), .Q(DP_pipe12[14]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_15_ ( .D(DP_pipe0_coeff_pipe02[15]), .CK(clk), 
        .RN(n1117), .Q(DP_pipe12[15]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_16_ ( .D(DP_pipe0_coeff_pipe02[16]), .CK(clk), 
        .RN(n1117), .Q(DP_pipe12[16]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_17_ ( .D(DP_pipe0_coeff_pipe02[17]), .CK(clk), 
        .RN(n1117), .Q(DP_pipe12[17]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_18_ ( .D(DP_pipe0_coeff_pipe02[18]), .CK(clk), 
        .RN(n1117), .Q(DP_pipe12[18]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_19_ ( .D(DP_pipe0_coeff_pipe02[19]), .CK(clk), 
        .RN(n1117), .Q(DP_pipe12[19]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_20_ ( .D(DP_pipe0_coeff_pipe02[20]), .CK(clk), 
        .RN(n1117), .Q(DP_pipe12[20]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_21_ ( .D(DP_pipe0_coeff_pipe02[21]), .CK(clk), 
        .RN(n1117), .Q(DP_pipe12[21]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_22_ ( .D(DP_pipe0_coeff_pipe02[22]), .CK(clk), 
        .RN(n1117), .Q(DP_pipe12[22]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_23_ ( .D(DP_pipe0_coeff_pipe02[23]), .CK(clk), 
        .RN(n1117), .Q(DP_pipe12[23]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_23_ ( .D(DP_sw0_23_), .CK(clk), .RN(n1117), .Q(
        DP_pipe01[23]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_0_ ( .D(DP_pipe0_coeff_pipe01[0]), .CK(clk), 
        .RN(n1118), .Q(DP_pipe11[0]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_1_ ( .D(DP_pipe0_coeff_pipe01[1]), .CK(clk), 
        .RN(n1118), .Q(DP_pipe11[1]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_2_ ( .D(DP_pipe0_coeff_pipe01[2]), .CK(clk), 
        .RN(n1118), .Q(DP_pipe11[2]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_3_ ( .D(DP_pipe0_coeff_pipe01[3]), .CK(clk), 
        .RN(n1118), .Q(DP_pipe11[3]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_4_ ( .D(DP_pipe0_coeff_pipe01[4]), .CK(clk), 
        .RN(n1118), .Q(DP_pipe11[4]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_5_ ( .D(DP_pipe0_coeff_pipe01[5]), .CK(clk), 
        .RN(n1118), .Q(DP_pipe11[5]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_6_ ( .D(DP_pipe0_coeff_pipe01[6]), .CK(clk), 
        .RN(n1118), .Q(DP_pipe11[6]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_7_ ( .D(DP_pipe0_coeff_pipe01[7]), .CK(clk), 
        .RN(n1118), .Q(DP_pipe11[7]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_8_ ( .D(DP_pipe0_coeff_pipe01[8]), .CK(clk), 
        .RN(n1118), .Q(DP_pipe11[8]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_9_ ( .D(DP_pipe0_coeff_pipe01[9]), .CK(clk), 
        .RN(n1118), .Q(DP_pipe11[9]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_10_ ( .D(DP_pipe0_coeff_pipe01[10]), .CK(clk), 
        .RN(n1118), .Q(DP_pipe11[10]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_11_ ( .D(DP_pipe0_coeff_pipe01[11]), .CK(clk), 
        .RN(n1118), .Q(DP_pipe11[11]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_12_ ( .D(DP_pipe0_coeff_pipe01[12]), .CK(clk), 
        .RN(n1119), .Q(DP_pipe11[12]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_13_ ( .D(DP_pipe0_coeff_pipe01[13]), .CK(clk), 
        .RN(n1119), .Q(DP_pipe11[13]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_14_ ( .D(DP_pipe0_coeff_pipe01[14]), .CK(clk), 
        .RN(n1119), .Q(DP_pipe11[14]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_15_ ( .D(DP_pipe0_coeff_pipe01[15]), .CK(clk), 
        .RN(n1119), .Q(DP_pipe11[15]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_16_ ( .D(DP_pipe0_coeff_pipe01[16]), .CK(clk), 
        .RN(n1119), .Q(DP_pipe11[16]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_17_ ( .D(DP_pipe0_coeff_pipe01[17]), .CK(clk), 
        .RN(n1119), .Q(DP_pipe11[17]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_18_ ( .D(DP_pipe0_coeff_pipe01[18]), .CK(clk), 
        .RN(n1119), .Q(DP_pipe11[18]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_19_ ( .D(DP_pipe0_coeff_pipe01[19]), .CK(clk), 
        .RN(n1119), .Q(DP_pipe11[19]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_20_ ( .D(DP_pipe0_coeff_pipe01[20]), .CK(clk), 
        .RN(n1119), .Q(DP_pipe11[20]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_21_ ( .D(DP_pipe0_coeff_pipe01[21]), .CK(clk), 
        .RN(n1119), .Q(DP_pipe11[21]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_22_ ( .D(DP_pipe0_coeff_pipe01[22]), .CK(clk), 
        .RN(n1119), .Q(DP_pipe11[22]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_23_ ( .D(DP_pipe0_coeff_pipe01[23]), .CK(clk), 
        .RN(n1119), .Q(DP_pipe11[23]) );
  DFFR_X1 DP_reg_ret0_Q_reg_0_ ( .D(DP_sw0_coeff_ret0[0]), .CK(clk), .RN(n1120), .Q(DP_ret0[0]) );
  DFFR_X1 DP_reg_ret0_Q_reg_1_ ( .D(DP_sw0_coeff_ret0[1]), .CK(clk), .RN(n1120), .Q(DP_ret0[1]) );
  DFFR_X1 DP_reg_ret0_Q_reg_2_ ( .D(DP_sw0_coeff_ret0[2]), .CK(clk), .RN(n1120), .Q(DP_ret0[2]) );
  DFFR_X1 DP_reg_ret0_Q_reg_3_ ( .D(DP_sw0_coeff_ret0[3]), .CK(clk), .RN(n1120), .Q(DP_ret0[3]) );
  DFFR_X1 DP_reg_ret0_Q_reg_4_ ( .D(DP_sw0_coeff_ret0[4]), .CK(clk), .RN(n1120), .Q(DP_ret0[4]) );
  DFFR_X1 DP_reg_ret0_Q_reg_5_ ( .D(DP_sw0_coeff_ret0[5]), .CK(clk), .RN(n1120), .Q(DP_ret0[5]) );
  DFFR_X1 DP_reg_ret0_Q_reg_6_ ( .D(DP_sw0_coeff_ret0[6]), .CK(clk), .RN(n1120), .Q(DP_ret0[6]) );
  DFFR_X1 DP_reg_ret0_Q_reg_7_ ( .D(DP_sw0_coeff_ret0[7]), .CK(clk), .RN(n1120), .Q(DP_ret0[7]) );
  DFFR_X1 DP_reg_ret0_Q_reg_8_ ( .D(DP_sw0_coeff_ret0[8]), .CK(clk), .RN(n1120), .Q(DP_ret0[8]) );
  DFFR_X1 DP_reg_ret0_Q_reg_9_ ( .D(DP_sw0_coeff_ret0[9]), .CK(clk), .RN(n1120), .Q(DP_ret0[9]) );
  DFFR_X1 DP_reg_ret0_Q_reg_10_ ( .D(DP_sw0_coeff_ret0[10]), .CK(clk), .RN(
        n1120), .Q(DP_ret0[10]) );
  DFFR_X1 DP_reg_ret0_Q_reg_11_ ( .D(DP_sw0_coeff_ret0[11]), .CK(clk), .RN(
        n1120), .Q(DP_ret0[11]) );
  DFFR_X1 DP_reg_ret0_Q_reg_12_ ( .D(DP_sw0_coeff_ret0[12]), .CK(clk), .RN(
        n1121), .Q(DP_ret0[12]) );
  DFFR_X1 DP_reg_ret0_Q_reg_13_ ( .D(DP_sw0_coeff_ret0[13]), .CK(clk), .RN(
        n1121), .Q(DP_ret0[13]) );
  DFFR_X1 DP_reg_ret0_Q_reg_14_ ( .D(DP_sw0_coeff_ret0[14]), .CK(clk), .RN(
        n1121), .Q(DP_ret0[14]) );
  DFFR_X1 DP_reg_ret0_Q_reg_15_ ( .D(DP_sw0_coeff_ret0[15]), .CK(clk), .RN(
        n1121), .Q(DP_ret0[15]) );
  DFFR_X1 DP_reg_ret0_Q_reg_16_ ( .D(DP_sw0_coeff_ret0[16]), .CK(clk), .RN(
        n1121), .Q(DP_ret0[16]) );
  DFFR_X1 DP_reg_ret0_Q_reg_17_ ( .D(DP_sw0_coeff_ret0[17]), .CK(clk), .RN(
        n1121), .Q(DP_ret0[17]) );
  DFFR_X1 DP_reg_ret0_Q_reg_18_ ( .D(DP_sw0_coeff_ret0[18]), .CK(clk), .RN(
        n1121), .Q(DP_ret0[18]) );
  DFFR_X1 DP_reg_ret0_Q_reg_19_ ( .D(DP_sw0_coeff_ret0[19]), .CK(clk), .RN(
        n1121), .Q(DP_ret0[19]) );
  DFFR_X1 DP_reg_ret0_Q_reg_20_ ( .D(DP_sw0_coeff_ret0[20]), .CK(clk), .RN(
        n1121), .Q(DP_ret0[20]) );
  DFFR_X1 DP_reg_ret0_Q_reg_21_ ( .D(DP_sw0_coeff_ret0[21]), .CK(clk), .RN(
        n1121), .Q(DP_ret0[21]) );
  DFFR_X1 DP_reg_ret0_Q_reg_22_ ( .D(DP_sw0_coeff_ret0[22]), .CK(clk), .RN(
        n1121), .Q(DP_ret0[22]) );
  DFFR_X1 DP_reg_ret0_Q_reg_23_ ( .D(DP_sw0_coeff_ret0[23]), .CK(clk), .RN(
        n1121), .Q(DP_ret0[23]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_23_ ( .D(DP_w_23_), .CK(clk), .RN(n1122), .Q(
        DP_pipe00[23]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_0_ ( .D(DP_pipe0_coeff_pipe00[0]), .CK(clk), 
        .RN(n1122), .Q(DP_pipe10[0]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_1_ ( .D(DP_pipe0_coeff_pipe00[1]), .CK(clk), 
        .RN(n1122), .Q(DP_pipe10[1]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_2_ ( .D(DP_pipe0_coeff_pipe00[2]), .CK(clk), 
        .RN(n1122), .Q(DP_pipe10[2]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_3_ ( .D(DP_pipe0_coeff_pipe00[3]), .CK(clk), 
        .RN(n1122), .Q(DP_pipe10[3]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_4_ ( .D(DP_pipe0_coeff_pipe00[4]), .CK(clk), 
        .RN(n1122), .Q(DP_pipe10[4]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_5_ ( .D(DP_pipe0_coeff_pipe00[5]), .CK(clk), 
        .RN(n1122), .Q(DP_pipe10[5]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_6_ ( .D(DP_pipe0_coeff_pipe00[6]), .CK(clk), 
        .RN(n1122), .Q(DP_pipe10[6]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_7_ ( .D(DP_pipe0_coeff_pipe00[7]), .CK(clk), 
        .RN(n1122), .Q(DP_pipe10[7]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_8_ ( .D(DP_pipe0_coeff_pipe00[8]), .CK(clk), 
        .RN(n1122), .Q(DP_pipe10[8]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_9_ ( .D(DP_pipe0_coeff_pipe00[9]), .CK(clk), 
        .RN(n1122), .Q(DP_pipe10[9]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_10_ ( .D(DP_pipe0_coeff_pipe00[10]), .CK(clk), 
        .RN(n1122), .Q(DP_pipe10[10]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_11_ ( .D(DP_pipe0_coeff_pipe00[11]), .CK(clk), 
        .RN(n1123), .Q(DP_pipe10[11]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_12_ ( .D(DP_pipe0_coeff_pipe00[12]), .CK(clk), 
        .RN(n1123), .Q(DP_pipe10[12]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_13_ ( .D(DP_pipe0_coeff_pipe00[13]), .CK(clk), 
        .RN(n1123), .Q(DP_pipe10[13]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_14_ ( .D(DP_pipe0_coeff_pipe00[14]), .CK(clk), 
        .RN(n1123), .Q(DP_pipe10[14]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_15_ ( .D(DP_pipe0_coeff_pipe00[15]), .CK(clk), 
        .RN(n1123), .Q(DP_pipe10[15]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_16_ ( .D(DP_pipe0_coeff_pipe00[16]), .CK(clk), 
        .RN(n1123), .Q(DP_pipe10[16]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_17_ ( .D(DP_pipe0_coeff_pipe00[17]), .CK(clk), 
        .RN(n1123), .Q(DP_pipe10[17]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_18_ ( .D(DP_pipe0_coeff_pipe00[18]), .CK(clk), 
        .RN(n1123), .Q(DP_pipe10[18]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_19_ ( .D(DP_pipe0_coeff_pipe00[19]), .CK(clk), 
        .RN(n1123), .Q(DP_pipe10[19]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_20_ ( .D(DP_pipe0_coeff_pipe00[20]), .CK(clk), 
        .RN(n1123), .Q(DP_pipe10[20]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_21_ ( .D(DP_pipe0_coeff_pipe00[21]), .CK(clk), 
        .RN(n1123), .Q(DP_pipe10[21]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_22_ ( .D(DP_pipe0_coeff_pipe00[22]), .CK(clk), 
        .RN(n1123), .Q(DP_pipe10[22]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_23_ ( .D(DP_pipe0_coeff_pipe00[23]), .CK(clk), 
        .RN(n1124), .Q(DP_pipe10[23]) );
  DFFR_X1 DP_reg_sw2_Q_reg_23_ ( .D(n606), .CK(clk), .RN(n1124), .Q(DP_sw2[23]), .QN(n339) );
  DFFR_X1 DP_reg_pipe03_Q_reg_23_ ( .D(DP_sw2[23]), .CK(clk), .RN(n1124), .Q(
        DP_pipe03[23]) );
  DFFR_X1 DP_reg_sw2_Q_reg_22_ ( .D(n604), .CK(clk), .RN(n1124), .Q(DP_sw2[22]), .QN(n338) );
  DFFR_X1 DP_reg_pipe03_Q_reg_22_ ( .D(DP_sw2[22]), .CK(clk), .RN(n1124), .Q(
        DP_pipe03[22]) );
  DFFR_X1 DP_reg_sw2_Q_reg_21_ ( .D(n602), .CK(clk), .RN(n1124), .Q(DP_sw2[21]), .QN(n337) );
  DFFR_X1 DP_reg_pipe03_Q_reg_21_ ( .D(DP_sw2[21]), .CK(clk), .RN(n1124), .Q(
        DP_pipe03[21]) );
  DFFR_X1 DP_reg_sw2_Q_reg_20_ ( .D(n600), .CK(clk), .RN(n1124), .Q(DP_sw2[20]), .QN(n336) );
  DFFR_X1 DP_reg_pipe03_Q_reg_20_ ( .D(DP_sw2[20]), .CK(clk), .RN(n1124), .Q(
        DP_pipe03[20]) );
  DFFR_X1 DP_reg_sw2_Q_reg_19_ ( .D(n598), .CK(clk), .RN(n1124), .Q(DP_sw2[19]), .QN(n335) );
  DFFR_X1 DP_reg_pipe03_Q_reg_19_ ( .D(DP_sw2[19]), .CK(clk), .RN(n1124), .Q(
        DP_pipe03[19]) );
  DFFR_X1 DP_reg_sw2_Q_reg_18_ ( .D(n596), .CK(clk), .RN(n1124), .Q(DP_sw2[18]), .QN(n334) );
  DFFR_X1 DP_reg_pipe03_Q_reg_18_ ( .D(DP_sw2[18]), .CK(clk), .RN(n1125), .Q(
        DP_pipe03[18]) );
  DFFR_X1 DP_reg_sw2_Q_reg_17_ ( .D(n594), .CK(clk), .RN(n1125), .Q(DP_sw2[17]), .QN(n333) );
  DFFR_X1 DP_reg_pipe03_Q_reg_17_ ( .D(DP_sw2[17]), .CK(clk), .RN(n1125), .Q(
        DP_pipe03[17]) );
  DFFR_X1 DP_reg_sw2_Q_reg_16_ ( .D(n592), .CK(clk), .RN(n1125), .Q(DP_sw2[16]), .QN(n332) );
  DFFR_X1 DP_reg_pipe03_Q_reg_16_ ( .D(DP_sw2[16]), .CK(clk), .RN(n1125), .Q(
        DP_pipe03[16]) );
  DFFR_X1 DP_reg_sw2_Q_reg_15_ ( .D(n590), .CK(clk), .RN(n1125), .Q(DP_sw2[15]), .QN(n331) );
  DFFR_X1 DP_reg_pipe03_Q_reg_15_ ( .D(DP_sw2[15]), .CK(clk), .RN(n1125), .Q(
        DP_pipe03[15]) );
  DFFR_X1 DP_reg_sw2_Q_reg_14_ ( .D(n588), .CK(clk), .RN(n1125), .Q(DP_sw2[14]), .QN(n330) );
  DFFR_X1 DP_reg_pipe03_Q_reg_14_ ( .D(DP_sw2[14]), .CK(clk), .RN(n1125), .Q(
        DP_pipe03[14]) );
  DFFR_X1 DP_reg_sw2_Q_reg_13_ ( .D(n586), .CK(clk), .RN(n1125), .Q(DP_sw2[13]), .QN(n329) );
  DFFR_X1 DP_reg_pipe03_Q_reg_13_ ( .D(DP_sw2[13]), .CK(clk), .RN(n1125), .Q(
        DP_pipe03[13]) );
  DFFR_X1 DP_reg_sw2_Q_reg_12_ ( .D(n584), .CK(clk), .RN(n1125), .Q(DP_sw2[12]), .QN(n328) );
  DFFR_X1 DP_reg_pipe03_Q_reg_12_ ( .D(DP_sw2[12]), .CK(clk), .RN(n1126), .Q(
        DP_pipe03[12]) );
  DFFR_X1 DP_reg_sw2_Q_reg_11_ ( .D(n582), .CK(clk), .RN(n1126), .Q(DP_sw2[11]), .QN(n327) );
  DFFR_X1 DP_reg_pipe03_Q_reg_11_ ( .D(DP_sw2[11]), .CK(clk), .RN(n1126), .Q(
        DP_pipe03[11]) );
  DFFR_X1 DP_reg_sw2_Q_reg_10_ ( .D(n580), .CK(clk), .RN(n1126), .Q(DP_sw2[10]), .QN(n326) );
  DFFR_X1 DP_reg_pipe03_Q_reg_10_ ( .D(DP_sw2[10]), .CK(clk), .RN(n1126), .Q(
        DP_pipe03[10]) );
  DFFR_X1 DP_reg_sw2_Q_reg_9_ ( .D(n578), .CK(clk), .RN(n1126), .Q(DP_sw2[9]), 
        .QN(n325) );
  DFFR_X1 DP_reg_pipe03_Q_reg_9_ ( .D(DP_sw2[9]), .CK(clk), .RN(n1126), .Q(
        DP_pipe03[9]) );
  DFFR_X1 DP_reg_sw2_Q_reg_8_ ( .D(n576), .CK(clk), .RN(n1126), .Q(DP_sw2[8]), 
        .QN(n324) );
  DFFR_X1 DP_reg_pipe03_Q_reg_8_ ( .D(DP_sw2[8]), .CK(clk), .RN(n1126), .Q(
        DP_pipe03[8]) );
  DFFR_X1 DP_reg_sw2_Q_reg_7_ ( .D(n574), .CK(clk), .RN(n1126), .Q(DP_sw2[7]), 
        .QN(n323) );
  DFFR_X1 DP_reg_pipe03_Q_reg_7_ ( .D(DP_sw2[7]), .CK(clk), .RN(n1126), .Q(
        DP_pipe03[7]) );
  DFFR_X1 DP_reg_sw2_Q_reg_6_ ( .D(n572), .CK(clk), .RN(n1126), .Q(DP_sw2[6]), 
        .QN(n322) );
  DFFR_X1 DP_reg_pipe03_Q_reg_6_ ( .D(DP_sw2[6]), .CK(clk), .RN(n1127), .Q(
        DP_pipe03[6]) );
  DFFR_X1 DP_reg_sw2_Q_reg_5_ ( .D(n570), .CK(clk), .RN(n1127), .Q(DP_sw2[5]), 
        .QN(n321) );
  DFFR_X1 DP_reg_pipe03_Q_reg_5_ ( .D(DP_sw2[5]), .CK(clk), .RN(n1127), .Q(
        DP_pipe03[5]) );
  DFFR_X1 DP_reg_sw2_Q_reg_4_ ( .D(n568), .CK(clk), .RN(n1127), .Q(DP_sw2[4]), 
        .QN(n320) );
  DFFR_X1 DP_reg_pipe03_Q_reg_4_ ( .D(DP_sw2[4]), .CK(clk), .RN(n1127), .Q(
        DP_pipe03[4]) );
  DFFR_X1 DP_reg_sw2_Q_reg_3_ ( .D(n566), .CK(clk), .RN(n1127), .Q(DP_sw2[3]), 
        .QN(n319) );
  DFFR_X1 DP_reg_pipe03_Q_reg_3_ ( .D(DP_sw2[3]), .CK(clk), .RN(n1127), .Q(
        DP_pipe03[3]) );
  DFFR_X1 DP_reg_sw2_Q_reg_2_ ( .D(n564), .CK(clk), .RN(n1127), .Q(DP_sw2[2]), 
        .QN(n318) );
  DFFR_X1 DP_reg_pipe03_Q_reg_2_ ( .D(DP_sw2[2]), .CK(clk), .RN(n1127), .Q(
        DP_pipe03[2]) );
  DFFR_X1 DP_reg_sw2_Q_reg_1_ ( .D(n562), .CK(clk), .RN(n1127), .Q(DP_sw2[1]), 
        .QN(n317) );
  DFFR_X1 DP_reg_pipe03_Q_reg_1_ ( .D(DP_sw2[1]), .CK(clk), .RN(n1127), .Q(
        DP_pipe03[1]) );
  DFFR_X1 DP_reg_sw2_Q_reg_0_ ( .D(n560), .CK(clk), .RN(n1127), .Q(DP_sw2[0]), 
        .QN(n316) );
  DFFR_X1 DP_reg_pipe03_Q_reg_0_ ( .D(DP_sw2[0]), .CK(clk), .RN(n1128), .Q(
        DP_pipe03[0]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_0_ ( .D(DP_pipe0_coeff_pipe03[0]), .CK(clk), 
        .RN(n1128), .Q(DP_pipe13[0]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_1_ ( .D(DP_pipe0_coeff_pipe03[1]), .CK(clk), 
        .RN(n1128), .Q(DP_pipe13[1]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_2_ ( .D(DP_pipe0_coeff_pipe03[2]), .CK(clk), 
        .RN(n1128), .Q(DP_pipe13[2]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_3_ ( .D(DP_pipe0_coeff_pipe03[3]), .CK(clk), 
        .RN(n1128), .Q(DP_pipe13[3]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_4_ ( .D(DP_pipe0_coeff_pipe03[4]), .CK(clk), 
        .RN(n1128), .Q(DP_pipe13[4]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_5_ ( .D(DP_pipe0_coeff_pipe03[5]), .CK(clk), 
        .RN(n1128), .Q(DP_pipe13[5]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_6_ ( .D(DP_pipe0_coeff_pipe03[6]), .CK(clk), 
        .RN(n1128), .Q(DP_pipe13[6]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_7_ ( .D(DP_pipe0_coeff_pipe03[7]), .CK(clk), 
        .RN(n1128), .Q(DP_pipe13[7]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_8_ ( .D(DP_pipe0_coeff_pipe03[8]), .CK(clk), 
        .RN(n1128), .Q(DP_pipe13[8]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_9_ ( .D(DP_pipe0_coeff_pipe03[9]), .CK(clk), 
        .RN(n1128), .Q(DP_pipe13[9]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_10_ ( .D(DP_pipe0_coeff_pipe03[10]), .CK(clk), 
        .RN(n1128), .Q(DP_pipe13[10]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_11_ ( .D(DP_pipe0_coeff_pipe03[11]), .CK(clk), 
        .RN(n1129), .Q(DP_pipe13[11]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_12_ ( .D(DP_pipe0_coeff_pipe03[12]), .CK(clk), 
        .RN(n1129), .Q(DP_pipe13[12]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_13_ ( .D(DP_pipe0_coeff_pipe03[13]), .CK(clk), 
        .RN(n1129), .Q(DP_pipe13[13]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_14_ ( .D(DP_pipe0_coeff_pipe03[14]), .CK(clk), 
        .RN(n1129), .Q(DP_pipe13[14]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_15_ ( .D(DP_pipe0_coeff_pipe03[15]), .CK(clk), 
        .RN(n1129), .Q(DP_pipe13[15]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_16_ ( .D(DP_pipe0_coeff_pipe03[16]), .CK(clk), 
        .RN(n1129), .Q(DP_pipe13[16]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_17_ ( .D(DP_pipe0_coeff_pipe03[17]), .CK(clk), 
        .RN(n1129), .Q(DP_pipe13[17]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_18_ ( .D(DP_pipe0_coeff_pipe03[18]), .CK(clk), 
        .RN(n1129), .Q(DP_pipe13[18]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_19_ ( .D(DP_pipe0_coeff_pipe03[19]), .CK(clk), 
        .RN(n1129), .Q(DP_pipe13[19]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_20_ ( .D(DP_pipe0_coeff_pipe03[20]), .CK(clk), 
        .RN(n1129), .Q(DP_pipe13[20]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_21_ ( .D(DP_pipe0_coeff_pipe03[21]), .CK(clk), 
        .RN(n1129), .Q(DP_pipe13[21]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_22_ ( .D(DP_pipe0_coeff_pipe03[22]), .CK(clk), 
        .RN(n1129), .Q(DP_pipe13[22]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_23_ ( .D(DP_pipe0_coeff_pipe03[23]), .CK(clk), 
        .RN(n1130), .Q(DP_pipe13[23]) );
  DFFR_X1 CU_presentState_reg_0_ ( .D(CU_nextState_0_), .CK(clk), .RN(n1130), 
        .QN(n315) );
  DFFR_X1 reg_delay_0_Q_reg_0_ ( .D(delayed_controls_0__1_), .CK(clk), .RN(
        n1130), .Q(delayed_controls_1__1_) );
  DFFR_X1 reg_delay_0_Q_reg_1_ ( .D(n1034), .CK(clk), .RN(n1130), .Q(
        delayed_controls_1__0_) );
  DFFR_X1 reg_delay_1_Q_reg_0_ ( .D(delayed_controls_1__1_), .CK(clk), .RN(
        n1130), .Q(vOut) );
  DFFR_X1 reg_delay_1_Q_reg_1_ ( .D(delayed_controls_1__0_), .CK(clk), .RN(
        n1130), .Q(delayed_controls_2__0_), .QN(n1028) );
  DFFR_X1 DP_reg_out_Q_reg_11_ ( .D(n531), .CK(clk), .RN(n1130), .Q(dOut[11]), 
        .QN(n313) );
  DFFR_X1 DP_reg_out_Q_reg_10_ ( .D(n530), .CK(clk), .RN(n1130), .Q(dOut[10]), 
        .QN(n312) );
  DFFR_X1 DP_reg_out_Q_reg_9_ ( .D(n529), .CK(clk), .RN(n1130), .Q(dOut[9]), 
        .QN(n311) );
  DFFR_X1 DP_reg_out_Q_reg_8_ ( .D(n528), .CK(clk), .RN(n1130), .Q(dOut[8]), 
        .QN(n310) );
  DFFR_X1 DP_reg_out_Q_reg_7_ ( .D(n527), .CK(clk), .RN(n1130), .Q(dOut[7]), 
        .QN(n309) );
  DFFR_X1 DP_reg_out_Q_reg_6_ ( .D(n526), .CK(clk), .RN(n1130), .Q(dOut[6]), 
        .QN(n308) );
  DFFR_X1 DP_reg_out_Q_reg_5_ ( .D(n525), .CK(clk), .RN(n1131), .Q(dOut[5]), 
        .QN(n307) );
  DFFR_X1 DP_reg_out_Q_reg_4_ ( .D(n524), .CK(clk), .RN(n1131), .Q(dOut[4]), 
        .QN(n306) );
  DFFR_X1 DP_reg_out_Q_reg_3_ ( .D(n523), .CK(clk), .RN(n1131), .Q(dOut[3]), 
        .QN(n305) );
  DFFR_X1 DP_reg_out_Q_reg_2_ ( .D(n522), .CK(clk), .RN(n1131), .Q(dOut[2]), 
        .QN(n304) );
  DFFR_X1 DP_reg_out_Q_reg_1_ ( .D(n521), .CK(clk), .RN(n1131), .Q(dOut[1]), 
        .QN(n303) );
  DFFR_X1 DP_reg_out_Q_reg_0_ ( .D(n520), .CK(clk), .RN(n1131), .Q(dOut[0]), 
        .QN(n302) );
  XOR2_X1 U501 ( .A(n1085), .B(n1034), .Z(CU_nextState_0_) );
  XOR2_X1 U503 ( .A(n315), .B(delayed_controls_0__1_), .Z(n74) );
  iir_filter_DW01_add_0 DP_add_223 ( .A({DP_pipe10[23], DP_pipe10[22], 
        DP_pipe10[21], DP_pipe10[20], DP_pipe10[19], DP_pipe10[18], 
        DP_pipe10[17], DP_pipe10[16], DP_pipe10[15], DP_pipe10[14], 
        DP_pipe10[13], DP_pipe10[12], DP_pipe10[11], DP_pipe10[10], 
        DP_pipe10[9], DP_pipe10[8], DP_pipe10[7], DP_pipe10[6], DP_pipe10[5], 
        DP_pipe10[4], DP_pipe10[3], DP_pipe10[2], DP_pipe10[1], DP_pipe10[0]}), 
        .B({DP_ff[23], DP_ff[22], DP_ff[21], DP_ff[20], DP_ff[19], DP_ff[18], 
        DP_ff[17], DP_ff[16], DP_ff[15], DP_ff[14], DP_ff[13], DP_ff[12], 
        DP_ff[11], DP_ff[10], DP_ff[9], DP_ff[8], DP_ff[7], DP_ff[6], DP_ff[5], 
        DP_ff[4], DP_ff[3], DP_ff[2], DP_ff[1], DP_ff[0]}), .CI(1'b0), .SUM({
        DP_y_23, DP_y_11_, DP_y_10_, DP_y_9_, DP_y_8_, DP_y_7_, DP_y_6_, 
        DP_y_5_, DP_y_4_, DP_y_3_, DP_y_2_, DP_y_1_, DP_y_0_, 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10}) );
  iir_filter_DW01_sub_0 DP_sub_217 ( .A({DP_x[11], DP_x[11], DP_x[10], DP_x[9], 
        DP_x[8], DP_x[7], DP_x[6], DP_x[5], DP_x[4], DP_x[3], DP_x[2], DP_x[1], 
        DP_x[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({DP_fb[23], DP_fb[22], DP_fb[21], DP_fb[20], DP_fb[19], 
        DP_fb[18], DP_fb[17], DP_fb[16], DP_fb[15], DP_fb[14], DP_fb[13], 
        DP_fb[12], DP_fb[11], DP_fb[10], DP_fb[9], DP_fb[8], DP_fb[7], 
        DP_fb[6], DP_fb[5], DP_fb[4], DP_fb[3], DP_fb[2], DP_fb[1], DP_fb[0]}), 
        .CI(1'b0), .DIFF({DP_w_23_, DP_w_22_, DP_w_21_, DP_w_20_, DP_w_19_, 
        DP_w_18_, DP_w_17_, DP_w_16_, DP_w_15_, DP_w_14_, DP_w_13_, DP_w_12_, 
        DP_w_11_, DP_w_10_, DP_w_9_, DP_w_8_, DP_w_7_, DP_w_6_, DP_w_5_, 
        DP_w_4_, DP_w_3_, DP_w_2_, DP_w_1_, DP_w_0_}) );
  iir_filter_DW01_add_1 DP_add_216 ( .A({DP_pipe11[23], DP_pipe11[22], 
        DP_pipe11[21], DP_pipe11[20], DP_pipe11[19], DP_pipe11[18], 
        DP_pipe11[17], DP_pipe11[16], DP_pipe11[15], DP_pipe11[14], 
        DP_pipe11[13], DP_pipe11[12], DP_pipe11[11], DP_pipe11[10], 
        DP_pipe11[9], DP_pipe11[8], DP_pipe11[7], DP_pipe11[6], DP_pipe11[5], 
        DP_pipe11[4], DP_pipe11[3], DP_pipe11[2], DP_pipe11[1], DP_pipe11[0]}), 
        .B({DP_ff_part[23], DP_ff_part[22], DP_ff_part[21], DP_ff_part[20], 
        DP_ff_part[19], DP_ff_part[18], DP_ff_part[17], DP_ff_part[16], 
        DP_ff_part[15], DP_ff_part[14], DP_ff_part[13], DP_ff_part[12], 
        DP_ff_part[11], DP_ff_part[10], DP_ff_part[9], DP_ff_part[8], 
        DP_ff_part[7], DP_ff_part[6], DP_ff_part[5], DP_ff_part[4], 
        DP_ff_part[3], DP_ff_part[2], DP_ff_part[1], DP_ff_part[0]}), .CI(1'b0), .SUM({DP_ff[23], DP_ff[22], DP_ff[21], DP_ff[20], DP_ff[19], DP_ff[18], 
        DP_ff[17], DP_ff[16], DP_ff[15], DP_ff[14], DP_ff[13], DP_ff[12], 
        DP_ff[11], DP_ff[10], DP_ff[9], DP_ff[8], DP_ff[7], DP_ff[6], DP_ff[5], 
        DP_ff[4], DP_ff[3], DP_ff[2], DP_ff[1], DP_ff[0]}) );
  iir_filter_DW01_add_2 DP_add_215 ( .A({DP_pipe12[23], DP_pipe12[22], 
        DP_pipe12[21], DP_pipe12[20], DP_pipe12[19], DP_pipe12[18], 
        DP_pipe12[17], DP_pipe12[16], DP_pipe12[15], DP_pipe12[14], 
        DP_pipe12[13], DP_pipe12[12], DP_pipe12[11], DP_pipe12[10], 
        DP_pipe12[9], DP_pipe12[8], DP_pipe12[7], DP_pipe12[6], DP_pipe12[5], 
        DP_pipe12[4], DP_pipe12[3], DP_pipe12[2], DP_pipe12[1], DP_pipe12[0]}), 
        .B({DP_pipe13[23], DP_pipe13[22], DP_pipe13[21], DP_pipe13[20], 
        DP_pipe13[19], DP_pipe13[18], DP_pipe13[17], DP_pipe13[16], 
        DP_pipe13[15], DP_pipe13[14], DP_pipe13[13], DP_pipe13[12], 
        DP_pipe13[11], DP_pipe13[10], DP_pipe13[9], DP_pipe13[8], DP_pipe13[7], 
        DP_pipe13[6], DP_pipe13[5], DP_pipe13[4], DP_pipe13[3], DP_pipe13[2], 
        DP_pipe13[1], DP_pipe13[0]}), .CI(1'b0), .SUM({DP_ff_part[23], 
        DP_ff_part[22], DP_ff_part[21], DP_ff_part[20], DP_ff_part[19], 
        DP_ff_part[18], DP_ff_part[17], DP_ff_part[16], DP_ff_part[15], 
        DP_ff_part[14], DP_ff_part[13], DP_ff_part[12], DP_ff_part[11], 
        DP_ff_part[10], DP_ff_part[9], DP_ff_part[8], DP_ff_part[7], 
        DP_ff_part[6], DP_ff_part[5], DP_ff_part[4], DP_ff_part[3], 
        DP_ff_part[2], DP_ff_part[1], DP_ff_part[0]}) );
  iir_filter_DW01_add_3 DP_add_214 ( .A({DP_ret0[23], DP_ret0[22], DP_ret0[21], 
        DP_ret0[20], DP_ret0[19], DP_ret0[18], DP_ret0[17], DP_ret0[16], 
        DP_ret0[15], DP_ret0[14], DP_ret0[13], DP_ret0[12], DP_ret0[11], 
        DP_ret0[10], DP_ret0[9], DP_ret0[8], DP_ret0[7], DP_ret0[6], 
        DP_ret0[5], DP_ret0[4], DP_ret0[3], DP_ret0[2], DP_ret0[1], DP_ret0[0]}), .B({DP_ret1[23], DP_ret1[22], DP_ret1[21], DP_ret1[20], DP_ret1[19], 
        DP_ret1[18], DP_ret1[17], DP_ret1[16], DP_ret1[15], DP_ret1[14], 
        DP_ret1[13], DP_ret1[12], DP_ret1[11], DP_ret1[10], DP_ret1[9], 
        DP_ret1[8], DP_ret1[7], DP_ret1[6], DP_ret1[5], DP_ret1[4], DP_ret1[3], 
        DP_ret1[2], DP_ret1[1], DP_ret1[0]}), .CI(1'b0), .SUM({DP_fb[23], 
        DP_fb[22], DP_fb[21], DP_fb[20], DP_fb[19], DP_fb[18], DP_fb[17], 
        DP_fb[16], DP_fb[15], DP_fb[14], DP_fb[13], DP_fb[12], DP_fb[11], 
        DP_fb[10], DP_fb[9], DP_fb[8], DP_fb[7], DP_fb[6], DP_fb[5], DP_fb[4], 
        DP_fb[3], DP_fb[2], DP_fb[1], DP_fb[0]}) );
  iir_filter_DW02_mult_0 DP_mult_209 ( .A({DP_coeffs_ff_int[72], 
        DP_coeffs_ff_int[73], DP_coeffs_ff_int[74], DP_coeffs_ff_int[75], 
        DP_coeffs_ff_int[76], DP_coeffs_ff_int[77], DP_coeffs_ff_int[78], 
        DP_coeffs_ff_int[79], DP_coeffs_ff_int[80], DP_coeffs_ff_int[81], 
        DP_coeffs_ff_int[82], DP_coeffs_ff_int[83], DP_coeffs_ff_int[84], 
        DP_coeffs_ff_int[85], DP_coeffs_ff_int[86], DP_coeffs_ff_int[87], 
        DP_coeffs_ff_int[88], DP_coeffs_ff_int[89], DP_coeffs_ff_int[90], 
        DP_coeffs_ff_int[91], DP_coeffs_ff_int[92], DP_coeffs_ff_int[93], 
        DP_coeffs_ff_int[94], DP_coeffs_ff_int[95]}), .B({DP_pipe03[23], 
        DP_pipe03[22], DP_pipe03[21], DP_pipe03[20], DP_pipe03[19], 
        DP_pipe03[18], DP_pipe03[17], DP_pipe03[16], DP_pipe03[15], 
        DP_pipe03[14], DP_pipe03[13], DP_pipe03[12], DP_pipe03[11], 
        DP_pipe03[10], DP_pipe03[9], DP_pipe03[8], DP_pipe03[7], DP_pipe03[6], 
        DP_pipe03[5], DP_pipe03[4], DP_pipe03[3], DP_pipe03[2], DP_pipe03[1], 
        DP_pipe03[0]}), .TC(1'b1), .PRODUCT({DP_pipe0_coeff_pipe03[23], 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        DP_pipe0_coeff_pipe03[22], DP_pipe0_coeff_pipe03[21], 
        DP_pipe0_coeff_pipe03[20], DP_pipe0_coeff_pipe03[19], 
        DP_pipe0_coeff_pipe03[18], DP_pipe0_coeff_pipe03[17], 
        DP_pipe0_coeff_pipe03[16], DP_pipe0_coeff_pipe03[15], 
        DP_pipe0_coeff_pipe03[14], DP_pipe0_coeff_pipe03[13], 
        DP_pipe0_coeff_pipe03[12], DP_pipe0_coeff_pipe03[11], 
        DP_pipe0_coeff_pipe03[10], DP_pipe0_coeff_pipe03[9], 
        DP_pipe0_coeff_pipe03[8], DP_pipe0_coeff_pipe03[7], 
        DP_pipe0_coeff_pipe03[6], DP_pipe0_coeff_pipe03[5], 
        DP_pipe0_coeff_pipe03[4], DP_pipe0_coeff_pipe03[3], 
        DP_pipe0_coeff_pipe03[2], DP_pipe0_coeff_pipe03[1], 
        DP_pipe0_coeff_pipe03[0], SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34}) );
  iir_filter_DW02_mult_1 DP_mult_208 ( .A({DP_coeffs_ff_int[48], 
        DP_coeffs_ff_int[49], DP_coeffs_ff_int[50], DP_coeffs_ff_int[51], 
        DP_coeffs_ff_int[52], DP_coeffs_ff_int[53], DP_coeffs_ff_int[54], 
        DP_coeffs_ff_int[55], DP_coeffs_ff_int[56], DP_coeffs_ff_int[57], 
        DP_coeffs_ff_int[58], DP_coeffs_ff_int[59], DP_coeffs_ff_int[60], 
        DP_coeffs_ff_int[61], DP_coeffs_ff_int[62], DP_coeffs_ff_int[63], 
        DP_coeffs_ff_int[64], DP_coeffs_ff_int[65], DP_coeffs_ff_int[66], 
        DP_coeffs_ff_int[67], DP_coeffs_ff_int[68], DP_coeffs_ff_int[69], 
        DP_coeffs_ff_int[70], DP_coeffs_ff_int[71]}), .B({DP_pipe02[23], 
        DP_pipe02[22], DP_pipe02[21], DP_pipe02[20], DP_pipe02[19], 
        DP_pipe02[18], DP_pipe02[17], DP_pipe02[16], DP_pipe02[15], 
        DP_pipe02[14], DP_pipe02[13], DP_pipe02[12], DP_pipe02[11], 
        DP_pipe02[10], DP_pipe02[9], DP_pipe02[8], DP_pipe02[7], DP_pipe02[6], 
        DP_pipe02[5], DP_pipe02[4], DP_pipe02[3], DP_pipe02[2], DP_pipe02[1], 
        DP_pipe02[0]}), .TC(1'b1), .PRODUCT({DP_pipe0_coeff_pipe02[23], 
        SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, 
        DP_pipe0_coeff_pipe02[22], DP_pipe0_coeff_pipe02[21], 
        DP_pipe0_coeff_pipe02[20], DP_pipe0_coeff_pipe02[19], 
        DP_pipe0_coeff_pipe02[18], DP_pipe0_coeff_pipe02[17], 
        DP_pipe0_coeff_pipe02[16], DP_pipe0_coeff_pipe02[15], 
        DP_pipe0_coeff_pipe02[14], DP_pipe0_coeff_pipe02[13], 
        DP_pipe0_coeff_pipe02[12], DP_pipe0_coeff_pipe02[11], 
        DP_pipe0_coeff_pipe02[10], DP_pipe0_coeff_pipe02[9], 
        DP_pipe0_coeff_pipe02[8], DP_pipe0_coeff_pipe02[7], 
        DP_pipe0_coeff_pipe02[6], DP_pipe0_coeff_pipe02[5], 
        DP_pipe0_coeff_pipe02[4], DP_pipe0_coeff_pipe02[3], 
        DP_pipe0_coeff_pipe02[2], DP_pipe0_coeff_pipe02[1], 
        DP_pipe0_coeff_pipe02[0], SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58}) );
  iir_filter_DW02_mult_2 DP_mult_207 ( .A({DP_coeffs_ff_int[24], 
        DP_coeffs_ff_int[25], DP_coeffs_ff_int[26], DP_coeffs_ff_int[27], 
        DP_coeffs_ff_int[28], DP_coeffs_ff_int[29], DP_coeffs_ff_int[30], 
        DP_coeffs_ff_int[31], DP_coeffs_ff_int[32], DP_coeffs_ff_int[33], 
        DP_coeffs_ff_int[34], DP_coeffs_ff_int[35], DP_coeffs_ff_int[36], 
        DP_coeffs_ff_int[37], DP_coeffs_ff_int[38], DP_coeffs_ff_int[39], 
        DP_coeffs_ff_int[40], DP_coeffs_ff_int[41], DP_coeffs_ff_int[42], 
        DP_coeffs_ff_int[43], DP_coeffs_ff_int[44], DP_coeffs_ff_int[45], 
        DP_coeffs_ff_int[46], DP_coeffs_ff_int[47]}), .B({DP_pipe01[23], 
        DP_pipe01[22], DP_pipe01[21], DP_pipe01[20], DP_pipe01[19], 
        DP_pipe01[18], DP_pipe01[17], DP_pipe01[16], DP_pipe01[15], 
        DP_pipe01[14], DP_pipe01[13], DP_pipe01[12], DP_pipe01[11], 
        DP_pipe01[10], DP_pipe01[9], DP_pipe01[8], DP_pipe01[7], DP_pipe01[6], 
        DP_pipe01[5], DP_pipe01[4], DP_pipe01[3], DP_pipe01[2], DP_pipe01[1], 
        DP_pipe01[0]}), .TC(1'b1), .PRODUCT({DP_pipe0_coeff_pipe01[23], 
        SYNOPSYS_UNCONNECTED__59, SYNOPSYS_UNCONNECTED__60, 
        DP_pipe0_coeff_pipe01[22], DP_pipe0_coeff_pipe01[21], 
        DP_pipe0_coeff_pipe01[20], DP_pipe0_coeff_pipe01[19], 
        DP_pipe0_coeff_pipe01[18], DP_pipe0_coeff_pipe01[17], 
        DP_pipe0_coeff_pipe01[16], DP_pipe0_coeff_pipe01[15], 
        DP_pipe0_coeff_pipe01[14], DP_pipe0_coeff_pipe01[13], 
        DP_pipe0_coeff_pipe01[12], DP_pipe0_coeff_pipe01[11], 
        DP_pipe0_coeff_pipe01[10], DP_pipe0_coeff_pipe01[9], 
        DP_pipe0_coeff_pipe01[8], DP_pipe0_coeff_pipe01[7], 
        DP_pipe0_coeff_pipe01[6], DP_pipe0_coeff_pipe01[5], 
        DP_pipe0_coeff_pipe01[4], DP_pipe0_coeff_pipe01[3], 
        DP_pipe0_coeff_pipe01[2], DP_pipe0_coeff_pipe01[1], 
        DP_pipe0_coeff_pipe01[0], SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82}) );
  iir_filter_DW02_mult_3 DP_mult_206 ( .A({DP_coeffs_ff_int[0], 
        DP_coeffs_ff_int[1], DP_coeffs_ff_int[2], DP_coeffs_ff_int[3], 
        DP_coeffs_ff_int[4], DP_coeffs_ff_int[5], DP_coeffs_ff_int[6], 
        DP_coeffs_ff_int[7], DP_coeffs_ff_int[8], DP_coeffs_ff_int[9], 
        DP_coeffs_ff_int[10], DP_coeffs_ff_int[11], DP_coeffs_ff_int[12], 
        DP_coeffs_ff_int[13], DP_coeffs_ff_int[14], DP_coeffs_ff_int[15], 
        DP_coeffs_ff_int[16], DP_coeffs_ff_int[17], DP_coeffs_ff_int[18], 
        DP_coeffs_ff_int[19], DP_coeffs_ff_int[20], DP_coeffs_ff_int[21], 
        DP_coeffs_ff_int[22], DP_coeffs_ff_int[23]}), .B({DP_pipe00[23], 
        DP_pipe00[22], DP_pipe00[21], DP_pipe00[20], DP_pipe00[19], 
        DP_pipe00[18], DP_pipe00[17], DP_pipe00[16], DP_pipe00[15], 
        DP_pipe00[14], DP_pipe00[13], DP_pipe00[12], DP_pipe00[11], 
        DP_pipe00[10], DP_pipe00[9], DP_pipe00[8], DP_pipe00[7], DP_pipe00[6], 
        DP_pipe00[5], DP_pipe00[4], DP_pipe00[3], DP_pipe00[2], DP_pipe00[1], 
        DP_pipe00[0]}), .TC(1'b1), .PRODUCT({DP_pipe0_coeff_pipe00[23], 
        SYNOPSYS_UNCONNECTED__83, SYNOPSYS_UNCONNECTED__84, 
        DP_pipe0_coeff_pipe00[22], DP_pipe0_coeff_pipe00[21], 
        DP_pipe0_coeff_pipe00[20], DP_pipe0_coeff_pipe00[19], 
        DP_pipe0_coeff_pipe00[18], DP_pipe0_coeff_pipe00[17], 
        DP_pipe0_coeff_pipe00[16], DP_pipe0_coeff_pipe00[15], 
        DP_pipe0_coeff_pipe00[14], DP_pipe0_coeff_pipe00[13], 
        DP_pipe0_coeff_pipe00[12], DP_pipe0_coeff_pipe00[11], 
        DP_pipe0_coeff_pipe00[10], DP_pipe0_coeff_pipe00[9], 
        DP_pipe0_coeff_pipe00[8], DP_pipe0_coeff_pipe00[7], 
        DP_pipe0_coeff_pipe00[6], DP_pipe0_coeff_pipe00[5], 
        DP_pipe0_coeff_pipe00[4], DP_pipe0_coeff_pipe00[3], 
        DP_pipe0_coeff_pipe00[2], DP_pipe0_coeff_pipe00[1], 
        DP_pipe0_coeff_pipe00[0], SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106}) );
  iir_filter_DW02_mult_4 DP_mult_205 ( .A({DP_coeffs_fb_int[24], 
        DP_coeffs_fb_int[25], DP_coeffs_fb_int[26], DP_coeffs_fb_int[27], 
        DP_coeffs_fb_int[28], DP_coeffs_fb_int[29], DP_coeffs_fb_int[30], 
        DP_coeffs_fb_int[31], DP_coeffs_fb_int[32], DP_coeffs_fb_int[33], 
        DP_coeffs_fb_int[34], DP_coeffs_fb_int[35], DP_coeffs_fb_int[36], 
        DP_coeffs_fb_int[37], DP_coeffs_fb_int[38], DP_coeffs_fb_int[39], 
        DP_coeffs_fb_int[40], DP_coeffs_fb_int[41], DP_coeffs_fb_int[42], 
        DP_coeffs_fb_int[43], DP_coeffs_fb_int[44], DP_coeffs_fb_int[45], 
        DP_coeffs_fb_int[46], DP_coeffs_fb_int[47]}), .B({DP_sw1_23_, 
        DP_sw1_22_, DP_sw1_21_, DP_sw1_20_, DP_sw1_19_, DP_sw1_18_, DP_sw1_17_, 
        DP_sw1_16_, DP_sw1_15_, DP_sw1_14_, DP_sw1_13_, DP_sw1_12_, DP_sw1_11_, 
        DP_sw1_10_, DP_sw1_9_, DP_sw1_8_, DP_sw1_7_, DP_sw1_6_, DP_sw1_5_, 
        DP_sw1_4_, DP_sw1_3_, DP_sw1_2_, DP_sw1_1_, DP_sw1_0_}), .TC(1'b1), 
        .PRODUCT({DP_sw1_coeff_ret1[23], SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, DP_sw1_coeff_ret1[22], 
        DP_sw1_coeff_ret1[21], DP_sw1_coeff_ret1[20], DP_sw1_coeff_ret1[19], 
        DP_sw1_coeff_ret1[18], DP_sw1_coeff_ret1[17], DP_sw1_coeff_ret1[16], 
        DP_sw1_coeff_ret1[15], DP_sw1_coeff_ret1[14], DP_sw1_coeff_ret1[13], 
        DP_sw1_coeff_ret1[12], DP_sw1_coeff_ret1[11], DP_sw1_coeff_ret1[10], 
        DP_sw1_coeff_ret1[9], DP_sw1_coeff_ret1[8], DP_sw1_coeff_ret1[7], 
        DP_sw1_coeff_ret1[6], DP_sw1_coeff_ret1[5], DP_sw1_coeff_ret1[4], 
        DP_sw1_coeff_ret1[3], DP_sw1_coeff_ret1[2], DP_sw1_coeff_ret1[1], 
        DP_sw1_coeff_ret1[0], SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130}) );
  iir_filter_DW02_mult_5 DP_mult_204 ( .A({DP_coeffs_fb_int[0], 
        DP_coeffs_fb_int[1], DP_coeffs_fb_int[2], DP_coeffs_fb_int[3], 
        DP_coeffs_fb_int[4], DP_coeffs_fb_int[5], DP_coeffs_fb_int[6], 
        DP_coeffs_fb_int[7], DP_coeffs_fb_int[8], DP_coeffs_fb_int[9], 
        DP_coeffs_fb_int[10], DP_coeffs_fb_int[11], DP_coeffs_fb_int[12], 
        DP_coeffs_fb_int[13], DP_coeffs_fb_int[14], DP_coeffs_fb_int[15], 
        DP_coeffs_fb_int[16], DP_coeffs_fb_int[17], DP_coeffs_fb_int[18], 
        DP_coeffs_fb_int[19], DP_coeffs_fb_int[20], DP_coeffs_fb_int[21], 
        DP_coeffs_fb_int[22], DP_coeffs_fb_int[23]}), .B({DP_sw0_23_, 
        DP_sw0_22_, DP_sw0_21_, DP_sw0_20_, DP_sw0_19_, DP_sw0_18_, DP_sw0_17_, 
        DP_sw0_16_, DP_sw0_15_, DP_sw0_14_, DP_sw0_13_, DP_sw0_12_, DP_sw0_11_, 
        DP_sw0_10_, DP_sw0_9_, DP_sw0_8_, DP_sw0_7_, DP_sw0_6_, DP_sw0_5_, 
        DP_sw0_4_, DP_sw0_3_, DP_sw0_2_, DP_sw0_1_, DP_sw0_0_}), .TC(1'b1), 
        .PRODUCT({DP_sw0_coeff_ret0[23], SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, DP_sw0_coeff_ret0[22], 
        DP_sw0_coeff_ret0[21], DP_sw0_coeff_ret0[20], DP_sw0_coeff_ret0[19], 
        DP_sw0_coeff_ret0[18], DP_sw0_coeff_ret0[17], DP_sw0_coeff_ret0[16], 
        DP_sw0_coeff_ret0[15], DP_sw0_coeff_ret0[14], DP_sw0_coeff_ret0[13], 
        DP_sw0_coeff_ret0[12], DP_sw0_coeff_ret0[11], DP_sw0_coeff_ret0[10], 
        DP_sw0_coeff_ret0[9], DP_sw0_coeff_ret0[8], DP_sw0_coeff_ret0[7], 
        DP_sw0_coeff_ret0[6], DP_sw0_coeff_ret0[5], DP_sw0_coeff_ret0[4], 
        DP_sw0_coeff_ret0[3], DP_sw0_coeff_ret0[2], DP_sw0_coeff_ret0[1], 
        DP_sw0_coeff_ret0[0], SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154}) );
  INV_X1 U504 ( .A(n1049), .ZN(n1033) );
  BUF_X1 U505 ( .A(n1051), .Z(n1049) );
  BUF_X1 U506 ( .A(n1058), .Z(n1036) );
  BUF_X1 U507 ( .A(n1057), .Z(n1037) );
  BUF_X1 U508 ( .A(n1058), .Z(n1035) );
  BUF_X1 U509 ( .A(n1057), .Z(n1038) );
  BUF_X1 U510 ( .A(n1056), .Z(n1039) );
  BUF_X1 U511 ( .A(n1052), .Z(n1048) );
  BUF_X1 U512 ( .A(n1052), .Z(n1047) );
  BUF_X1 U513 ( .A(n1053), .Z(n1046) );
  BUF_X1 U514 ( .A(n1054), .Z(n1044) );
  BUF_X1 U515 ( .A(n1053), .Z(n1045) );
  BUF_X1 U516 ( .A(n1054), .Z(n1043) );
  BUF_X1 U517 ( .A(n1055), .Z(n1042) );
  BUF_X1 U518 ( .A(n1056), .Z(n1040) );
  BUF_X1 U519 ( .A(n1055), .Z(n1041) );
  BUF_X1 U520 ( .A(n1051), .Z(n1050) );
  BUF_X1 U521 ( .A(n1087), .Z(n1061) );
  BUF_X1 U522 ( .A(n1087), .Z(n1062) );
  BUF_X1 U523 ( .A(n1087), .Z(n1063) );
  BUF_X1 U524 ( .A(n1087), .Z(n1064) );
  BUF_X1 U525 ( .A(n1086), .Z(n1067) );
  BUF_X1 U526 ( .A(n1086), .Z(n1068) );
  BUF_X1 U527 ( .A(n1086), .Z(n1070) );
  BUF_X1 U528 ( .A(n1086), .Z(n1069) );
  BUF_X1 U529 ( .A(n1087), .Z(n1066) );
  BUF_X1 U530 ( .A(n1087), .Z(n1065) );
  BUF_X1 U531 ( .A(n1088), .Z(n1059) );
  BUF_X1 U532 ( .A(n1088), .Z(n1060) );
  BUF_X1 U533 ( .A(n1085), .Z(n1078) );
  BUF_X1 U534 ( .A(n1085), .Z(n1077) );
  BUF_X1 U535 ( .A(n1085), .Z(n1076) );
  BUF_X1 U536 ( .A(n1085), .Z(n1073) );
  BUF_X1 U537 ( .A(n1086), .Z(n1072) );
  BUF_X1 U538 ( .A(n1085), .Z(n1074) );
  BUF_X1 U539 ( .A(n1085), .Z(n1075) );
  BUF_X1 U540 ( .A(n1084), .Z(n1082) );
  BUF_X1 U541 ( .A(n1084), .Z(n1081) );
  BUF_X1 U542 ( .A(n1084), .Z(n1080) );
  BUF_X1 U543 ( .A(n1084), .Z(n1079) );
  BUF_X1 U544 ( .A(n1084), .Z(n1083) );
  BUF_X1 U545 ( .A(n1086), .Z(n1071) );
  BUF_X1 U546 ( .A(n1029), .Z(n1051) );
  BUF_X1 U547 ( .A(n1029), .Z(n1052) );
  BUF_X1 U548 ( .A(n1029), .Z(n1053) );
  BUF_X1 U549 ( .A(n1030), .Z(n1054) );
  BUF_X1 U550 ( .A(n1030), .Z(n1056) );
  BUF_X1 U551 ( .A(n1030), .Z(n1055) );
  BUF_X1 U552 ( .A(n1031), .Z(n1058) );
  BUF_X1 U553 ( .A(n1031), .Z(n1057) );
  BUF_X1 U554 ( .A(n1089), .Z(n1086) );
  BUF_X1 U555 ( .A(n1089), .Z(n1087) );
  BUF_X1 U556 ( .A(n1090), .Z(n1085) );
  BUF_X1 U557 ( .A(n1090), .Z(n1084) );
  BUF_X1 U558 ( .A(n1089), .Z(n1088) );
  BUF_X1 U559 ( .A(n74), .Z(n1029) );
  BUF_X1 U560 ( .A(n74), .Z(n1030) );
  BUF_X1 U561 ( .A(n74), .Z(n1031) );
  OR2_X1 U562 ( .A1(n1028), .A2(DP_N4), .ZN(n58) );
  OAI221_X1 U563 ( .B1(n58), .B2(n59), .C1(delayed_controls_2__0_), .C2(n302), 
        .A(n60), .ZN(n520) );
  INV_X1 U564 ( .A(DP_y_0_), .ZN(n59) );
  OAI221_X1 U565 ( .B1(n58), .B2(n61), .C1(delayed_controls_2__0_), .C2(n303), 
        .A(n60), .ZN(n521) );
  INV_X1 U566 ( .A(DP_y_1_), .ZN(n61) );
  OAI221_X1 U567 ( .B1(n58), .B2(n62), .C1(delayed_controls_2__0_), .C2(n304), 
        .A(n60), .ZN(n522) );
  INV_X1 U568 ( .A(DP_y_2_), .ZN(n62) );
  OAI221_X1 U569 ( .B1(n58), .B2(n63), .C1(delayed_controls_2__0_), .C2(n305), 
        .A(n60), .ZN(n523) );
  INV_X1 U570 ( .A(DP_y_3_), .ZN(n63) );
  OAI221_X1 U571 ( .B1(n58), .B2(n64), .C1(delayed_controls_2__0_), .C2(n306), 
        .A(n60), .ZN(n524) );
  INV_X1 U572 ( .A(DP_y_4_), .ZN(n64) );
  OAI221_X1 U573 ( .B1(n58), .B2(n65), .C1(delayed_controls_2__0_), .C2(n307), 
        .A(n60), .ZN(n525) );
  INV_X1 U574 ( .A(DP_y_5_), .ZN(n65) );
  OAI221_X1 U575 ( .B1(n58), .B2(n66), .C1(delayed_controls_2__0_), .C2(n308), 
        .A(n60), .ZN(n526) );
  INV_X1 U576 ( .A(DP_y_6_), .ZN(n66) );
  OAI221_X1 U577 ( .B1(n58), .B2(n67), .C1(delayed_controls_2__0_), .C2(n309), 
        .A(n60), .ZN(n527) );
  INV_X1 U578 ( .A(DP_y_7_), .ZN(n67) );
  OAI221_X1 U579 ( .B1(n58), .B2(n68), .C1(delayed_controls_2__0_), .C2(n310), 
        .A(n60), .ZN(n528) );
  INV_X1 U580 ( .A(DP_y_8_), .ZN(n68) );
  OAI221_X1 U581 ( .B1(n58), .B2(n69), .C1(delayed_controls_2__0_), .C2(n311), 
        .A(n60), .ZN(n529) );
  INV_X1 U582 ( .A(DP_y_9_), .ZN(n69) );
  OAI221_X1 U583 ( .B1(n58), .B2(n70), .C1(delayed_controls_2__0_), .C2(n312), 
        .A(n60), .ZN(n530) );
  INV_X1 U584 ( .A(DP_y_10_), .ZN(n70) );
  NAND2_X1 U585 ( .A1(delayed_controls_2__0_), .A2(DP_N2), .ZN(n60) );
  OAI21_X1 U586 ( .B1(delayed_controls_2__0_), .B2(n313), .A(n72), .ZN(n531)
         );
  OAI211_X1 U587 ( .C1(DP_N4), .C2(DP_y_23), .A(n73), .B(
        delayed_controls_2__0_), .ZN(n72) );
  INV_X1 U588 ( .A(DP_N2), .ZN(n73) );
  INV_X1 U589 ( .A(n102), .ZN(n712) );
  AOI22_X1 U590 ( .A1(n1033), .A2(DP_w_22_), .B1(n1048), .B2(DP_sw0_22_), .ZN(
        n102) );
  INV_X1 U591 ( .A(n108), .ZN(n727) );
  AOI22_X1 U592 ( .A1(n1034), .A2(DP_w_19_), .B1(n1047), .B2(DP_sw0_19_), .ZN(
        n108) );
  INV_X1 U593 ( .A(n110), .ZN(n732) );
  AOI22_X1 U594 ( .A1(n1032), .A2(DP_w_18_), .B1(n1047), .B2(DP_sw0_18_), .ZN(
        n110) );
  INV_X1 U595 ( .A(n112), .ZN(n737) );
  AOI22_X1 U596 ( .A1(n1032), .A2(DP_w_17_), .B1(n1046), .B2(DP_sw0_17_), .ZN(
        n112) );
  INV_X1 U597 ( .A(n104), .ZN(n717) );
  AOI22_X1 U598 ( .A1(n1032), .A2(DP_w_21_), .B1(n1048), .B2(DP_sw0_21_), .ZN(
        n104) );
  INV_X1 U599 ( .A(n106), .ZN(n722) );
  AOI22_X1 U600 ( .A1(n1033), .A2(DP_w_20_), .B1(n1047), .B2(DP_sw0_20_), .ZN(
        n106) );
  INV_X1 U601 ( .A(n100), .ZN(n707) );
  AOI22_X1 U602 ( .A1(n1034), .A2(DP_w_23_), .B1(n1049), .B2(DP_sw0_23_), .ZN(
        n100) );
  INV_X1 U603 ( .A(n114), .ZN(n742) );
  AOI22_X1 U604 ( .A1(n1033), .A2(DP_w_16_), .B1(n1046), .B2(DP_sw0_16_), .ZN(
        n114) );
  INV_X1 U605 ( .A(n124), .ZN(n767) );
  AOI22_X1 U606 ( .A1(n1034), .A2(DP_w_11_), .B1(n1044), .B2(DP_sw0_11_), .ZN(
        n124) );
  INV_X1 U607 ( .A(n126), .ZN(n772) );
  AOI22_X1 U608 ( .A1(n1033), .A2(DP_w_10_), .B1(n1043), .B2(DP_sw0_10_), .ZN(
        n126) );
  INV_X1 U609 ( .A(n128), .ZN(n777) );
  AOI22_X1 U610 ( .A1(n1033), .A2(DP_w_9_), .B1(n1045), .B2(DP_sw0_9_), .ZN(
        n128) );
  INV_X1 U611 ( .A(n130), .ZN(n782) );
  AOI22_X1 U612 ( .A1(n1033), .A2(DP_w_8_), .B1(n1043), .B2(DP_sw0_8_), .ZN(
        n130) );
  INV_X1 U613 ( .A(n132), .ZN(n787) );
  AOI22_X1 U614 ( .A1(n1033), .A2(DP_w_7_), .B1(n1042), .B2(DP_sw0_7_), .ZN(
        n132) );
  INV_X1 U615 ( .A(n134), .ZN(n792) );
  AOI22_X1 U616 ( .A1(n1033), .A2(DP_w_6_), .B1(n1042), .B2(DP_sw0_6_), .ZN(
        n134) );
  INV_X1 U617 ( .A(n116), .ZN(n747) );
  AOI22_X1 U618 ( .A1(n1033), .A2(DP_w_15_), .B1(n1045), .B2(DP_sw0_15_), .ZN(
        n116) );
  INV_X1 U619 ( .A(n118), .ZN(n752) );
  AOI22_X1 U620 ( .A1(n1034), .A2(DP_w_14_), .B1(n1045), .B2(DP_sw0_14_), .ZN(
        n118) );
  INV_X1 U621 ( .A(n120), .ZN(n757) );
  AOI22_X1 U622 ( .A1(n1033), .A2(DP_w_13_), .B1(n1044), .B2(DP_sw0_13_), .ZN(
        n120) );
  INV_X1 U623 ( .A(n122), .ZN(n762) );
  AOI22_X1 U624 ( .A1(n1034), .A2(DP_w_12_), .B1(n1044), .B2(DP_sw0_12_), .ZN(
        n122) );
  OAI22_X1 U625 ( .A1(n1035), .A2(n1003), .B1(n1032), .B2(n316), .ZN(n560) );
  OAI22_X1 U626 ( .A1(n1035), .A2(n1006), .B1(n1032), .B2(n317), .ZN(n562) );
  OAI22_X1 U627 ( .A1(n1036), .A2(n1007), .B1(n1032), .B2(n318), .ZN(n564) );
  OAI22_X1 U628 ( .A1(n1035), .A2(n1008), .B1(n1032), .B2(n319), .ZN(n566) );
  OAI22_X1 U629 ( .A1(n1036), .A2(n1009), .B1(n1032), .B2(n320), .ZN(n568) );
  OAI22_X1 U630 ( .A1(n1036), .A2(n1010), .B1(n1032), .B2(n321), .ZN(n570) );
  OAI22_X1 U631 ( .A1(n1036), .A2(n1011), .B1(n1032), .B2(n322), .ZN(n572) );
  OAI22_X1 U632 ( .A1(n1036), .A2(n1012), .B1(n1032), .B2(n323), .ZN(n574) );
  OAI22_X1 U633 ( .A1(n1037), .A2(n1013), .B1(n1032), .B2(n324), .ZN(n576) );
  OAI22_X1 U634 ( .A1(n1037), .A2(n1014), .B1(n1032), .B2(n325), .ZN(n578) );
  OAI22_X1 U635 ( .A1(n1037), .A2(n1015), .B1(n1032), .B2(n326), .ZN(n580) );
  OAI22_X1 U636 ( .A1(n1037), .A2(n1016), .B1(n1032), .B2(n327), .ZN(n582) );
  OAI22_X1 U637 ( .A1(n1038), .A2(n1017), .B1(n1034), .B2(n328), .ZN(n584) );
  OAI22_X1 U638 ( .A1(n1035), .A2(n1018), .B1(n1033), .B2(n329), .ZN(n586) );
  OAI22_X1 U639 ( .A1(n1038), .A2(n1019), .B1(n1032), .B2(n330), .ZN(n588) );
  OAI22_X1 U640 ( .A1(n1037), .A2(n1020), .B1(n1034), .B2(n331), .ZN(n590) );
  OAI22_X1 U641 ( .A1(n1038), .A2(n1021), .B1(n1033), .B2(n332), .ZN(n592) );
  OAI22_X1 U642 ( .A1(n1039), .A2(n1022), .B1(n1033), .B2(n333), .ZN(n594) );
  OAI22_X1 U643 ( .A1(n1039), .A2(n1023), .B1(n1032), .B2(n334), .ZN(n596) );
  OAI22_X1 U644 ( .A1(n1038), .A2(n1024), .B1(n1032), .B2(n335), .ZN(n598) );
  OAI22_X1 U645 ( .A1(n1039), .A2(n1025), .B1(n1032), .B2(n336), .ZN(n600) );
  OAI22_X1 U646 ( .A1(n1035), .A2(n1026), .B1(n1032), .B2(n337), .ZN(n602) );
  OAI22_X1 U647 ( .A1(n1039), .A2(n1027), .B1(n1032), .B2(n338), .ZN(n604) );
  OAI22_X1 U648 ( .A1(n1038), .A2(n1004), .B1(n1032), .B2(n339), .ZN(n606) );
  OAI22_X1 U649 ( .A1(n1039), .A2(n1005), .B1(n1034), .B2(n1003), .ZN(n846) );
  INV_X1 U650 ( .A(n136), .ZN(n797) );
  AOI22_X1 U651 ( .A1(n1033), .A2(DP_w_5_), .B1(n1041), .B2(DP_sw0_5_), .ZN(
        n136) );
  INV_X1 U652 ( .A(n138), .ZN(n802) );
  AOI22_X1 U653 ( .A1(n1034), .A2(DP_w_4_), .B1(n1041), .B2(DP_sw0_4_), .ZN(
        n138) );
  OAI21_X1 U654 ( .B1(n1074), .B2(n389), .A(n147), .ZN(n847) );
  NAND2_X1 U655 ( .A1(coeffs_ff[23]), .A2(n1065), .ZN(n147) );
  OAI21_X1 U656 ( .B1(n1074), .B2(n390), .A(n148), .ZN(n848) );
  NAND2_X1 U657 ( .A1(coeffs_ff[22]), .A2(n1065), .ZN(n148) );
  OAI21_X1 U658 ( .B1(n1073), .B2(n391), .A(n149), .ZN(n849) );
  NAND2_X1 U659 ( .A1(coeffs_ff[21]), .A2(n1064), .ZN(n149) );
  OAI21_X1 U660 ( .B1(n1073), .B2(n392), .A(n150), .ZN(n850) );
  NAND2_X1 U661 ( .A1(coeffs_ff[20]), .A2(n1064), .ZN(n150) );
  OAI21_X1 U662 ( .B1(n1073), .B2(n393), .A(n151), .ZN(n851) );
  NAND2_X1 U663 ( .A1(coeffs_ff[19]), .A2(n1064), .ZN(n151) );
  OAI21_X1 U664 ( .B1(n1072), .B2(n394), .A(n152), .ZN(n852) );
  NAND2_X1 U665 ( .A1(coeffs_ff[18]), .A2(n1064), .ZN(n152) );
  OAI21_X1 U666 ( .B1(n1072), .B2(n395), .A(n153), .ZN(n853) );
  NAND2_X1 U667 ( .A1(coeffs_ff[17]), .A2(n1063), .ZN(n153) );
  OAI21_X1 U668 ( .B1(n1072), .B2(n396), .A(n154), .ZN(n854) );
  NAND2_X1 U669 ( .A1(coeffs_ff[16]), .A2(n1063), .ZN(n154) );
  OAI21_X1 U670 ( .B1(n1072), .B2(n397), .A(n155), .ZN(n855) );
  NAND2_X1 U671 ( .A1(coeffs_ff[15]), .A2(n1063), .ZN(n155) );
  OAI21_X1 U672 ( .B1(n1072), .B2(n398), .A(n156), .ZN(n856) );
  NAND2_X1 U673 ( .A1(coeffs_ff[14]), .A2(n1063), .ZN(n156) );
  OAI21_X1 U674 ( .B1(n1073), .B2(n399), .A(n157), .ZN(n857) );
  NAND2_X1 U675 ( .A1(coeffs_ff[13]), .A2(n1062), .ZN(n157) );
  OAI21_X1 U676 ( .B1(n1072), .B2(n400), .A(n158), .ZN(n858) );
  NAND2_X1 U677 ( .A1(coeffs_ff[12]), .A2(n1062), .ZN(n158) );
  OAI21_X1 U678 ( .B1(n1072), .B2(n401), .A(n159), .ZN(n859) );
  NAND2_X1 U679 ( .A1(coeffs_ff[11]), .A2(n1062), .ZN(n159) );
  OAI21_X1 U680 ( .B1(n1073), .B2(n402), .A(n160), .ZN(n860) );
  NAND2_X1 U681 ( .A1(coeffs_ff[10]), .A2(n1062), .ZN(n160) );
  OAI21_X1 U682 ( .B1(n1073), .B2(n403), .A(n161), .ZN(n861) );
  NAND2_X1 U683 ( .A1(coeffs_ff[9]), .A2(n1061), .ZN(n161) );
  OAI21_X1 U684 ( .B1(n1073), .B2(n404), .A(n162), .ZN(n862) );
  NAND2_X1 U685 ( .A1(coeffs_ff[8]), .A2(n1061), .ZN(n162) );
  OAI21_X1 U686 ( .B1(n1073), .B2(n405), .A(n163), .ZN(n863) );
  NAND2_X1 U687 ( .A1(coeffs_ff[7]), .A2(n1061), .ZN(n163) );
  OAI21_X1 U688 ( .B1(n1073), .B2(n406), .A(n164), .ZN(n864) );
  NAND2_X1 U689 ( .A1(coeffs_ff[6]), .A2(n1061), .ZN(n164) );
  OAI21_X1 U690 ( .B1(n1073), .B2(n407), .A(n165), .ZN(n865) );
  NAND2_X1 U691 ( .A1(coeffs_ff[5]), .A2(n1060), .ZN(n165) );
  OAI21_X1 U692 ( .B1(n1075), .B2(n408), .A(n166), .ZN(n866) );
  NAND2_X1 U693 ( .A1(coeffs_ff[4]), .A2(n1060), .ZN(n166) );
  OAI21_X1 U694 ( .B1(n1074), .B2(n409), .A(n167), .ZN(n867) );
  NAND2_X1 U695 ( .A1(coeffs_ff[3]), .A2(n1060), .ZN(n167) );
  OAI21_X1 U696 ( .B1(n1074), .B2(n410), .A(n168), .ZN(n868) );
  NAND2_X1 U697 ( .A1(coeffs_ff[2]), .A2(n1060), .ZN(n168) );
  OAI21_X1 U698 ( .B1(n1074), .B2(n411), .A(n169), .ZN(n869) );
  NAND2_X1 U699 ( .A1(coeffs_ff[1]), .A2(n1059), .ZN(n169) );
  OAI21_X1 U700 ( .B1(n1075), .B2(n412), .A(n170), .ZN(n870) );
  NAND2_X1 U701 ( .A1(coeffs_ff[0]), .A2(n1059), .ZN(n170) );
  OAI21_X1 U702 ( .B1(n1075), .B2(n413), .A(n171), .ZN(n871) );
  NAND2_X1 U703 ( .A1(coeffs_ff[47]), .A2(n1059), .ZN(n171) );
  OAI21_X1 U704 ( .B1(n1075), .B2(n414), .A(n172), .ZN(n872) );
  NAND2_X1 U705 ( .A1(coeffs_ff[46]), .A2(n1059), .ZN(n172) );
  OAI21_X1 U706 ( .B1(n1075), .B2(n415), .A(n173), .ZN(n873) );
  NAND2_X1 U707 ( .A1(coeffs_ff[45]), .A2(n1060), .ZN(n173) );
  OAI21_X1 U708 ( .B1(n1078), .B2(n479), .A(n237), .ZN(n937) );
  NAND2_X1 U709 ( .A1(coeffs_ff[77]), .A2(n1070), .ZN(n237) );
  OAI21_X1 U710 ( .B1(n1078), .B2(n480), .A(n238), .ZN(n938) );
  NAND2_X1 U711 ( .A1(coeffs_ff[76]), .A2(n1070), .ZN(n238) );
  OAI21_X1 U712 ( .B1(n1078), .B2(n481), .A(n239), .ZN(n939) );
  NAND2_X1 U713 ( .A1(coeffs_ff[75]), .A2(n1071), .ZN(n239) );
  OAI21_X1 U714 ( .B1(n1078), .B2(n482), .A(n240), .ZN(n940) );
  NAND2_X1 U715 ( .A1(coeffs_ff[74]), .A2(n1071), .ZN(n240) );
  OAI21_X1 U716 ( .B1(n1078), .B2(n483), .A(n241), .ZN(n941) );
  NAND2_X1 U717 ( .A1(coeffs_ff[73]), .A2(n1071), .ZN(n241) );
  OAI21_X1 U718 ( .B1(n1078), .B2(n484), .A(n242), .ZN(n942) );
  NAND2_X1 U719 ( .A1(coeffs_ff[72]), .A2(n1070), .ZN(n242) );
  OAI21_X1 U720 ( .B1(n1078), .B2(n485), .A(n243), .ZN(n943) );
  NAND2_X1 U721 ( .A1(coeffs_fb[23]), .A2(n1070), .ZN(n243) );
  OAI21_X1 U722 ( .B1(n1078), .B2(n486), .A(n244), .ZN(n944) );
  NAND2_X1 U723 ( .A1(coeffs_fb[22]), .A2(n1070), .ZN(n244) );
  OAI21_X1 U724 ( .B1(n1078), .B2(n487), .A(n245), .ZN(n945) );
  NAND2_X1 U725 ( .A1(coeffs_fb[21]), .A2(n1070), .ZN(n245) );
  OAI21_X1 U726 ( .B1(n1078), .B2(n488), .A(n246), .ZN(n946) );
  NAND2_X1 U727 ( .A1(coeffs_fb[20]), .A2(n1070), .ZN(n246) );
  OAI21_X1 U728 ( .B1(n1078), .B2(n489), .A(n247), .ZN(n947) );
  NAND2_X1 U729 ( .A1(coeffs_fb[19]), .A2(n1070), .ZN(n247) );
  OAI21_X1 U730 ( .B1(n1078), .B2(n490), .A(n248), .ZN(n948) );
  NAND2_X1 U731 ( .A1(coeffs_fb[18]), .A2(n1070), .ZN(n248) );
  OAI21_X1 U732 ( .B1(n1078), .B2(n491), .A(n249), .ZN(n949) );
  NAND2_X1 U733 ( .A1(coeffs_fb[17]), .A2(n1069), .ZN(n249) );
  OAI21_X1 U734 ( .B1(n1077), .B2(n492), .A(n250), .ZN(n950) );
  NAND2_X1 U735 ( .A1(coeffs_fb[16]), .A2(n1069), .ZN(n250) );
  OAI21_X1 U736 ( .B1(n1077), .B2(n493), .A(n251), .ZN(n951) );
  NAND2_X1 U737 ( .A1(coeffs_fb[15]), .A2(n1069), .ZN(n251) );
  OAI21_X1 U738 ( .B1(n1077), .B2(n495), .A(n253), .ZN(n953) );
  NAND2_X1 U739 ( .A1(coeffs_fb[13]), .A2(n1069), .ZN(n253) );
  OAI21_X1 U740 ( .B1(n1077), .B2(n496), .A(n254), .ZN(n954) );
  NAND2_X1 U741 ( .A1(coeffs_fb[12]), .A2(n1069), .ZN(n254) );
  OAI21_X1 U742 ( .B1(n1077), .B2(n497), .A(n255), .ZN(n955) );
  NAND2_X1 U743 ( .A1(coeffs_fb[11]), .A2(n1069), .ZN(n255) );
  OAI21_X1 U744 ( .B1(n1077), .B2(n498), .A(n256), .ZN(n956) );
  NAND2_X1 U745 ( .A1(coeffs_fb[10]), .A2(n1068), .ZN(n256) );
  OAI21_X1 U746 ( .B1(n1077), .B2(n499), .A(n257), .ZN(n957) );
  NAND2_X1 U747 ( .A1(coeffs_fb[9]), .A2(n1068), .ZN(n257) );
  OAI21_X1 U748 ( .B1(n1077), .B2(n500), .A(n258), .ZN(n958) );
  NAND2_X1 U749 ( .A1(coeffs_fb[8]), .A2(n1068), .ZN(n258) );
  OAI21_X1 U750 ( .B1(n1077), .B2(n501), .A(n259), .ZN(n959) );
  NAND2_X1 U751 ( .A1(coeffs_fb[7]), .A2(n1068), .ZN(n259) );
  OAI21_X1 U752 ( .B1(n1077), .B2(n502), .A(n260), .ZN(n960) );
  NAND2_X1 U753 ( .A1(coeffs_fb[6]), .A2(n1068), .ZN(n260) );
  OAI21_X1 U754 ( .B1(n1077), .B2(n503), .A(n261), .ZN(n961) );
  NAND2_X1 U755 ( .A1(coeffs_fb[5]), .A2(n1068), .ZN(n261) );
  OAI21_X1 U756 ( .B1(n1077), .B2(n504), .A(n262), .ZN(n962) );
  NAND2_X1 U757 ( .A1(coeffs_fb[4]), .A2(n1068), .ZN(n262) );
  OAI21_X1 U758 ( .B1(n1077), .B2(n505), .A(n263), .ZN(n963) );
  NAND2_X1 U759 ( .A1(coeffs_fb[3]), .A2(n1068), .ZN(n263) );
  OAI21_X1 U760 ( .B1(n1076), .B2(n506), .A(n264), .ZN(n964) );
  NAND2_X1 U761 ( .A1(coeffs_fb[2]), .A2(n1067), .ZN(n264) );
  OAI21_X1 U762 ( .B1(n1076), .B2(n507), .A(n265), .ZN(n965) );
  NAND2_X1 U763 ( .A1(coeffs_fb[1]), .A2(n1067), .ZN(n265) );
  OAI21_X1 U764 ( .B1(n1076), .B2(n508), .A(n266), .ZN(n966) );
  NAND2_X1 U765 ( .A1(coeffs_fb[0]), .A2(n1067), .ZN(n266) );
  OAI21_X1 U766 ( .B1(n1076), .B2(n509), .A(n267), .ZN(n967) );
  NAND2_X1 U767 ( .A1(coeffs_fb[47]), .A2(n1067), .ZN(n267) );
  OAI21_X1 U768 ( .B1(n1076), .B2(n510), .A(n268), .ZN(n968) );
  NAND2_X1 U769 ( .A1(coeffs_fb[46]), .A2(n1067), .ZN(n268) );
  OAI21_X1 U770 ( .B1(n1076), .B2(n511), .A(n269), .ZN(n969) );
  NAND2_X1 U771 ( .A1(coeffs_fb[45]), .A2(n1067), .ZN(n269) );
  OAI21_X1 U772 ( .B1(n1076), .B2(n512), .A(n270), .ZN(n970) );
  NAND2_X1 U773 ( .A1(coeffs_fb[44]), .A2(n1067), .ZN(n270) );
  OAI21_X1 U774 ( .B1(n1076), .B2(n513), .A(n271), .ZN(n971) );
  NAND2_X1 U775 ( .A1(coeffs_fb[43]), .A2(n1067), .ZN(n271) );
  OAI21_X1 U776 ( .B1(n1076), .B2(n514), .A(n272), .ZN(n972) );
  NAND2_X1 U777 ( .A1(coeffs_fb[42]), .A2(n1066), .ZN(n272) );
  OAI21_X1 U778 ( .B1(n1076), .B2(n515), .A(n273), .ZN(n973) );
  NAND2_X1 U779 ( .A1(coeffs_fb[41]), .A2(n1066), .ZN(n273) );
  OAI21_X1 U780 ( .B1(n1076), .B2(n516), .A(n274), .ZN(n974) );
  NAND2_X1 U781 ( .A1(coeffs_fb[40]), .A2(n1066), .ZN(n274) );
  OAI21_X1 U782 ( .B1(n1076), .B2(n517), .A(n275), .ZN(n975) );
  NAND2_X1 U783 ( .A1(coeffs_fb[39]), .A2(n1066), .ZN(n275) );
  OAI21_X1 U784 ( .B1(n1076), .B2(n518), .A(n276), .ZN(n976) );
  NAND2_X1 U785 ( .A1(coeffs_fb[38]), .A2(n1066), .ZN(n276) );
  OAI21_X1 U786 ( .B1(n1074), .B2(n277), .A(n33), .ZN(n978) );
  NAND2_X1 U787 ( .A1(coeffs_fb[36]), .A2(n1066), .ZN(n33) );
  OAI21_X1 U788 ( .B1(n1075), .B2(n278), .A(n34), .ZN(n979) );
  NAND2_X1 U789 ( .A1(coeffs_fb[35]), .A2(n1066), .ZN(n34) );
  OAI21_X1 U790 ( .B1(n1075), .B2(n279), .A(n35), .ZN(n980) );
  NAND2_X1 U791 ( .A1(coeffs_fb[34]), .A2(n1067), .ZN(n35) );
  OAI21_X1 U792 ( .B1(n1075), .B2(n280), .A(n36), .ZN(n981) );
  NAND2_X1 U793 ( .A1(coeffs_fb[33]), .A2(n1067), .ZN(n36) );
  OAI21_X1 U794 ( .B1(n1074), .B2(n281), .A(n37), .ZN(n982) );
  NAND2_X1 U795 ( .A1(coeffs_fb[32]), .A2(n1067), .ZN(n37) );
  OAI21_X1 U796 ( .B1(n1074), .B2(n282), .A(n38), .ZN(n983) );
  NAND2_X1 U797 ( .A1(coeffs_fb[31]), .A2(n1067), .ZN(n38) );
  OAI21_X1 U798 ( .B1(n1074), .B2(n283), .A(n39), .ZN(n984) );
  NAND2_X1 U799 ( .A1(coeffs_fb[30]), .A2(n1068), .ZN(n39) );
  OAI21_X1 U800 ( .B1(n1073), .B2(n284), .A(n40), .ZN(n985) );
  NAND2_X1 U801 ( .A1(coeffs_fb[29]), .A2(n1068), .ZN(n40) );
  OAI21_X1 U802 ( .B1(n1073), .B2(n285), .A(n41), .ZN(n986) );
  NAND2_X1 U803 ( .A1(coeffs_fb[28]), .A2(n1068), .ZN(n41) );
  OAI21_X1 U804 ( .B1(n1073), .B2(n286), .A(n42), .ZN(n987) );
  NAND2_X1 U805 ( .A1(coeffs_fb[27]), .A2(n1068), .ZN(n42) );
  OAI21_X1 U806 ( .B1(n1072), .B2(n287), .A(n43), .ZN(n988) );
  NAND2_X1 U807 ( .A1(coeffs_fb[26]), .A2(n1069), .ZN(n43) );
  OAI21_X1 U808 ( .B1(n1072), .B2(n288), .A(n44), .ZN(n989) );
  NAND2_X1 U809 ( .A1(coeffs_fb[25]), .A2(n1069), .ZN(n44) );
  OAI21_X1 U810 ( .B1(n1072), .B2(n289), .A(n45), .ZN(n990) );
  NAND2_X1 U811 ( .A1(coeffs_fb[24]), .A2(n1069), .ZN(n45) );
  OAI21_X1 U812 ( .B1(n1072), .B2(n290), .A(n46), .ZN(n991) );
  NAND2_X1 U813 ( .A1(dIn[11]), .A2(n1069), .ZN(n46) );
  OAI21_X1 U814 ( .B1(n1072), .B2(n292), .A(n48), .ZN(n993) );
  NAND2_X1 U815 ( .A1(dIn[9]), .A2(n1070), .ZN(n48) );
  OAI21_X1 U816 ( .B1(n1072), .B2(n293), .A(n49), .ZN(n994) );
  NAND2_X1 U817 ( .A1(dIn[8]), .A2(n1070), .ZN(n49) );
  OAI21_X1 U818 ( .B1(n1074), .B2(n294), .A(n50), .ZN(n995) );
  NAND2_X1 U819 ( .A1(dIn[7]), .A2(n1071), .ZN(n50) );
  OAI21_X1 U820 ( .B1(n1074), .B2(n295), .A(n51), .ZN(n996) );
  NAND2_X1 U821 ( .A1(dIn[6]), .A2(n1071), .ZN(n51) );
  OAI21_X1 U822 ( .B1(n1074), .B2(n296), .A(n52), .ZN(n997) );
  NAND2_X1 U823 ( .A1(dIn[5]), .A2(n1069), .ZN(n52) );
  OAI21_X1 U824 ( .B1(n1074), .B2(n297), .A(n53), .ZN(n998) );
  NAND2_X1 U825 ( .A1(dIn[4]), .A2(n1071), .ZN(n53) );
  OAI21_X1 U826 ( .B1(n1075), .B2(n298), .A(n54), .ZN(n999) );
  NAND2_X1 U827 ( .A1(dIn[3]), .A2(n1071), .ZN(n54) );
  OAI21_X1 U828 ( .B1(n1075), .B2(n299), .A(n55), .ZN(n1000) );
  NAND2_X1 U829 ( .A1(dIn[2]), .A2(n1066), .ZN(n55) );
  OAI21_X1 U830 ( .B1(n1075), .B2(n300), .A(n56), .ZN(n1001) );
  NAND2_X1 U831 ( .A1(dIn[1]), .A2(n1065), .ZN(n56) );
  OAI21_X1 U832 ( .B1(n1075), .B2(n301), .A(n57), .ZN(n1002) );
  NAND2_X1 U833 ( .A1(dIn[0]), .A2(n1065), .ZN(n57) );
  OAI21_X1 U834 ( .B1(n1071), .B2(n291), .A(n47), .ZN(n992) );
  NAND2_X1 U835 ( .A1(dIn[10]), .A2(n1070), .ZN(n47) );
  OAI21_X1 U836 ( .B1(n1082), .B2(n428), .A(n186), .ZN(n886) );
  NAND2_X1 U837 ( .A1(coeffs_ff[32]), .A2(n1066), .ZN(n186) );
  OAI21_X1 U838 ( .B1(n1082), .B2(n429), .A(n187), .ZN(n887) );
  NAND2_X1 U839 ( .A1(coeffs_ff[31]), .A2(n1060), .ZN(n187) );
  OAI21_X1 U840 ( .B1(n1082), .B2(n430), .A(n188), .ZN(n888) );
  NAND2_X1 U841 ( .A1(coeffs_ff[30]), .A2(n1060), .ZN(n188) );
  OAI21_X1 U842 ( .B1(n1082), .B2(n431), .A(n189), .ZN(n889) );
  NAND2_X1 U843 ( .A1(coeffs_ff[29]), .A2(n1060), .ZN(n189) );
  OAI21_X1 U844 ( .B1(n1082), .B2(n432), .A(n190), .ZN(n890) );
  NAND2_X1 U845 ( .A1(coeffs_ff[28]), .A2(n1061), .ZN(n190) );
  OAI21_X1 U846 ( .B1(n1082), .B2(n433), .A(n191), .ZN(n891) );
  NAND2_X1 U847 ( .A1(coeffs_ff[27]), .A2(n1061), .ZN(n191) );
  OAI21_X1 U848 ( .B1(n1082), .B2(n434), .A(n192), .ZN(n892) );
  NAND2_X1 U849 ( .A1(coeffs_ff[26]), .A2(n1061), .ZN(n192) );
  OAI21_X1 U850 ( .B1(n1082), .B2(n435), .A(n193), .ZN(n893) );
  NAND2_X1 U851 ( .A1(coeffs_ff[25]), .A2(n1061), .ZN(n193) );
  OAI21_X1 U852 ( .B1(n1082), .B2(n436), .A(n194), .ZN(n894) );
  NAND2_X1 U853 ( .A1(coeffs_ff[24]), .A2(n1061), .ZN(n194) );
  OAI21_X1 U854 ( .B1(n1082), .B2(n437), .A(n195), .ZN(n895) );
  NAND2_X1 U855 ( .A1(coeffs_ff[71]), .A2(n1061), .ZN(n195) );
  OAI21_X1 U856 ( .B1(n1082), .B2(n438), .A(n196), .ZN(n896) );
  NAND2_X1 U857 ( .A1(coeffs_ff[70]), .A2(n1061), .ZN(n196) );
  OAI21_X1 U858 ( .B1(n1082), .B2(n439), .A(n197), .ZN(n897) );
  NAND2_X1 U859 ( .A1(coeffs_ff[69]), .A2(n1061), .ZN(n197) );
  OAI21_X1 U860 ( .B1(n1082), .B2(n440), .A(n198), .ZN(n898) );
  NAND2_X1 U861 ( .A1(coeffs_ff[68]), .A2(n1062), .ZN(n198) );
  OAI21_X1 U862 ( .B1(n1081), .B2(n441), .A(n199), .ZN(n899) );
  NAND2_X1 U863 ( .A1(coeffs_ff[67]), .A2(n1062), .ZN(n199) );
  OAI21_X1 U864 ( .B1(n1081), .B2(n442), .A(n200), .ZN(n900) );
  NAND2_X1 U865 ( .A1(coeffs_ff[66]), .A2(n1062), .ZN(n200) );
  OAI21_X1 U866 ( .B1(n1081), .B2(n443), .A(n201), .ZN(n901) );
  NAND2_X1 U867 ( .A1(coeffs_ff[65]), .A2(n1062), .ZN(n201) );
  OAI21_X1 U868 ( .B1(n1081), .B2(n444), .A(n202), .ZN(n902) );
  NAND2_X1 U869 ( .A1(coeffs_ff[64]), .A2(n1062), .ZN(n202) );
  OAI21_X1 U870 ( .B1(n1081), .B2(n445), .A(n203), .ZN(n903) );
  NAND2_X1 U871 ( .A1(coeffs_ff[63]), .A2(n1062), .ZN(n203) );
  OAI21_X1 U872 ( .B1(n1081), .B2(n446), .A(n204), .ZN(n904) );
  NAND2_X1 U873 ( .A1(coeffs_ff[62]), .A2(n1062), .ZN(n204) );
  OAI21_X1 U874 ( .B1(n1081), .B2(n447), .A(n205), .ZN(n905) );
  NAND2_X1 U875 ( .A1(coeffs_ff[61]), .A2(n1062), .ZN(n205) );
  OAI21_X1 U876 ( .B1(n1081), .B2(n448), .A(n206), .ZN(n906) );
  NAND2_X1 U877 ( .A1(coeffs_ff[60]), .A2(n1063), .ZN(n206) );
  OAI21_X1 U878 ( .B1(n1081), .B2(n449), .A(n207), .ZN(n907) );
  NAND2_X1 U879 ( .A1(coeffs_ff[59]), .A2(n1063), .ZN(n207) );
  OAI21_X1 U880 ( .B1(n1081), .B2(n450), .A(n208), .ZN(n908) );
  NAND2_X1 U881 ( .A1(coeffs_ff[58]), .A2(n1063), .ZN(n208) );
  OAI21_X1 U882 ( .B1(n1081), .B2(n451), .A(n209), .ZN(n909) );
  NAND2_X1 U883 ( .A1(coeffs_ff[57]), .A2(n1063), .ZN(n209) );
  OAI21_X1 U884 ( .B1(n1081), .B2(n452), .A(n210), .ZN(n910) );
  NAND2_X1 U885 ( .A1(coeffs_ff[56]), .A2(n1063), .ZN(n210) );
  OAI21_X1 U886 ( .B1(n1081), .B2(n453), .A(n211), .ZN(n911) );
  NAND2_X1 U887 ( .A1(coeffs_ff[55]), .A2(n1063), .ZN(n211) );
  OAI21_X1 U888 ( .B1(n1080), .B2(n454), .A(n212), .ZN(n912) );
  NAND2_X1 U889 ( .A1(coeffs_ff[54]), .A2(n1063), .ZN(n212) );
  OAI21_X1 U890 ( .B1(n1080), .B2(n455), .A(n213), .ZN(n913) );
  NAND2_X1 U891 ( .A1(coeffs_ff[53]), .A2(n1063), .ZN(n213) );
  OAI21_X1 U892 ( .B1(n1080), .B2(n456), .A(n214), .ZN(n914) );
  NAND2_X1 U893 ( .A1(coeffs_ff[52]), .A2(n1064), .ZN(n214) );
  OAI21_X1 U894 ( .B1(n1080), .B2(n457), .A(n215), .ZN(n915) );
  NAND2_X1 U895 ( .A1(coeffs_ff[51]), .A2(n1064), .ZN(n215) );
  OAI21_X1 U896 ( .B1(n1080), .B2(n458), .A(n216), .ZN(n916) );
  NAND2_X1 U897 ( .A1(coeffs_ff[50]), .A2(n1064), .ZN(n216) );
  OAI21_X1 U898 ( .B1(n1080), .B2(n459), .A(n217), .ZN(n917) );
  NAND2_X1 U899 ( .A1(coeffs_ff[49]), .A2(n1064), .ZN(n217) );
  OAI21_X1 U900 ( .B1(n1080), .B2(n460), .A(n218), .ZN(n918) );
  NAND2_X1 U901 ( .A1(coeffs_ff[48]), .A2(n1064), .ZN(n218) );
  OAI21_X1 U902 ( .B1(n1080), .B2(n461), .A(n219), .ZN(n919) );
  NAND2_X1 U903 ( .A1(coeffs_ff[95]), .A2(n1064), .ZN(n219) );
  OAI21_X1 U904 ( .B1(n1080), .B2(n462), .A(n220), .ZN(n920) );
  NAND2_X1 U905 ( .A1(coeffs_ff[94]), .A2(n1064), .ZN(n220) );
  OAI21_X1 U906 ( .B1(n1080), .B2(n463), .A(n221), .ZN(n921) );
  NAND2_X1 U907 ( .A1(coeffs_ff[93]), .A2(n1064), .ZN(n221) );
  OAI21_X1 U908 ( .B1(n1080), .B2(n464), .A(n222), .ZN(n922) );
  NAND2_X1 U909 ( .A1(coeffs_ff[92]), .A2(n1065), .ZN(n222) );
  OAI21_X1 U910 ( .B1(n1080), .B2(n465), .A(n223), .ZN(n923) );
  NAND2_X1 U911 ( .A1(coeffs_ff[91]), .A2(n1065), .ZN(n223) );
  OAI21_X1 U912 ( .B1(n1080), .B2(n466), .A(n224), .ZN(n924) );
  NAND2_X1 U913 ( .A1(coeffs_ff[90]), .A2(n1065), .ZN(n224) );
  OAI21_X1 U914 ( .B1(n1079), .B2(n467), .A(n225), .ZN(n925) );
  NAND2_X1 U915 ( .A1(coeffs_ff[89]), .A2(n1065), .ZN(n225) );
  OAI21_X1 U916 ( .B1(n1079), .B2(n468), .A(n226), .ZN(n926) );
  NAND2_X1 U917 ( .A1(coeffs_ff[88]), .A2(n1065), .ZN(n226) );
  OAI21_X1 U918 ( .B1(n1079), .B2(n469), .A(n227), .ZN(n927) );
  NAND2_X1 U919 ( .A1(coeffs_ff[87]), .A2(n1065), .ZN(n227) );
  OAI21_X1 U920 ( .B1(n1079), .B2(n470), .A(n228), .ZN(n928) );
  NAND2_X1 U921 ( .A1(coeffs_ff[86]), .A2(n1065), .ZN(n228) );
  OAI21_X1 U922 ( .B1(n1079), .B2(n471), .A(n229), .ZN(n929) );
  NAND2_X1 U923 ( .A1(coeffs_ff[85]), .A2(n1065), .ZN(n229) );
  OAI21_X1 U924 ( .B1(n1079), .B2(n472), .A(n230), .ZN(n930) );
  NAND2_X1 U925 ( .A1(coeffs_ff[84]), .A2(n1066), .ZN(n230) );
  OAI21_X1 U926 ( .B1(n1079), .B2(n473), .A(n231), .ZN(n931) );
  NAND2_X1 U927 ( .A1(coeffs_ff[83]), .A2(n1066), .ZN(n231) );
  OAI21_X1 U928 ( .B1(n1079), .B2(n474), .A(n232), .ZN(n932) );
  NAND2_X1 U929 ( .A1(coeffs_ff[82]), .A2(n1066), .ZN(n232) );
  OAI21_X1 U930 ( .B1(n1079), .B2(n475), .A(n233), .ZN(n933) );
  NAND2_X1 U931 ( .A1(coeffs_ff[81]), .A2(n1071), .ZN(n233) );
  OAI21_X1 U932 ( .B1(n1079), .B2(n476), .A(n234), .ZN(n934) );
  NAND2_X1 U933 ( .A1(coeffs_ff[80]), .A2(n1071), .ZN(n234) );
  OAI21_X1 U934 ( .B1(n1079), .B2(n477), .A(n235), .ZN(n935) );
  NAND2_X1 U935 ( .A1(coeffs_ff[79]), .A2(n1071), .ZN(n235) );
  OAI21_X1 U936 ( .B1(n1079), .B2(n478), .A(n236), .ZN(n936) );
  NAND2_X1 U937 ( .A1(coeffs_ff[78]), .A2(n1071), .ZN(n236) );
  OAI21_X1 U938 ( .B1(n1079), .B2(n494), .A(n252), .ZN(n952) );
  NAND2_X1 U939 ( .A1(coeffs_fb[14]), .A2(n1069), .ZN(n252) );
  OAI21_X1 U940 ( .B1(n1083), .B2(n416), .A(n174), .ZN(n874) );
  NAND2_X1 U941 ( .A1(coeffs_ff[44]), .A2(n1059), .ZN(n174) );
  OAI21_X1 U942 ( .B1(n1083), .B2(n417), .A(n175), .ZN(n875) );
  NAND2_X1 U943 ( .A1(coeffs_ff[43]), .A2(n1059), .ZN(n175) );
  OAI21_X1 U944 ( .B1(n1083), .B2(n418), .A(n176), .ZN(n876) );
  NAND2_X1 U945 ( .A1(coeffs_ff[42]), .A2(n1059), .ZN(n176) );
  OAI21_X1 U946 ( .B1(n1083), .B2(n419), .A(n177), .ZN(n877) );
  NAND2_X1 U947 ( .A1(coeffs_ff[41]), .A2(n1059), .ZN(n177) );
  OAI21_X1 U948 ( .B1(n1083), .B2(n420), .A(n178), .ZN(n878) );
  NAND2_X1 U949 ( .A1(coeffs_ff[40]), .A2(n1059), .ZN(n178) );
  OAI21_X1 U950 ( .B1(n1083), .B2(n421), .A(n179), .ZN(n879) );
  NAND2_X1 U951 ( .A1(coeffs_ff[39]), .A2(n1059), .ZN(n179) );
  OAI21_X1 U952 ( .B1(n1083), .B2(n422), .A(n180), .ZN(n880) );
  NAND2_X1 U953 ( .A1(coeffs_ff[38]), .A2(n1059), .ZN(n180) );
  OAI21_X1 U954 ( .B1(n1083), .B2(n423), .A(n181), .ZN(n881) );
  NAND2_X1 U955 ( .A1(coeffs_ff[37]), .A2(n1059), .ZN(n181) );
  OAI21_X1 U956 ( .B1(n1083), .B2(n424), .A(n182), .ZN(n882) );
  NAND2_X1 U957 ( .A1(coeffs_ff[36]), .A2(n1060), .ZN(n182) );
  OAI21_X1 U958 ( .B1(n1083), .B2(n425), .A(n183), .ZN(n883) );
  NAND2_X1 U959 ( .A1(coeffs_ff[35]), .A2(n1060), .ZN(n183) );
  OAI21_X1 U960 ( .B1(n1083), .B2(n426), .A(n184), .ZN(n884) );
  NAND2_X1 U961 ( .A1(coeffs_ff[34]), .A2(n1060), .ZN(n184) );
  OAI21_X1 U962 ( .B1(n1083), .B2(n427), .A(n185), .ZN(n885) );
  NAND2_X1 U963 ( .A1(coeffs_ff[33]), .A2(n1060), .ZN(n185) );
  OAI21_X1 U964 ( .B1(n1075), .B2(n519), .A(n32), .ZN(n977) );
  NAND2_X1 U965 ( .A1(n1083), .A2(coeffs_fb[37]), .ZN(n32) );
  BUF_X1 U966 ( .A(vIn), .Z(n1089) );
  BUF_X1 U967 ( .A(vIn), .Z(n1090) );
  INV_X1 U968 ( .A(n103), .ZN(n716) );
  AOI22_X1 U969 ( .A1(n1033), .A2(DP_sw0_21_), .B1(n1048), .B2(DP_sw1_21_), 
        .ZN(n103) );
  INV_X1 U970 ( .A(n105), .ZN(n721) );
  AOI22_X1 U971 ( .A1(n1034), .A2(DP_sw0_20_), .B1(n1048), .B2(DP_sw1_20_), 
        .ZN(n105) );
  INV_X1 U972 ( .A(n107), .ZN(n726) );
  AOI22_X1 U973 ( .A1(n1034), .A2(DP_sw0_19_), .B1(n1047), .B2(DP_sw1_19_), 
        .ZN(n107) );
  INV_X1 U974 ( .A(n109), .ZN(n731) );
  AOI22_X1 U975 ( .A1(n1033), .A2(DP_sw0_18_), .B1(n1047), .B2(DP_sw1_18_), 
        .ZN(n109) );
  INV_X1 U976 ( .A(n111), .ZN(n736) );
  AOI22_X1 U977 ( .A1(n1032), .A2(DP_sw0_17_), .B1(n1046), .B2(DP_sw1_17_), 
        .ZN(n111) );
  INV_X1 U978 ( .A(n101), .ZN(n711) );
  AOI22_X1 U979 ( .A1(n1033), .A2(DP_sw0_22_), .B1(n1048), .B2(DP_sw1_22_), 
        .ZN(n101) );
  INV_X1 U980 ( .A(n113), .ZN(n741) );
  AOI22_X1 U981 ( .A1(n1033), .A2(DP_sw0_16_), .B1(n1046), .B2(DP_sw1_16_), 
        .ZN(n113) );
  INV_X1 U982 ( .A(n115), .ZN(n746) );
  AOI22_X1 U983 ( .A1(n1034), .A2(DP_sw0_15_), .B1(n1046), .B2(DP_sw1_15_), 
        .ZN(n115) );
  INV_X1 U984 ( .A(n117), .ZN(n751) );
  AOI22_X1 U985 ( .A1(n1032), .A2(DP_sw0_14_), .B1(n1045), .B2(DP_sw1_14_), 
        .ZN(n117) );
  INV_X1 U986 ( .A(n119), .ZN(n756) );
  AOI22_X1 U987 ( .A1(n1032), .A2(DP_sw0_13_), .B1(n1045), .B2(DP_sw1_13_), 
        .ZN(n119) );
  INV_X1 U988 ( .A(n121), .ZN(n761) );
  AOI22_X1 U989 ( .A1(n1033), .A2(DP_sw0_12_), .B1(n1044), .B2(DP_sw1_12_), 
        .ZN(n121) );
  INV_X1 U990 ( .A(n125), .ZN(n771) );
  AOI22_X1 U991 ( .A1(n1033), .A2(DP_sw0_10_), .B1(n1043), .B2(DP_sw1_10_), 
        .ZN(n125) );
  INV_X1 U992 ( .A(n127), .ZN(n776) );
  AOI22_X1 U993 ( .A1(n1033), .A2(DP_sw0_9_), .B1(n1043), .B2(DP_sw1_9_), .ZN(
        n127) );
  INV_X1 U994 ( .A(n129), .ZN(n781) );
  AOI22_X1 U995 ( .A1(n1033), .A2(DP_sw0_8_), .B1(n1043), .B2(DP_sw1_8_), .ZN(
        n129) );
  INV_X1 U996 ( .A(n131), .ZN(n786) );
  AOI22_X1 U997 ( .A1(n1033), .A2(DP_sw0_7_), .B1(n1042), .B2(DP_sw1_7_), .ZN(
        n131) );
  INV_X1 U998 ( .A(n133), .ZN(n791) );
  AOI22_X1 U999 ( .A1(n1033), .A2(DP_sw0_6_), .B1(n1042), .B2(DP_sw1_6_), .ZN(
        n133) );
  INV_X1 U1000 ( .A(n135), .ZN(n796) );
  AOI22_X1 U1001 ( .A1(n1033), .A2(DP_sw0_5_), .B1(n1042), .B2(DP_sw1_5_), 
        .ZN(n135) );
  INV_X1 U1002 ( .A(n145), .ZN(n820) );
  AOI22_X1 U1003 ( .A1(n1034), .A2(DP_w_0_), .B1(n1041), .B2(DP_sw0_0_), .ZN(
        n145) );
  INV_X1 U1004 ( .A(n140), .ZN(n807) );
  AOI22_X1 U1005 ( .A1(n1034), .A2(DP_w_3_), .B1(n1040), .B2(DP_sw0_3_), .ZN(
        n140) );
  INV_X1 U1006 ( .A(n142), .ZN(n812) );
  AOI22_X1 U1007 ( .A1(n1034), .A2(DP_w_2_), .B1(n1040), .B2(DP_sw0_2_), .ZN(
        n142) );
  INV_X1 U1008 ( .A(n144), .ZN(n817) );
  AOI22_X1 U1009 ( .A1(n1034), .A2(DP_w_1_), .B1(n1040), .B2(DP_sw0_1_), .ZN(
        n144) );
  INV_X1 U1010 ( .A(n99), .ZN(n706) );
  AOI22_X1 U1011 ( .A1(n1034), .A2(DP_sw0_23_), .B1(n1049), .B2(DP_sw1_23_), 
        .ZN(n99) );
  INV_X1 U1012 ( .A(n123), .ZN(n766) );
  AOI22_X1 U1013 ( .A1(n1034), .A2(DP_sw0_11_), .B1(n1044), .B2(DP_sw1_11_), 
        .ZN(n123) );
  INV_X1 U1014 ( .A(n137), .ZN(n801) );
  AOI22_X1 U1015 ( .A1(n1034), .A2(DP_sw0_4_), .B1(n1041), .B2(DP_sw1_4_), 
        .ZN(n137) );
  INV_X1 U1016 ( .A(n139), .ZN(n806) );
  AOI22_X1 U1017 ( .A1(n1034), .A2(DP_sw0_3_), .B1(n1041), .B2(DP_sw1_3_), 
        .ZN(n139) );
  INV_X1 U1018 ( .A(n141), .ZN(n811) );
  AOI22_X1 U1019 ( .A1(n1034), .A2(DP_sw0_2_), .B1(n1040), .B2(DP_sw1_2_), 
        .ZN(n141) );
  INV_X1 U1020 ( .A(n143), .ZN(n816) );
  AOI22_X1 U1021 ( .A1(n1034), .A2(DP_sw0_1_), .B1(n1040), .B2(DP_sw1_1_), 
        .ZN(n143) );
  BUF_X1 U1022 ( .A(rst_n), .Z(n1132) );
  BUF_X1 U1023 ( .A(rst_n), .Z(n1133) );
  BUF_X1 U1024 ( .A(rst_n), .Z(n1134) );
  BUF_X1 U1025 ( .A(rst_n), .Z(n1135) );
  BUF_X1 U1026 ( .A(rst_n), .Z(n1136) );
  BUF_X1 U1027 ( .A(rst_n), .Z(n1137) );
  BUF_X1 U1028 ( .A(rst_n), .Z(n1138) );
  INV_X1 U1029 ( .A(n1049), .ZN(n1032) );
  INV_X1 U1030 ( .A(n1050), .ZN(n1034) );
  CLKBUF_X1 U1031 ( .A(n1138), .Z(n1091) );
  CLKBUF_X1 U1032 ( .A(n1138), .Z(n1092) );
  CLKBUF_X1 U1033 ( .A(n1138), .Z(n1093) );
  CLKBUF_X1 U1034 ( .A(n1138), .Z(n1094) );
  CLKBUF_X1 U1035 ( .A(n1138), .Z(n1095) );
  CLKBUF_X1 U1036 ( .A(n1137), .Z(n1096) );
  CLKBUF_X1 U1037 ( .A(n1137), .Z(n1097) );
  CLKBUF_X1 U1038 ( .A(n1137), .Z(n1098) );
  CLKBUF_X1 U1039 ( .A(n1137), .Z(n1099) );
  CLKBUF_X1 U1040 ( .A(n1137), .Z(n1100) );
  CLKBUF_X1 U1041 ( .A(n1137), .Z(n1101) );
  CLKBUF_X1 U1042 ( .A(n1136), .Z(n1102) );
  CLKBUF_X1 U1043 ( .A(n1136), .Z(n1103) );
  CLKBUF_X1 U1044 ( .A(n1136), .Z(n1104) );
  CLKBUF_X1 U1045 ( .A(n1136), .Z(n1105) );
  CLKBUF_X1 U1046 ( .A(n1136), .Z(n1106) );
  CLKBUF_X1 U1047 ( .A(n1136), .Z(n1107) );
  CLKBUF_X1 U1048 ( .A(n1135), .Z(n1108) );
  CLKBUF_X1 U1049 ( .A(n1135), .Z(n1109) );
  CLKBUF_X1 U1050 ( .A(n1135), .Z(n1110) );
  CLKBUF_X1 U1051 ( .A(n1135), .Z(n1111) );
  CLKBUF_X1 U1052 ( .A(n1135), .Z(n1112) );
  CLKBUF_X1 U1053 ( .A(n1135), .Z(n1113) );
  CLKBUF_X1 U1054 ( .A(n1134), .Z(n1114) );
  CLKBUF_X1 U1055 ( .A(n1134), .Z(n1115) );
  CLKBUF_X1 U1056 ( .A(n1134), .Z(n1116) );
  CLKBUF_X1 U1057 ( .A(n1134), .Z(n1117) );
  CLKBUF_X1 U1058 ( .A(n1134), .Z(n1118) );
  CLKBUF_X1 U1059 ( .A(n1134), .Z(n1119) );
  CLKBUF_X1 U1060 ( .A(n1133), .Z(n1120) );
  CLKBUF_X1 U1061 ( .A(n1133), .Z(n1121) );
  CLKBUF_X1 U1062 ( .A(n1133), .Z(n1122) );
  CLKBUF_X1 U1063 ( .A(n1133), .Z(n1123) );
  CLKBUF_X1 U1064 ( .A(n1133), .Z(n1124) );
  CLKBUF_X1 U1065 ( .A(n1133), .Z(n1125) );
  CLKBUF_X1 U1066 ( .A(n1132), .Z(n1126) );
  CLKBUF_X1 U1067 ( .A(n1132), .Z(n1127) );
  CLKBUF_X1 U1068 ( .A(n1132), .Z(n1128) );
  CLKBUF_X1 U1069 ( .A(n1132), .Z(n1129) );
  CLKBUF_X1 U1070 ( .A(n1132), .Z(n1130) );
  CLKBUF_X1 U1071 ( .A(n1132), .Z(n1131) );
  INV_X1 U1072 ( .A(DP_y_23), .ZN(n1139) );
  NOR2_X1 U1073 ( .A1(DP_y_11_), .A2(n1139), .ZN(DP_N4) );
  INV_X1 U1074 ( .A(DP_y_11_), .ZN(n1140) );
  NOR2_X1 U1075 ( .A1(DP_y_23), .A2(n1140), .ZN(DP_N2) );
endmodule

