
module iir_filter_DW_mult_tc_5 ( a, b, product );
  input [23:0] a;
  input [23:0] b;
  output [47:0] product;
  wire   n251, n293, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n325, n326, n327, n332, n333, n334, n335, n336, n337, n339,
         n341, n342, n343, n344, n345, n346, n347, n348, n350, n352, n353,
         n354, n355, n356, n359, n360, n361, n362, n363, n364, n365, n367,
         n369, n370, n371, n372, n376, n378, n379, n380, n381, n382, n383,
         n384, n387, n388, n389, n390, n394, n396, n397, n398, n399, n400,
         n401, n402, n405, n407, n409, n410, n411, n412, n416, n418, n419,
         n420, n421, n422, n423, n426, n427, n428, n429, n430, n431, n432,
         n434, n435, n436, n437, n438, n439, n445, n450, n451, n452, n453,
         n454, n455, n456, n457, n459, n461, n462, n463, n464, n465, n466,
         n467, n468, n474, n475, n476, n477, n478, n479, n480, n481, n483,
         n486, n487, n488, n489, n490, n492, n495, n496, n497, n498, n499,
         n501, n502, n503, n504, n505, n506, n507, n508, n511, n512, n513,
         n514, n515, n516, n517, n519, n520, n521, n522, n524, n525, n526,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n550, n551, n552, n553, n554,
         n555, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n581, n582, n583, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n609,
         n610, n611, n620, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n643, n644, n645, n646, n657,
         n661, n662, n663, n666, n667, n668, n670, n671, n673, n674, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1817, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376;

  FA_X1 U546 ( .A(n1195), .B(n682), .CI(n1218), .CO(n678), .S(n679) );
  FA_X1 U547 ( .A(n683), .B(n1196), .CI(n686), .CO(n680), .S(n681) );
  FA_X1 U549 ( .A(n690), .B(n1242), .CI(n687), .CO(n684), .S(n685) );
  FA_X1 U550 ( .A(n1219), .B(n692), .CI(n1197), .CO(n686), .S(n687) );
  FA_X1 U551 ( .A(n691), .B(n698), .CI(n696), .CO(n688), .S(n689) );
  FA_X1 U552 ( .A(n1198), .B(n1220), .CI(n693), .CO(n690), .S(n691) );
  FA_X1 U554 ( .A(n702), .B(n699), .CI(n697), .CO(n694), .S(n695) );
  FA_X1 U555 ( .A(n1266), .B(n1243), .CI(n704), .CO(n696), .S(n697) );
  FA_X1 U556 ( .A(n1221), .B(n1199), .CI(n706), .CO(n698), .S(n699) );
  FA_X1 U557 ( .A(n710), .B(n712), .CI(n703), .CO(n700), .S(n701) );
  FA_X1 U558 ( .A(n714), .B(n1244), .CI(n705), .CO(n702), .S(n703) );
  FA_X1 U559 ( .A(n1222), .B(n1200), .CI(n707), .CO(n704), .S(n705) );
  FA_X1 U561 ( .A(n718), .B(n713), .CI(n711), .CO(n708), .S(n709) );
  FA_X1 U562 ( .A(n715), .B(n722), .CI(n720), .CO(n710), .S(n711) );
  FA_X1 U563 ( .A(n1245), .B(n1223), .CI(n1290), .CO(n712), .S(n713) );
  FA_X1 U564 ( .A(n1267), .B(n1201), .CI(n724), .CO(n714), .S(n715) );
  FA_X1 U565 ( .A(n728), .B(n721), .CI(n719), .CO(n716), .S(n717) );
  FA_X1 U566 ( .A(n723), .B(n732), .CI(n730), .CO(n718), .S(n719) );
  FA_X1 U567 ( .A(n1202), .B(n1246), .CI(n734), .CO(n720), .S(n721) );
  FA_X1 U568 ( .A(n1268), .B(n1224), .CI(n725), .CO(n722), .S(n723) );
  FA_X1 U570 ( .A(n738), .B(n731), .CI(n729), .CO(n726), .S(n727) );
  FA_X1 U571 ( .A(n735), .B(n733), .CI(n740), .CO(n728), .S(n729) );
  FA_X1 U572 ( .A(n744), .B(n1314), .CI(n742), .CO(n730), .S(n731) );
  FA_X1 U573 ( .A(n1225), .B(n1291), .CI(n1269), .CO(n732), .S(n733) );
  FA_X1 U574 ( .A(n746), .B(n1203), .CI(n1247), .CO(n734), .S(n735) );
  FA_X1 U575 ( .A(n750), .B(n741), .CI(n739), .CO(n736), .S(n737) );
  FA_X1 U576 ( .A(n754), .B(n745), .CI(n752), .CO(n738), .S(n739) );
  FA_X1 U577 ( .A(n756), .B(n758), .CI(n743), .CO(n740), .S(n741) );
  FA_X1 U578 ( .A(n1226), .B(n1270), .CI(n1204), .CO(n742), .S(n743) );
  FA_X1 U579 ( .A(n1292), .B(n1248), .CI(n747), .CO(n744), .S(n745) );
  FA_X1 U581 ( .A(n762), .B(n753), .CI(n751), .CO(n748), .S(n749) );
  FA_X1 U582 ( .A(n755), .B(n766), .CI(n764), .CO(n750), .S(n751) );
  FA_X1 U583 ( .A(n757), .B(n768), .CI(n759), .CO(n752), .S(n753) );
  FA_X1 U584 ( .A(n1338), .B(n1271), .CI(n770), .CO(n754), .S(n755) );
  FA_X1 U585 ( .A(n1249), .B(n1293), .CI(n1315), .CO(n756), .S(n757) );
  FA_X1 U586 ( .A(n772), .B(n1205), .CI(n1227), .CO(n758), .S(n759) );
  FA_X1 U587 ( .A(n776), .B(n765), .CI(n763), .CO(n760), .S(n761) );
  FA_X1 U588 ( .A(n767), .B(n780), .CI(n778), .CO(n762), .S(n763) );
  FA_X1 U589 ( .A(n771), .B(n769), .CI(n782), .CO(n764), .S(n765) );
  FA_X1 U590 ( .A(n786), .B(n1228), .CI(n784), .CO(n766), .S(n767) );
  FA_X1 U591 ( .A(n1294), .B(n1206), .CI(n1272), .CO(n768), .S(n769) );
  FA_X1 U592 ( .A(n1316), .B(n1250), .CI(n773), .CO(n770), .S(n771) );
  FA_X1 U594 ( .A(n790), .B(n779), .CI(n777), .CO(n774), .S(n775) );
  FA_X1 U595 ( .A(n781), .B(n794), .CI(n792), .CO(n776), .S(n777) );
  FA_X1 U596 ( .A(n796), .B(n787), .CI(n783), .CO(n778), .S(n779) );
  FA_X1 U597 ( .A(n798), .B(n800), .CI(n785), .CO(n780), .S(n781) );
  FA_X1 U598 ( .A(n1339), .B(n1229), .CI(n1362), .CO(n782), .S(n783) );
  FA_X1 U599 ( .A(n1273), .B(n1317), .CI(n1295), .CO(n784), .S(n785) );
  FA_X1 U600 ( .A(n802), .B(n1207), .CI(n1251), .CO(n786), .S(n787) );
  FA_X1 U601 ( .A(n806), .B(n793), .CI(n791), .CO(n788), .S(n789) );
  FA_X1 U602 ( .A(n795), .B(n810), .CI(n808), .CO(n790), .S(n791) );
  FA_X1 U604 ( .A(n814), .B(n816), .CI(n799), .CO(n794), .S(n795) );
  FA_X1 U606 ( .A(n1208), .B(n1318), .CI(n1230), .CO(n798), .S(n799) );
  FA_X1 U607 ( .A(n1340), .B(n1252), .CI(n803), .CO(n800), .S(n801) );
  FA_X1 U609 ( .A(n822), .B(n809), .CI(n807), .CO(n804), .S(n805) );
  FA_X1 U610 ( .A(n811), .B(n826), .CI(n824), .CO(n806), .S(n807) );
  FA_X1 U611 ( .A(n828), .B(n819), .CI(n813), .CO(n808), .S(n809) );
  FA_X1 U612 ( .A(n815), .B(n832), .CI(n817), .CO(n810), .S(n811) );
  FA_X1 U614 ( .A(n1319), .B(n1253), .CI(n1341), .CO(n814), .S(n815) );
  FA_X1 U615 ( .A(n1231), .B(n1297), .CI(n1275), .CO(n816), .S(n817) );
  FA_X1 U616 ( .A(n1363), .B(n2039), .CI(n1209), .CO(n818), .S(n819) );
  FA_X1 U618 ( .A(n827), .B(n844), .CI(n842), .CO(n822), .S(n823) );
  FA_X1 U619 ( .A(n846), .B(n848), .CI(n829), .CO(n824), .S(n825) );
  FA_X1 U620 ( .A(n835), .B(n831), .CI(n833), .CO(n826), .S(n827) );
  FA_X1 U621 ( .A(n850), .B(n854), .CI(n852), .CO(n828), .S(n829) );
  FA_X1 U622 ( .A(n1254), .B(n1320), .CI(n1298), .CO(n830), .S(n831) );
  FA_X1 U623 ( .A(n1232), .B(n1364), .CI(n1342), .CO(n832), .S(n833) );
  FA_X1 U624 ( .A(n1210), .B(n1276), .CI(n837), .CO(n834), .S(n835) );
  FA_X1 U626 ( .A(n858), .B(n843), .CI(n841), .CO(n838), .S(n839) );
  FA_X1 U627 ( .A(n845), .B(n847), .CI(n860), .CO(n840), .S(n841) );
  FA_X1 U628 ( .A(n864), .B(n849), .CI(n862), .CO(n842), .S(n843) );
  FA_X1 U629 ( .A(n855), .B(n853), .CI(n866), .CO(n844), .S(n845) );
  FA_X1 U630 ( .A(n868), .B(n870), .CI(n851), .CO(n846), .S(n847) );
  FA_X1 U631 ( .A(n1410), .B(n1365), .CI(n872), .CO(n848), .S(n849) );
  FA_X1 U632 ( .A(n1299), .B(n1277), .CI(n1343), .CO(n850), .S(n851) );
  FA_X1 U633 ( .A(n1255), .B(n1321), .CI(n874), .CO(n852), .S(n853) );
  FA_X1 U634 ( .A(n1387), .B(n1211), .CI(n1233), .CO(n854), .S(n855) );
  FA_X1 U635 ( .A(n878), .B(n861), .CI(n859), .CO(n856), .S(n857) );
  FA_X1 U636 ( .A(n863), .B(n882), .CI(n880), .CO(n858), .S(n859) );
  FA_X1 U637 ( .A(n884), .B(n867), .CI(n865), .CO(n860), .S(n861) );
  FA_X1 U638 ( .A(n888), .B(n873), .CI(n886), .CO(n862), .S(n863) );
  FA_X1 U639 ( .A(n869), .B(n890), .CI(n871), .CO(n864), .S(n865) );
  FA_X1 U640 ( .A(n894), .B(n1300), .CI(n892), .CO(n866), .S(n867) );
  FA_X1 U641 ( .A(n1234), .B(n1322), .CI(n1256), .CO(n868), .S(n869) );
  FA_X1 U642 ( .A(n1212), .B(n1366), .CI(n1344), .CO(n870), .S(n871) );
  FA_X1 U643 ( .A(n1388), .B(n1278), .CI(n875), .CO(n872), .S(n873) );
  FA_X1 U647 ( .A(n887), .B(n904), .CI(n902), .CO(n880), .S(n881) );
  FA_X1 U649 ( .A(n891), .B(n908), .CI(n895), .CO(n884), .S(n885) );
  FA_X1 U650 ( .A(n914), .B(n910), .CI(n912), .CO(n886), .S(n887) );
  FA_X1 U651 ( .A(n1367), .B(n1389), .CI(n1434), .CO(n888), .S(n889) );
  FA_X1 U652 ( .A(n1301), .B(n1257), .CI(n1345), .CO(n890), .S(n891) );
  FA_X1 U653 ( .A(n2066), .B(n1323), .CI(n1279), .CO(n892), .S(n893) );
  FA_X1 U654 ( .A(n1235), .B(n1411), .CI(n1213), .CO(n894), .S(n895) );
  FA_X1 U657 ( .A(n907), .B(n926), .CI(n905), .CO(n900), .S(n901) );
  FA_X1 U658 ( .A(n909), .B(n930), .CI(n928), .CO(n902), .S(n903) );
  FA_X1 U659 ( .A(n915), .B(n911), .CI(n913), .CO(n904), .S(n905) );
  FA_X1 U660 ( .A(n932), .B(n936), .CI(n934), .CO(n906), .S(n907) );
  FA_X1 U662 ( .A(n1280), .B(n1346), .CI(n1324), .CO(n910), .S(n911) );
  FA_X1 U664 ( .A(n1302), .B(n917), .CI(n1214), .CO(n914), .S(n915) );
  FA_X1 U666 ( .A(n942), .B(n923), .CI(n921), .CO(n918), .S(n919) );
  FA_X1 U667 ( .A(n925), .B(n927), .CI(n944), .CO(n920), .S(n921) );
  FA_X1 U668 ( .A(n929), .B(n948), .CI(n946), .CO(n922), .S(n923) );
  FA_X1 U670 ( .A(n933), .B(n952), .CI(n937), .CO(n926), .S(n927) );
  FA_X1 U672 ( .A(n939), .B(n960), .CI(n1458), .CO(n930), .S(n931) );
  FA_X1 U673 ( .A(n1325), .B(n1435), .CI(n1413), .CO(n932), .S(n933) );
  FA_X1 U674 ( .A(n1281), .B(n1369), .CI(n1391), .CO(n934), .S(n935) );
  FA_X1 U675 ( .A(n1259), .B(n1347), .CI(n1303), .CO(n936), .S(n937) );
  FA_X1 U680 ( .A(n951), .B(n970), .CI(n968), .CO(n944), .S(n945) );
  FA_X1 U681 ( .A(n972), .B(n959), .CI(n953), .CO(n946), .S(n947) );
  FA_X1 U682 ( .A(n955), .B(n974), .CI(n957), .CO(n948), .S(n949) );
  FA_X1 U683 ( .A(n976), .B(n980), .CI(n978), .CO(n950), .S(n951) );
  FA_X1 U684 ( .A(n1326), .B(n1392), .CI(n961), .CO(n952), .S(n953) );
  FA_X1 U686 ( .A(n1459), .B(n1370), .CI(n1436), .CO(n956), .S(n957) );
  FA_X1 U687 ( .A(n1260), .B(n1348), .CI(n1182), .CO(n958), .S(n959) );
  HA_X1 U688 ( .A(n1238), .B(n1216), .CO(n960), .S(n961) );
  FA_X1 U689 ( .A(n984), .B(n967), .CI(n965), .CO(n962), .S(n963) );
  FA_X1 U690 ( .A(n969), .B(n971), .CI(n986), .CO(n964), .S(n965) );
  FA_X1 U691 ( .A(n973), .B(n990), .CI(n988), .CO(n966), .S(n967) );
  FA_X1 U697 ( .A(n1283), .B(n1460), .CI(n1371), .CO(n978), .S(n979) );
  FA_X1 U698 ( .A(n1239), .B(n1349), .CI(n1261), .CO(n980), .S(n981) );
  FA_X1 U699 ( .A(n1004), .B(n987), .CI(n985), .CO(n982), .S(n983) );
  FA_X1 U700 ( .A(n989), .B(n991), .CI(n1006), .CO(n984), .S(n985) );
  FA_X1 U701 ( .A(n993), .B(n1010), .CI(n1008), .CO(n986), .S(n987) );
  FA_X1 U702 ( .A(n999), .B(n997), .CI(n1012), .CO(n988), .S(n989) );
  FA_X1 U703 ( .A(n1014), .B(n1016), .CI(n995), .CO(n990), .S(n991) );
  FA_X1 U706 ( .A(n1284), .B(n1438), .CI(n1372), .CO(n996), .S(n997) );
  FA_X1 U707 ( .A(n1461), .B(n1350), .CI(n1183), .CO(n998), .S(n999) );
  HA_X1 U708 ( .A(n1240), .B(n1262), .CO(n1000), .S(n1001) );
  FA_X1 U709 ( .A(n1022), .B(n1007), .CI(n1005), .CO(n1002), .S(n1003) );
  FA_X1 U710 ( .A(n1009), .B(n1011), .CI(n1024), .CO(n1004), .S(n1005) );
  FA_X1 U711 ( .A(n1013), .B(n1028), .CI(n1026), .CO(n1006), .S(n1007) );
  FA_X1 U712 ( .A(n1019), .B(n1015), .CI(n1017), .CO(n1008), .S(n1009) );
  FA_X1 U713 ( .A(n1030), .B(n1034), .CI(n1241), .CO(n1010), .S(n1011) );
  FA_X1 U714 ( .A(n1036), .B(n1439), .CI(n1032), .CO(n1012), .S(n1013) );
  FA_X1 U715 ( .A(n1462), .B(n1395), .CI(n1417), .CO(n1014), .S(n1015) );
  FA_X1 U716 ( .A(n1307), .B(n1373), .CI(n1329), .CO(n1016), .S(n1017) );
  FA_X1 U718 ( .A(n1040), .B(n1025), .CI(n1023), .CO(n1020), .S(n1021) );
  FA_X1 U719 ( .A(n1027), .B(n1044), .CI(n1042), .CO(n1022), .S(n1023) );
  FA_X1 U720 ( .A(n1046), .B(n1035), .CI(n1029), .CO(n1024), .S(n1025) );
  FA_X1 U721 ( .A(n1033), .B(n1048), .CI(n1031), .CO(n1026), .S(n1027) );
  FA_X1 U722 ( .A(n1052), .B(n1050), .CI(n1037), .CO(n1028), .S(n1029) );
  FA_X1 U723 ( .A(n1418), .B(n1440), .CI(n1352), .CO(n1030), .S(n1031) );
  FA_X1 U724 ( .A(n1463), .B(n1330), .CI(n1396), .CO(n1032), .S(n1033) );
  FA_X1 U725 ( .A(n1308), .B(n1374), .CI(n1184), .CO(n1034), .S(n1035) );
  HA_X1 U726 ( .A(n1264), .B(n1286), .CO(n1036), .S(n1037) );
  FA_X1 U727 ( .A(n1056), .B(n1043), .CI(n1041), .CO(n1038), .S(n1039) );
  FA_X1 U728 ( .A(n1058), .B(n1047), .CI(n1045), .CO(n1040), .S(n1041) );
  FA_X1 U730 ( .A(n1049), .B(n1265), .CI(n1051), .CO(n1044), .S(n1045) );
  FA_X1 U731 ( .A(n1064), .B(n1068), .CI(n1066), .CO(n1046), .S(n1047) );
  FA_X1 U732 ( .A(n1397), .B(n1441), .CI(n1419), .CO(n1048), .S(n1049) );
  FA_X1 U733 ( .A(n1331), .B(n1353), .CI(n1375), .CO(n1050), .S(n1051) );
  FA_X1 U734 ( .A(n1287), .B(n1309), .CI(n1464), .CO(n1052), .S(n1053) );
  FA_X1 U735 ( .A(n1072), .B(n1059), .CI(n1057), .CO(n1054), .S(n1055) );
  FA_X1 U736 ( .A(n1074), .B(n1063), .CI(n1061), .CO(n1056), .S(n1057) );
  FA_X1 U737 ( .A(n1067), .B(n1065), .CI(n1076), .CO(n1058), .S(n1059) );
  FA_X1 U739 ( .A(n1398), .B(n1420), .CI(n1069), .CO(n1062), .S(n1063) );
  FA_X1 U740 ( .A(n1442), .B(n1354), .CI(n1332), .CO(n1064), .S(n1065) );
  FA_X1 U741 ( .A(n1465), .B(n1376), .CI(n1185), .CO(n1066), .S(n1067) );
  HA_X1 U742 ( .A(n1288), .B(n1310), .CO(n1068), .S(n1069) );
  FA_X1 U743 ( .A(n1086), .B(n1075), .CI(n1073), .CO(n1070), .S(n1071) );
  FA_X1 U744 ( .A(n1088), .B(n1090), .CI(n1077), .CO(n1072), .S(n1073) );
  FA_X1 U748 ( .A(n1355), .B(n1443), .CI(n1377), .CO(n1080), .S(n1081) );
  FA_X1 U749 ( .A(n1311), .B(n1333), .CI(n1466), .CO(n1082), .S(n1083) );
  FA_X1 U750 ( .A(n1100), .B(n1089), .CI(n1087), .CO(n1084), .S(n1085) );
  FA_X1 U751 ( .A(n1102), .B(n1104), .CI(n1091), .CO(n1086), .S(n1087) );
  FA_X1 U752 ( .A(n1093), .B(n1106), .CI(n1095), .CO(n1088), .S(n1089) );
  FA_X1 U753 ( .A(n1097), .B(n1422), .CI(n1108), .CO(n1090), .S(n1091) );
  FA_X1 U754 ( .A(n1378), .B(n1444), .CI(n1356), .CO(n1092), .S(n1093) );
  HA_X1 U756 ( .A(n1312), .B(n1334), .CO(n1096), .S(n1097) );
  FA_X1 U757 ( .A(n1103), .B(n1112), .CI(n1101), .CO(n1098), .S(n1099) );
  FA_X1 U758 ( .A(n1114), .B(n1109), .CI(n1105), .CO(n1100), .S(n1101) );
  FA_X1 U759 ( .A(n1313), .B(n1116), .CI(n1107), .CO(n1102), .S(n1103) );
  FA_X1 U760 ( .A(n1120), .B(n1423), .CI(n1118), .CO(n1104), .S(n1105) );
  FA_X1 U761 ( .A(n1379), .B(n1445), .CI(n1401), .CO(n1106), .S(n1107) );
  FA_X1 U762 ( .A(n1335), .B(n1468), .CI(n1357), .CO(n1108), .S(n1109) );
  FA_X1 U763 ( .A(n1124), .B(n1115), .CI(n1113), .CO(n1110), .S(n1111) );
  FA_X1 U764 ( .A(n1119), .B(n1117), .CI(n1126), .CO(n1112), .S(n1113) );
  FA_X1 U765 ( .A(n1130), .B(n1121), .CI(n1128), .CO(n1114), .S(n1115) );
  FA_X1 U766 ( .A(n1380), .B(n1446), .CI(n1424), .CO(n1116), .S(n1117) );
  FA_X1 U767 ( .A(n1469), .B(n1402), .CI(n1187), .CO(n1118), .S(n1119) );
  HA_X1 U768 ( .A(n1336), .B(n1358), .CO(n1120), .S(n1121) );
  FA_X1 U769 ( .A(n1127), .B(n1134), .CI(n1125), .CO(n1122), .S(n1123) );
  FA_X1 U770 ( .A(n1131), .B(n1129), .CI(n1136), .CO(n1124), .S(n1125) );
  FA_X1 U771 ( .A(n1337), .B(n1140), .CI(n1138), .CO(n1126), .S(n1127) );
  FA_X1 U772 ( .A(n1403), .B(n1447), .CI(n1425), .CO(n1128), .S(n1129) );
  FA_X1 U773 ( .A(n1359), .B(n1470), .CI(n1381), .CO(n1130), .S(n1131) );
  FA_X1 U774 ( .A(n1144), .B(n1137), .CI(n1135), .CO(n1132), .S(n1133) );
  FA_X1 U775 ( .A(n1146), .B(n1148), .CI(n1139), .CO(n1134), .S(n1135) );
  FA_X1 U776 ( .A(n1404), .B(n1448), .CI(n1141), .CO(n1136), .S(n1137) );
  FA_X1 U777 ( .A(n1188), .B(n1426), .CI(n1471), .CO(n1138), .S(n1139) );
  HA_X1 U778 ( .A(n1360), .B(n1382), .CO(n1140), .S(n1141) );
  FA_X1 U779 ( .A(n1152), .B(n1147), .CI(n1145), .CO(n1142), .S(n1143) );
  FA_X1 U780 ( .A(n1361), .B(n1154), .CI(n1149), .CO(n1144), .S(n1145) );
  FA_X1 U781 ( .A(n1427), .B(n1449), .CI(n1156), .CO(n1146), .S(n1147) );
  FA_X1 U782 ( .A(n1383), .B(n1472), .CI(n1405), .CO(n1148), .S(n1149) );
  FA_X1 U783 ( .A(n1160), .B(n1155), .CI(n1153), .CO(n1150), .S(n1151) );
  FA_X1 U784 ( .A(n1157), .B(n1473), .CI(n1162), .CO(n1152), .S(n1153) );
  FA_X1 U785 ( .A(n1450), .B(n1428), .CI(n1189), .CO(n1154), .S(n1155) );
  HA_X1 U786 ( .A(n1384), .B(n1406), .CO(n1156), .S(n1157) );
  FA_X1 U787 ( .A(n1163), .B(n1385), .CI(n1164), .CO(n1158), .S(n1159) );
  FA_X1 U788 ( .A(n1168), .B(n1429), .CI(n1166), .CO(n1160), .S(n1161) );
  FA_X1 U789 ( .A(n1451), .B(n1474), .CI(n1407), .CO(n1162), .S(n1163) );
  FA_X1 U790 ( .A(n1172), .B(n1169), .CI(n1167), .CO(n1164), .S(n1165) );
  FA_X1 U791 ( .A(n1452), .B(n1475), .CI(n1190), .CO(n1166), .S(n1167) );
  HA_X1 U792 ( .A(n1408), .B(n1430), .CO(n1168), .S(n1169) );
  FA_X1 U793 ( .A(n1409), .B(n1176), .CI(n1173), .CO(n1170), .S(n1171) );
  FA_X1 U794 ( .A(n1476), .B(n1453), .CI(n1431), .CO(n1172), .S(n1173) );
  FA_X1 U795 ( .A(n1191), .B(n1454), .CI(n1177), .CO(n1174), .S(n1175) );
  HA_X1 U796 ( .A(n1432), .B(n1477), .CO(n1176), .S(n1177) );
  FA_X1 U797 ( .A(n1455), .B(n1478), .CI(n1180), .CO(n1178), .S(n1179) );
  HA_X1 U798 ( .A(n1456), .B(n1479), .CO(n1180), .S(n1181) );
  XNOR2_X1 U1448 ( .A(n551), .B(n1929), .ZN(product[23]) );
  AND2_X1 U1449 ( .A1(n674), .A2(n550), .ZN(n1929) );
  XNOR2_X1 U1450 ( .A(a[18]), .B(a[19]), .ZN(n2156) );
  INV_X1 U1451 ( .A(a[13]), .ZN(n1930) );
  OR2_X2 U1452 ( .A1(n2026), .A2(n2018), .ZN(n1931) );
  INV_X1 U1453 ( .A(n2162), .ZN(n1932) );
  AND2_X1 U1454 ( .A1(n2273), .A2(n2272), .ZN(n1933) );
  OR2_X2 U1455 ( .A1(n2257), .A2(n2159), .ZN(n1998) );
  INV_X1 U1456 ( .A(n2257), .ZN(n2286) );
  INV_X1 U1457 ( .A(n2257), .ZN(n2285) );
  INV_X1 U1458 ( .A(n2162), .ZN(n2280) );
  XNOR2_X1 U1459 ( .A(n1080), .B(n1934), .ZN(n1061) );
  XNOR2_X1 U1460 ( .A(n2058), .B(n1082), .ZN(n1934) );
  INV_X1 U1461 ( .A(n2042), .ZN(n1935) );
  BUF_X2 U1462 ( .A(n2277), .Z(n2175) );
  XOR2_X2 U1463 ( .A(a[20]), .B(a[19]), .Z(n2257) );
  CLKBUF_X3 U1464 ( .A(n293), .Z(n1936) );
  NOR2_X1 U1465 ( .A1(n542), .A2(n547), .ZN(n1937) );
  NOR2_X2 U1466 ( .A1(n941), .A2(n962), .ZN(n547) );
  AND2_X2 U1467 ( .A1(n775), .A2(n788), .ZN(n1938) );
  INV_X4 U1468 ( .A(n1938), .ZN(n474) );
  OR2_X2 U1469 ( .A1(n2155), .A2(n2019), .ZN(n1939) );
  CLKBUF_X2 U1470 ( .A(n2070), .Z(n1941) );
  BUF_X2 U1471 ( .A(n2070), .Z(n1940) );
  CLKBUF_X1 U1472 ( .A(n2070), .Z(n2205) );
  XNOR2_X1 U1473 ( .A(a[0]), .B(n2362), .ZN(n1817) );
  BUF_X1 U1474 ( .A(n514), .Z(n1942) );
  BUF_X1 U1475 ( .A(n2265), .Z(n2054) );
  CLKBUF_X3 U1476 ( .A(n2055), .Z(n2179) );
  BUF_X1 U1477 ( .A(n2089), .Z(n1943) );
  XOR2_X1 U1478 ( .A(n924), .B(n903), .Z(n1944) );
  XOR2_X1 U1479 ( .A(n922), .B(n1944), .Z(n899) );
  NAND2_X1 U1480 ( .A1(n922), .A2(n924), .ZN(n1945) );
  NAND2_X1 U1481 ( .A1(n922), .A2(n903), .ZN(n1946) );
  NAND2_X1 U1482 ( .A1(n924), .A2(n903), .ZN(n1947) );
  NAND3_X1 U1483 ( .A1(n1945), .A2(n1946), .A3(n1947), .ZN(n898) );
  OR2_X1 U1484 ( .A1(n2159), .A2(n2257), .ZN(n2089) );
  CLKBUF_X1 U1485 ( .A(n1001), .Z(n2106) );
  CLKBUF_X1 U1486 ( .A(n2306), .Z(n1948) );
  BUF_X4 U1487 ( .A(n2306), .Z(n1949) );
  INV_X1 U1488 ( .A(n2307), .ZN(n2306) );
  XOR2_X1 U1489 ( .A(n840), .B(n825), .Z(n1950) );
  XOR2_X1 U1490 ( .A(n823), .B(n1950), .Z(n821) );
  NAND2_X1 U1491 ( .A1(n823), .A2(n840), .ZN(n1951) );
  NAND2_X1 U1492 ( .A1(n823), .A2(n825), .ZN(n1952) );
  NAND2_X1 U1493 ( .A1(n840), .A2(n825), .ZN(n1953) );
  NAND3_X1 U1494 ( .A1(n1951), .A2(n1952), .A3(n1953), .ZN(n820) );
  BUF_X1 U1495 ( .A(n1502), .Z(n1954) );
  NOR2_X1 U1496 ( .A1(n520), .A2(n513), .ZN(n1955) );
  XNOR2_X1 U1497 ( .A(a[22]), .B(n2313), .ZN(n1956) );
  NAND3_X1 U1498 ( .A1(n2099), .A2(n2100), .A3(n2101), .ZN(n1957) );
  INV_X1 U1499 ( .A(n2285), .ZN(n1958) );
  XOR2_X1 U1500 ( .A(n920), .B(n901), .Z(n1959) );
  XOR2_X1 U1501 ( .A(n899), .B(n1959), .Z(n897) );
  NAND2_X1 U1502 ( .A1(n899), .A2(n920), .ZN(n1960) );
  NAND2_X1 U1503 ( .A1(n899), .A2(n901), .ZN(n1961) );
  NAND2_X1 U1504 ( .A1(n920), .A2(n901), .ZN(n1962) );
  NAND3_X1 U1505 ( .A1(n1960), .A2(n1961), .A3(n1962), .ZN(n896) );
  CLKBUF_X1 U1506 ( .A(n506), .Z(n2042) );
  CLKBUF_X1 U1507 ( .A(n490), .Z(n2109) );
  CLKBUF_X3 U1508 ( .A(n2351), .Z(n2008) );
  INV_X1 U1509 ( .A(n2033), .ZN(n2164) );
  INV_X1 U1510 ( .A(n2072), .ZN(n2231) );
  INV_X1 U1511 ( .A(n2070), .ZN(n2166) );
  AND2_X1 U1512 ( .A1(n1193), .A2(n1481), .ZN(n1963) );
  OR2_X1 U1513 ( .A1(n1457), .A2(n1480), .ZN(n1964) );
  OR2_X1 U1514 ( .A1(n1179), .A2(n1433), .ZN(n1965) );
  AND2_X1 U1515 ( .A1(n1039), .A2(n1054), .ZN(n1966) );
  AND2_X1 U1516 ( .A1(n1123), .A2(n1132), .ZN(n1967) );
  AND2_X1 U1517 ( .A1(n1143), .A2(n1150), .ZN(n1968) );
  AND2_X1 U1518 ( .A1(n1151), .A2(n1158), .ZN(n1969) );
  OR2_X1 U1519 ( .A1(n2160), .A2(n2208), .ZN(n1970) );
  AND2_X1 U1520 ( .A1(n1457), .A2(n1480), .ZN(n1971) );
  AND2_X1 U1521 ( .A1(n1179), .A2(n1433), .ZN(n1972) );
  AND2_X1 U1522 ( .A1(n1111), .A2(n1122), .ZN(n1973) );
  AND2_X1 U1523 ( .A1(n1133), .A2(n1142), .ZN(n1974) );
  AND2_X1 U1524 ( .A1(n1055), .A2(n1070), .ZN(n1975) );
  AND2_X1 U1525 ( .A1(n1021), .A2(n1038), .ZN(n1976) );
  OR2_X1 U1526 ( .A1(n1151), .A2(n1158), .ZN(n1977) );
  OR2_X1 U1527 ( .A1(n1123), .A2(n1132), .ZN(n1978) );
  OR2_X1 U1528 ( .A1(n1039), .A2(n1054), .ZN(n1979) );
  OR2_X1 U1529 ( .A1(n1143), .A2(n1150), .ZN(n1980) );
  XNOR2_X1 U1530 ( .A(n560), .B(n1981), .ZN(product[22]) );
  AND2_X1 U1531 ( .A1(n2088), .A2(n559), .ZN(n1981) );
  XNOR2_X1 U1532 ( .A(n2054), .B(n1982), .ZN(product[34]) );
  AND2_X1 U1533 ( .A1(n663), .A2(n439), .ZN(n1982) );
  NOR2_X1 U1534 ( .A1(n1003), .A2(n1020), .ZN(n1983) );
  OR2_X2 U1535 ( .A1(n2148), .A2(n2149), .ZN(n1351) );
  BUF_X1 U1536 ( .A(n536), .Z(n1989) );
  BUF_X1 U1537 ( .A(n536), .Z(n1987) );
  CLKBUF_X1 U1538 ( .A(n251), .Z(n2303) );
  BUF_X4 U1539 ( .A(n251), .Z(n2304) );
  OR2_X2 U1540 ( .A1(n2169), .A2(n2194), .ZN(n1984) );
  BUF_X1 U1541 ( .A(n2294), .Z(n1986) );
  BUF_X2 U1542 ( .A(n2294), .Z(n1985) );
  BUF_X1 U1543 ( .A(n536), .Z(n1988) );
  INV_X1 U1544 ( .A(n508), .ZN(n1990) );
  CLKBUF_X1 U1545 ( .A(n521), .Z(n1991) );
  AND2_X2 U1546 ( .A1(n1817), .A2(n2303), .ZN(n2172) );
  CLKBUF_X1 U1547 ( .A(n520), .Z(n1992) );
  XNOR2_X1 U1548 ( .A(a[6]), .B(n2355), .ZN(n1993) );
  XNOR2_X1 U1549 ( .A(a[6]), .B(n2355), .ZN(n2194) );
  OR2_X1 U1550 ( .A1(n839), .A2(n856), .ZN(n1994) );
  BUF_X1 U1551 ( .A(n2237), .Z(n1995) );
  CLKBUF_X1 U1552 ( .A(n897), .Z(n1996) );
  BUF_X1 U1553 ( .A(n1528), .Z(n1997) );
  BUF_X2 U1554 ( .A(n2277), .Z(n2176) );
  INV_X1 U1555 ( .A(n2091), .ZN(n1999) );
  CLKBUF_X1 U1556 ( .A(n2283), .Z(n2000) );
  CLKBUF_X1 U1557 ( .A(n2305), .Z(n2002) );
  CLKBUF_X3 U1558 ( .A(n2305), .Z(n2001) );
  INV_X1 U1559 ( .A(n2307), .ZN(n2305) );
  NOR2_X1 U1560 ( .A1(n877), .A2(n896), .ZN(n2003) );
  NOR2_X1 U1561 ( .A1(n877), .A2(n896), .ZN(n531) );
  INV_X1 U1562 ( .A(n1970), .ZN(n2004) );
  CLKBUF_X1 U1563 ( .A(n2334), .Z(n2005) );
  CLKBUF_X1 U1564 ( .A(n552), .Z(n2006) );
  OR2_X2 U1565 ( .A1(n1215), .A2(n1237), .ZN(n938) );
  CLKBUF_X1 U1566 ( .A(n2351), .Z(n2007) );
  XNOR2_X1 U1567 ( .A(n1000), .B(n2152), .ZN(n2009) );
  OR2_X2 U1568 ( .A1(n2171), .A2(n2198), .ZN(n2010) );
  XNOR2_X2 U1569 ( .A(n2338), .B(a[12]), .ZN(n2198) );
  NOR2_X1 U1570 ( .A1(n558), .A2(n563), .ZN(n552) );
  INV_X1 U1571 ( .A(a[15]), .ZN(n2012) );
  INV_X1 U1572 ( .A(a[15]), .ZN(n2011) );
  CLKBUF_X1 U1573 ( .A(n2286), .Z(n2013) );
  CLKBUF_X1 U1574 ( .A(n2293), .Z(n2014) );
  BUF_X1 U1575 ( .A(n2293), .Z(n2016) );
  BUF_X2 U1576 ( .A(n2293), .Z(n2015) );
  XOR2_X1 U1577 ( .A(a[18]), .B(a[17]), .Z(n2017) );
  XNOR2_X1 U1578 ( .A(a[14]), .B(n2332), .ZN(n2019) );
  XNOR2_X1 U1579 ( .A(a[14]), .B(n1930), .ZN(n2018) );
  XNOR2_X1 U1580 ( .A(a[14]), .B(n1930), .ZN(n2153) );
  INV_X1 U1581 ( .A(n2011), .ZN(n2021) );
  INV_X1 U1582 ( .A(n2012), .ZN(n2020) );
  BUF_X1 U1583 ( .A(n1258), .Z(n2022) );
  INV_X1 U1584 ( .A(n2300), .ZN(n2023) );
  CLKBUF_X1 U1585 ( .A(n2292), .Z(n2024) );
  XNOR2_X1 U1586 ( .A(n950), .B(n2025), .ZN(n925) );
  XNOR2_X1 U1587 ( .A(n935), .B(n931), .ZN(n2025) );
  XOR2_X1 U1588 ( .A(a[14]), .B(n2325), .Z(n2026) );
  INV_X1 U1589 ( .A(n1939), .ZN(n2027) );
  INV_X1 U1590 ( .A(n2363), .ZN(n2029) );
  INV_X1 U1591 ( .A(n2363), .ZN(n2028) );
  OR2_X1 U1592 ( .A1(n2160), .A2(n2208), .ZN(n2030) );
  INV_X1 U1593 ( .A(n2162), .ZN(n2031) );
  NOR2_X2 U1594 ( .A1(n2163), .A2(n2157), .ZN(n2162) );
  BUF_X2 U1595 ( .A(n293), .Z(n2199) );
  INV_X1 U1596 ( .A(n2173), .ZN(n2032) );
  OR2_X2 U1597 ( .A1(n2158), .A2(n2165), .ZN(n2033) );
  OR2_X1 U1598 ( .A1(n2165), .A2(n2158), .ZN(n2055) );
  INV_X1 U1599 ( .A(n1984), .ZN(n2034) );
  CLKBUF_X1 U1600 ( .A(n2298), .Z(n2035) );
  BUF_X2 U1601 ( .A(n2298), .Z(n2036) );
  CLKBUF_X1 U1602 ( .A(n2313), .Z(n2037) );
  INV_X1 U1603 ( .A(n2061), .ZN(n2038) );
  BUF_X1 U1604 ( .A(n2030), .Z(n2046) );
  BUF_X2 U1605 ( .A(n2030), .Z(n2048) );
  INV_X2 U1606 ( .A(n2363), .ZN(n2360) );
  OAI22_X1 U1607 ( .A1(n1984), .A2(n1683), .B1(n1682), .B2(n2035), .ZN(n2039)
         );
  INV_X1 U1608 ( .A(n2172), .ZN(n2041) );
  INV_X1 U1609 ( .A(n2172), .ZN(n2040) );
  INV_X1 U1610 ( .A(n2172), .ZN(n2282) );
  INV_X1 U1611 ( .A(n2289), .ZN(n2043) );
  INV_X2 U1612 ( .A(n1995), .ZN(n2289) );
  XOR2_X1 U1613 ( .A(a[16]), .B(a[15]), .Z(n2237) );
  INV_X1 U1614 ( .A(n2331), .ZN(n2045) );
  INV_X1 U1615 ( .A(n2331), .ZN(n2044) );
  BUF_X2 U1616 ( .A(n2030), .Z(n2047) );
  BUF_X2 U1617 ( .A(n2055), .Z(n2180) );
  INV_X1 U1618 ( .A(n2295), .ZN(n2049) );
  OAI22_X1 U1619 ( .A1(n2040), .A2(n1766), .B1(n1765), .B2(n2304), .ZN(n2050)
         );
  AND2_X1 U1620 ( .A1(n2273), .A2(n2272), .ZN(n2051) );
  CLKBUF_X3 U1621 ( .A(a[17]), .Z(n2052) );
  INV_X2 U1622 ( .A(n2320), .ZN(n2317) );
  XNOR2_X1 U1623 ( .A(n1351), .B(n2053), .ZN(n1019) );
  XNOR2_X1 U1624 ( .A(n1263), .B(n1285), .ZN(n2053) );
  XOR2_X1 U1625 ( .A(a[10]), .B(a[9]), .Z(n2158) );
  INV_X2 U1626 ( .A(n2153), .ZN(n2291) );
  INV_X2 U1627 ( .A(n2019), .ZN(n2290) );
  INV_X2 U1628 ( .A(n2244), .ZN(n2284) );
  CLKBUF_X1 U1629 ( .A(n535), .Z(n2056) );
  XNOR2_X2 U1630 ( .A(a[16]), .B(a[15]), .ZN(n2057) );
  CLKBUF_X1 U1631 ( .A(n2087), .Z(n2068) );
  NAND3_X1 U1632 ( .A1(n2250), .A2(n2251), .A3(n2252), .ZN(n2058) );
  OR2_X2 U1633 ( .A1(n2171), .A2(n2198), .ZN(n2059) );
  OR2_X1 U1634 ( .A1(n2171), .A2(n2198), .ZN(n2081) );
  NOR2_X2 U1635 ( .A1(n727), .A2(n736), .ZN(n428) );
  AOI21_X2 U1636 ( .B1(n426), .B2(n445), .A(n427), .ZN(n421) );
  INV_X1 U1637 ( .A(n2059), .ZN(n2170) );
  INV_X2 U1638 ( .A(n2342), .ZN(n2339) );
  INV_X1 U1639 ( .A(n2090), .ZN(n2060) );
  NOR2_X1 U1640 ( .A1(n2174), .A2(n2237), .ZN(n2061) );
  INV_X2 U1641 ( .A(n2172), .ZN(n2281) );
  XNOR2_X1 U1642 ( .A(n2062), .B(n2106), .ZN(n993) );
  XNOR2_X1 U1643 ( .A(n1018), .B(n1394), .ZN(n2062) );
  XNOR2_X1 U1644 ( .A(n2063), .B(n943), .ZN(n941) );
  XNOR2_X1 U1645 ( .A(n964), .B(n945), .ZN(n2063) );
  INV_X2 U1646 ( .A(n2355), .ZN(n2352) );
  INV_X2 U1647 ( .A(n2312), .ZN(n2310) );
  CLKBUF_X1 U1648 ( .A(n505), .Z(n2064) );
  OR2_X1 U1649 ( .A1(n502), .A2(n495), .ZN(n2065) );
  INV_X1 U1650 ( .A(n917), .ZN(n2066) );
  OAI22_X1 U1651 ( .A1(n1970), .A2(n1733), .B1(n1732), .B2(n2302), .ZN(n916)
         );
  CLKBUF_X1 U1652 ( .A(n956), .Z(n2067) );
  CLKBUF_X1 U1653 ( .A(n977), .Z(n2069) );
  OR2_X2 U1654 ( .A1(n2167), .A2(n2080), .ZN(n2070) );
  XOR2_X1 U1655 ( .A(n2313), .B(a[20]), .Z(n2159) );
  XOR2_X1 U1656 ( .A(a[6]), .B(n2349), .Z(n2169) );
  INV_X1 U1657 ( .A(n2348), .ZN(n2345) );
  BUF_X1 U1658 ( .A(n2203), .Z(n2071) );
  XNOR2_X1 U1659 ( .A(a[8]), .B(a[7]), .ZN(n2072) );
  INV_X2 U1660 ( .A(n2231), .ZN(n2296) );
  NAND3_X1 U1661 ( .A1(n2211), .A2(n2212), .A3(n2213), .ZN(n2073) );
  NAND2_X1 U1662 ( .A1(n1080), .A2(n1078), .ZN(n2074) );
  NAND2_X1 U1663 ( .A1(n1080), .A2(n1082), .ZN(n2075) );
  NAND2_X1 U1664 ( .A1(n1078), .A2(n1082), .ZN(n2076) );
  NAND3_X1 U1665 ( .A1(n2074), .A2(n2075), .A3(n2076), .ZN(n1060) );
  XOR2_X1 U1666 ( .A(a[2]), .B(a[1]), .Z(n2077) );
  OR2_X1 U1667 ( .A1(n1970), .A2(n1742), .ZN(n2078) );
  OR2_X1 U1668 ( .A1(n2301), .A2(n1741), .ZN(n2079) );
  NAND2_X1 U1669 ( .A1(n2078), .A2(n2079), .ZN(n1443) );
  XOR2_X1 U1670 ( .A(a[2]), .B(a[1]), .Z(n2208) );
  INV_X2 U1671 ( .A(n2077), .ZN(n2301) );
  XNOR2_X1 U1672 ( .A(a[22]), .B(n2313), .ZN(n2080) );
  BUF_X2 U1673 ( .A(n2070), .Z(n2204) );
  XOR2_X1 U1674 ( .A(a[4]), .B(a[3]), .Z(n2157) );
  XOR2_X1 U1675 ( .A(n1274), .B(n1296), .Z(n2082) );
  XOR2_X1 U1676 ( .A(n818), .B(n2082), .Z(n797) );
  NAND2_X1 U1677 ( .A1(n818), .A2(n1274), .ZN(n2083) );
  NAND2_X1 U1678 ( .A1(n818), .A2(n1296), .ZN(n2084) );
  NAND2_X1 U1679 ( .A1(n1274), .A2(n1296), .ZN(n2085) );
  NAND3_X1 U1680 ( .A1(n2083), .A2(n2084), .A3(n2085), .ZN(n796) );
  OAI21_X1 U1681 ( .B1(n2003), .B2(n535), .A(n532), .ZN(n2086) );
  INV_X1 U1682 ( .A(n2359), .ZN(n2356) );
  INV_X2 U1683 ( .A(n2359), .ZN(n2357) );
  BUF_X2 U1684 ( .A(n2031), .Z(n2177) );
  NOR2_X1 U1685 ( .A1(n919), .A2(n940), .ZN(n2087) );
  NOR2_X1 U1686 ( .A1(n940), .A2(n919), .ZN(n542) );
  OR2_X1 U1687 ( .A1(n963), .A2(n982), .ZN(n2088) );
  INV_X2 U1688 ( .A(n2168), .ZN(n2108) );
  OR2_X1 U1689 ( .A1(n534), .A2(n2003), .ZN(n2090) );
  OR2_X1 U1690 ( .A1(n918), .A2(n1996), .ZN(n2091) );
  NOR2_X1 U1691 ( .A1(n2089), .A2(n1528), .ZN(n2092) );
  NOR2_X1 U1692 ( .A1(n1527), .A2(n2286), .ZN(n2093) );
  OR2_X1 U1693 ( .A1(n2092), .A2(n2093), .ZN(n1238) );
  NOR2_X1 U1694 ( .A1(n963), .A2(n982), .ZN(n558) );
  INV_X1 U1695 ( .A(n293), .ZN(n2094) );
  INV_X1 U1696 ( .A(n2316), .ZN(n2096) );
  INV_X1 U1697 ( .A(n2316), .ZN(n2095) );
  OR2_X2 U1698 ( .A1(n2156), .A2(n2154), .ZN(n293) );
  NOR2_X1 U1699 ( .A1(n805), .A2(n820), .ZN(n2097) );
  NOR2_X1 U1700 ( .A1(n805), .A2(n820), .ZN(n495) );
  INV_X1 U1701 ( .A(n555), .ZN(n2098) );
  NAND2_X1 U1702 ( .A1(n1018), .A2(n1394), .ZN(n2099) );
  NAND2_X1 U1703 ( .A1(n1018), .A2(n1001), .ZN(n2100) );
  NAND2_X1 U1704 ( .A1(n1001), .A2(n1394), .ZN(n2101) );
  NAND3_X1 U1705 ( .A1(n2101), .A2(n2100), .A3(n2099), .ZN(n992) );
  XOR2_X1 U1706 ( .A(n975), .B(n981), .Z(n2102) );
  XOR2_X1 U1707 ( .A(n2102), .B(n992), .Z(n969) );
  NAND2_X1 U1708 ( .A1(n2009), .A2(n981), .ZN(n2103) );
  NAND2_X1 U1709 ( .A1(n2009), .A2(n1957), .ZN(n2104) );
  NAND2_X1 U1710 ( .A1(n981), .A2(n992), .ZN(n2105) );
  NAND3_X1 U1711 ( .A1(n2103), .A2(n2104), .A3(n2105), .ZN(n968) );
  INV_X1 U1712 ( .A(n2208), .ZN(n2302) );
  AOI21_X1 U1713 ( .B1(n581), .B2(n567), .A(n568), .ZN(n2107) );
  INV_X1 U1714 ( .A(n2168), .ZN(n2278) );
  INV_X2 U1715 ( .A(n2337), .ZN(n2334) );
  NOR2_X1 U1716 ( .A1(n2174), .A2(n2237), .ZN(n2173) );
  INV_X1 U1717 ( .A(n1998), .ZN(n2110) );
  XOR2_X1 U1718 ( .A(n1412), .B(n1236), .Z(n2111) );
  XOR2_X1 U1719 ( .A(n2111), .B(n2022), .Z(n913) );
  NAND2_X1 U1720 ( .A1(n1258), .A2(n1412), .ZN(n2112) );
  NAND2_X1 U1721 ( .A1(n1258), .A2(n1236), .ZN(n2113) );
  NAND2_X1 U1722 ( .A1(n1412), .A2(n1236), .ZN(n2114) );
  NAND3_X1 U1723 ( .A1(n2113), .A2(n2112), .A3(n2114), .ZN(n912) );
  INV_X1 U1724 ( .A(n2065), .ZN(n2115) );
  NOR2_X1 U1725 ( .A1(n495), .A2(n502), .ZN(n489) );
  NOR2_X1 U1726 ( .A1(n2169), .A2(n1993), .ZN(n2168) );
  XOR2_X1 U1727 ( .A(n947), .B(n949), .Z(n2116) );
  XOR2_X1 U1728 ( .A(n2116), .B(n966), .Z(n943) );
  NAND2_X1 U1729 ( .A1(n947), .A2(n949), .ZN(n2117) );
  NAND2_X1 U1730 ( .A1(n947), .A2(n966), .ZN(n2118) );
  NAND2_X1 U1731 ( .A1(n949), .A2(n966), .ZN(n2119) );
  NAND3_X1 U1732 ( .A1(n2117), .A2(n2118), .A3(n2119), .ZN(n942) );
  NAND2_X1 U1733 ( .A1(n964), .A2(n945), .ZN(n2120) );
  NAND2_X1 U1734 ( .A1(n964), .A2(n943), .ZN(n2121) );
  NAND2_X1 U1735 ( .A1(n945), .A2(n943), .ZN(n2122) );
  NAND3_X1 U1736 ( .A1(n2120), .A2(n2121), .A3(n2122), .ZN(n940) );
  XOR2_X1 U1737 ( .A(a[14]), .B(n2011), .Z(n2155) );
  INV_X2 U1738 ( .A(n2326), .ZN(n2322) );
  AOI21_X1 U1739 ( .B1(n1955), .B2(n526), .A(n512), .ZN(n506) );
  INV_X2 U1740 ( .A(n2312), .ZN(n2309) );
  XOR2_X1 U1741 ( .A(n801), .B(n797), .Z(n2214) );
  XOR2_X1 U1742 ( .A(n2123), .B(n1094), .Z(n1077) );
  XOR2_X1 U1743 ( .A(n1092), .B(n1289), .Z(n2123) );
  XOR2_X1 U1744 ( .A(n1306), .B(n2245), .Z(n995) );
  XNOR2_X1 U1745 ( .A(n2067), .B(n2124), .ZN(n929) );
  XNOR2_X1 U1746 ( .A(n958), .B(n954), .ZN(n2124) );
  AND2_X1 U1747 ( .A1(n2125), .A2(n2072), .ZN(n2161) );
  XOR2_X1 U1748 ( .A(a[8]), .B(a[9]), .Z(n2125) );
  INV_X1 U1749 ( .A(n537), .ZN(n536) );
  INV_X1 U1750 ( .A(n435), .ZN(n662) );
  AOI21_X1 U1751 ( .B1(n565), .B2(n561), .A(n562), .ZN(n560) );
  NAND2_X1 U1752 ( .A1(n662), .A2(n436), .ZN(n311) );
  AOI21_X1 U1753 ( .B1(n662), .B2(n445), .A(n434), .ZN(n432) );
  INV_X1 U1754 ( .A(n436), .ZN(n434) );
  XNOR2_X1 U1755 ( .A(n504), .B(n317), .ZN(product[29]) );
  XNOR2_X1 U1756 ( .A(n497), .B(n316), .ZN(product[30]) );
  NAND2_X1 U1757 ( .A1(n667), .A2(n496), .ZN(n316) );
  XNOR2_X1 U1758 ( .A(n515), .B(n318), .ZN(product[28]) );
  NAND2_X1 U1759 ( .A1(n1994), .A2(n1942), .ZN(n318) );
  INV_X1 U1760 ( .A(n502), .ZN(n668) );
  INV_X1 U1761 ( .A(n563), .ZN(n561) );
  INV_X1 U1762 ( .A(n564), .ZN(n562) );
  INV_X1 U1763 ( .A(n438), .ZN(n663) );
  NAND2_X1 U1764 ( .A1(n2060), .A2(n670), .ZN(n516) );
  INV_X1 U1765 ( .A(n382), .ZN(n380) );
  NOR2_X1 U1766 ( .A1(n534), .A2(n531), .ZN(n525) );
  AOI21_X1 U1767 ( .B1(n581), .B2(n567), .A(n568), .ZN(n566) );
  AOI21_X1 U1768 ( .B1(n2130), .B2(n416), .A(n407), .ZN(n405) );
  INV_X1 U1769 ( .A(n409), .ZN(n407) );
  INV_X1 U1770 ( .A(n481), .ZN(n483) );
  INV_X1 U1771 ( .A(n521), .ZN(n519) );
  OAI21_X1 U1772 ( .B1(n600), .B2(n597), .A(n598), .ZN(n596) );
  OAI21_X1 U1773 ( .B1(n620), .B2(n610), .A(n611), .ZN(n609) );
  NAND2_X1 U1774 ( .A1(n671), .A2(n532), .ZN(n320) );
  NAND2_X1 U1775 ( .A1(n666), .A2(n481), .ZN(n315) );
  INV_X1 U1776 ( .A(n1992), .ZN(n670) );
  NAND2_X1 U1777 ( .A1(n941), .A2(n962), .ZN(n550) );
  NOR2_X1 U1778 ( .A1(n384), .A2(n364), .ZN(n362) );
  NAND2_X1 U1779 ( .A1(n2129), .A2(n378), .ZN(n305) );
  NAND2_X1 U1780 ( .A1(n2130), .A2(n409), .ZN(n308) );
  NAND2_X1 U1781 ( .A1(n422), .A2(n2128), .ZN(n411) );
  NAND2_X1 U1782 ( .A1(n657), .A2(n387), .ZN(n306) );
  INV_X1 U1783 ( .A(n384), .ZN(n657) );
  NAND2_X1 U1784 ( .A1(n2132), .A2(n396), .ZN(n307) );
  NAND2_X1 U1785 ( .A1(n661), .A2(n429), .ZN(n310) );
  INV_X1 U1786 ( .A(n428), .ZN(n661) );
  XOR2_X1 U1787 ( .A(n544), .B(n322), .Z(product[24]) );
  NAND2_X1 U1788 ( .A1(n673), .A2(n543), .ZN(n322) );
  AOI21_X1 U1789 ( .B1(n565), .B2(n545), .A(n546), .ZN(n544) );
  NOR2_X1 U1790 ( .A1(n737), .A2(n748), .ZN(n435) );
  AOI21_X1 U1791 ( .B1(n423), .B2(n2128), .A(n416), .ZN(n412) );
  INV_X1 U1792 ( .A(n480), .ZN(n666) );
  OAI21_X1 U1793 ( .B1(n492), .B2(n480), .A(n481), .ZN(n479) );
  NAND2_X1 U1794 ( .A1(n737), .A2(n748), .ZN(n436) );
  NOR2_X1 U1795 ( .A1(n1003), .A2(n1020), .ZN(n569) );
  XNOR2_X1 U1796 ( .A(n522), .B(n319), .ZN(product[27]) );
  NAND2_X1 U1797 ( .A1(n670), .A2(n1991), .ZN(n319) );
  INV_X1 U1798 ( .A(n378), .ZN(n376) );
  INV_X1 U1799 ( .A(n396), .ZN(n394) );
  NOR2_X1 U1800 ( .A1(n2065), .A2(n480), .ZN(n478) );
  NAND2_X1 U1801 ( .A1(n1003), .A2(n1020), .ZN(n570) );
  OR2_X1 U1802 ( .A1(n761), .A2(n774), .ZN(n2126) );
  NOR2_X1 U1803 ( .A1(n789), .A2(n804), .ZN(n480) );
  XNOR2_X1 U1804 ( .A(n2127), .B(n900), .ZN(n879) );
  XNOR2_X1 U1805 ( .A(n883), .B(n885), .ZN(n2127) );
  INV_X1 U1806 ( .A(n352), .ZN(n350) );
  NAND2_X1 U1807 ( .A1(n789), .A2(n804), .ZN(n481) );
  NOR2_X1 U1808 ( .A1(n695), .A2(n700), .ZN(n384) );
  NAND2_X1 U1809 ( .A1(n2133), .A2(n1978), .ZN(n599) );
  OR2_X1 U1810 ( .A1(n717), .A2(n726), .ZN(n2128) );
  OAI21_X1 U1811 ( .B1(n638), .B2(n636), .A(n637), .ZN(n635) );
  NAND2_X1 U1812 ( .A1(n2138), .A2(n369), .ZN(n304) );
  OR2_X1 U1813 ( .A1(n694), .A2(n689), .ZN(n2129) );
  AOI21_X1 U1814 ( .B1(n625), .B2(n1977), .A(n1969), .ZN(n620) );
  AOI21_X1 U1815 ( .B1(n2133), .B2(n1967), .A(n1973), .ZN(n600) );
  OAI21_X1 U1816 ( .B1(n405), .B2(n360), .A(n361), .ZN(n359) );
  AOI21_X1 U1817 ( .B1(n362), .B2(n394), .A(n363), .ZN(n361) );
  OAI21_X1 U1818 ( .B1(n364), .B2(n387), .A(n365), .ZN(n363) );
  AOI21_X1 U1819 ( .B1(n376), .B2(n2138), .A(n367), .ZN(n365) );
  AOI21_X1 U1820 ( .B1(n2131), .B2(n1968), .A(n1974), .ZN(n611) );
  OR2_X1 U1821 ( .A1(n709), .A2(n716), .ZN(n2130) );
  OR2_X1 U1822 ( .A1(n1133), .A2(n1142), .ZN(n2131) );
  NOR2_X1 U1823 ( .A1(n1071), .A2(n1084), .ZN(n590) );
  NAND2_X1 U1824 ( .A1(n2142), .A2(n341), .ZN(n302) );
  NAND2_X1 U1825 ( .A1(n2141), .A2(n352), .ZN(n303) );
  OR2_X1 U1826 ( .A1(n701), .A2(n708), .ZN(n2132) );
  NAND2_X1 U1827 ( .A1(n695), .A2(n700), .ZN(n387) );
  NOR2_X1 U1828 ( .A1(n1099), .A2(n1110), .ZN(n597) );
  NAND2_X1 U1829 ( .A1(n919), .A2(n940), .ZN(n543) );
  NAND2_X1 U1830 ( .A1(n727), .A2(n736), .ZN(n429) );
  NAND2_X1 U1831 ( .A1(n857), .A2(n876), .ZN(n521) );
  NAND2_X1 U1832 ( .A1(n701), .A2(n708), .ZN(n396) );
  OR2_X1 U1833 ( .A1(n1111), .A2(n1122), .ZN(n2133) );
  NAND2_X1 U1834 ( .A1(n2129), .A2(n2138), .ZN(n364) );
  OR2_X1 U1835 ( .A1(n1021), .A2(n1038), .ZN(n2256) );
  OR2_X1 U1836 ( .A1(n788), .A2(n775), .ZN(n2203) );
  INV_X1 U1837 ( .A(n369), .ZN(n367) );
  OR2_X1 U1838 ( .A1(n1055), .A2(n1070), .ZN(n2134) );
  NOR2_X1 U1839 ( .A1(n336), .A2(n334), .ZN(n332) );
  NAND2_X1 U1840 ( .A1(n1099), .A2(n1110), .ZN(n598) );
  NAND2_X1 U1841 ( .A1(n1980), .A2(n2131), .ZN(n610) );
  NAND2_X1 U1842 ( .A1(n2256), .A2(n1979), .ZN(n571) );
  XNOR2_X1 U1843 ( .A(n2135), .B(n1327), .ZN(n977) );
  XNOR2_X1 U1844 ( .A(n1305), .B(n1437), .ZN(n2135) );
  XNOR2_X1 U1845 ( .A(n906), .B(n2136), .ZN(n883) );
  XNOR2_X1 U1846 ( .A(n889), .B(n893), .ZN(n2136) );
  XNOR2_X1 U1847 ( .A(n2137), .B(n879), .ZN(n877) );
  XNOR2_X1 U1848 ( .A(n898), .B(n881), .ZN(n2137) );
  OR2_X1 U1849 ( .A1(n685), .A2(n688), .ZN(n2138) );
  BUF_X1 U1850 ( .A(n2072), .Z(n2178) );
  AOI21_X1 U1851 ( .B1(n643), .B2(n1965), .A(n1972), .ZN(n638) );
  OAI21_X1 U1852 ( .B1(n646), .B2(n644), .A(n645), .ZN(n643) );
  AOI21_X1 U1853 ( .B1(n1964), .B2(n1963), .A(n1971), .ZN(n646) );
  NAND2_X1 U1854 ( .A1(n678), .A2(n677), .ZN(n335) );
  INV_X1 U1855 ( .A(n341), .ZN(n339) );
  NOR2_X1 U1856 ( .A1(n1175), .A2(n1178), .ZN(n636) );
  XNOR2_X1 U1857 ( .A(n2139), .B(n1186), .ZN(n1095) );
  XNOR2_X1 U1858 ( .A(n1400), .B(n2050), .ZN(n2139) );
  XNOR2_X1 U1859 ( .A(n996), .B(n2140), .ZN(n973) );
  XNOR2_X1 U1860 ( .A(n994), .B(n1217), .ZN(n2140) );
  OR2_X1 U1861 ( .A1(n681), .A2(n684), .ZN(n2141) );
  OR2_X1 U1862 ( .A1(n679), .A2(n680), .ZN(n2142) );
  NAND2_X1 U1863 ( .A1(n681), .A2(n684), .ZN(n352) );
  NAND2_X1 U1864 ( .A1(n679), .A2(n680), .ZN(n341) );
  NAND2_X1 U1865 ( .A1(n1175), .A2(n1178), .ZN(n637) );
  NAND2_X1 U1866 ( .A1(n1159), .A2(n1161), .ZN(n627) );
  INV_X1 U1867 ( .A(n676), .ZN(n677) );
  NOR2_X1 U1868 ( .A1(n678), .A2(n677), .ZN(n334) );
  OR2_X1 U1869 ( .A1(n1194), .A2(n676), .ZN(n2143) );
  AND2_X1 U1870 ( .A1(n1194), .A2(n676), .ZN(n2144) );
  NAND2_X1 U1871 ( .A1(n2358), .A2(n2364), .ZN(n1756) );
  NAND2_X1 U1872 ( .A1(n2021), .A2(n2364), .ZN(n1606) );
  INV_X1 U1873 ( .A(n2343), .ZN(n2340) );
  INV_X1 U1874 ( .A(n2331), .ZN(n2329) );
  INV_X1 U1875 ( .A(n2338), .ZN(n2335) );
  INV_X1 U1876 ( .A(n2349), .ZN(n2346) );
  INV_X1 U1877 ( .A(n2011), .ZN(n2323) );
  INV_X1 U1878 ( .A(n1682), .ZN(n2368) );
  XOR2_X1 U1879 ( .A(n2145), .B(n1096), .Z(n1079) );
  XOR2_X1 U1880 ( .A(n1399), .B(n1421), .Z(n2145) );
  INV_X1 U1881 ( .A(n1956), .ZN(n2283) );
  INV_X1 U1882 ( .A(n2154), .ZN(n2288) );
  INV_X1 U1883 ( .A(n1507), .ZN(n2375) );
  NAND2_X1 U1884 ( .A1(n2352), .A2(n2364), .ZN(n1731) );
  INV_X1 U1885 ( .A(n682), .ZN(n683) );
  INV_X1 U1886 ( .A(n2198), .ZN(n2293) );
  INV_X1 U1887 ( .A(n2017), .ZN(n2287) );
  INV_X1 U1888 ( .A(n2194), .ZN(n2298) );
  INV_X1 U1889 ( .A(n1993), .ZN(n2297) );
  INV_X1 U1890 ( .A(n2198), .ZN(n2292) );
  INV_X1 U1891 ( .A(n2354), .ZN(n2351) );
  INV_X1 U1892 ( .A(n2331), .ZN(n2328) );
  NOR2_X1 U1893 ( .A1(n2289), .A2(n2364), .ZN(n1289) );
  NOR2_X1 U1894 ( .A1(n2296), .A2(n2364), .ZN(n1385) );
  NOR2_X1 U1895 ( .A1(n2300), .A2(n2364), .ZN(n1433) );
  NOR2_X1 U1896 ( .A1(n2301), .A2(n2364), .ZN(n1457) );
  OR2_X1 U1897 ( .A1(n2146), .A2(n2147), .ZN(n1390) );
  NOR2_X1 U1898 ( .A1(n1984), .A2(n1687), .ZN(n2146) );
  NOR2_X1 U1899 ( .A1(n1686), .A2(n2036), .ZN(n2147) );
  NOR2_X1 U1900 ( .A1(n2033), .A2(n1646), .ZN(n2148) );
  NOR2_X1 U1901 ( .A1(n1985), .A2(n1645), .ZN(n2149) );
  INV_X1 U1902 ( .A(n2161), .ZN(n2276) );
  NAND2_X1 U1903 ( .A1(n1181), .A2(n1192), .ZN(n645) );
  NOR2_X1 U1904 ( .A1(n1181), .A2(n1192), .ZN(n644) );
  INV_X1 U1905 ( .A(n1632), .ZN(n2370) );
  INV_X1 U1906 ( .A(n1532), .ZN(n2374) );
  NOR2_X1 U1907 ( .A1(n2297), .A2(n2364), .ZN(n1409) );
  NAND2_X1 U1908 ( .A1(n2335), .A2(n2364), .ZN(n1656) );
  NAND2_X1 U1909 ( .A1(n2328), .A2(n2364), .ZN(n1631) );
  NAND2_X1 U1910 ( .A1(n2317), .A2(n2364), .ZN(n1581) );
  NAND2_X1 U1911 ( .A1(n2096), .A2(n2364), .ZN(n1556) );
  NAND2_X1 U1912 ( .A1(n2310), .A2(n2364), .ZN(n1531) );
  NAND2_X1 U1913 ( .A1(n2346), .A2(n2364), .ZN(n1706) );
  NAND2_X1 U1914 ( .A1(n2340), .A2(n2364), .ZN(n1681) );
  OR2_X1 U1915 ( .A1(n2150), .A2(n2151), .ZN(n1306) );
  NOR2_X1 U1916 ( .A1(n1939), .A2(n1599), .ZN(n2150) );
  NOR2_X1 U1917 ( .A1(n1598), .A2(n2291), .ZN(n2151) );
  NOR2_X1 U1918 ( .A1(n2290), .A2(n2364), .ZN(n1313) );
  NOR2_X1 U1919 ( .A1(n2295), .A2(n2364), .ZN(n1361) );
  NOR2_X1 U1920 ( .A1(n2288), .A2(n2364), .ZN(n1265) );
  NOR2_X1 U1921 ( .A1(n2285), .A2(n2364), .ZN(n1241) );
  INV_X1 U1922 ( .A(n1707), .ZN(n2367) );
  INV_X1 U1923 ( .A(n802), .ZN(n803) );
  INV_X1 U1924 ( .A(n724), .ZN(n725) );
  NOR2_X1 U1925 ( .A1(n2024), .A2(n2364), .ZN(n1337) );
  OAI22_X1 U1926 ( .A1(n2241), .A2(n1534), .B1(n2287), .B2(n1533), .ZN(n1243)
         );
  INV_X1 U1927 ( .A(n1557), .ZN(n2373) );
  INV_X1 U1928 ( .A(n1607), .ZN(n2371) );
  OAI22_X1 U1929 ( .A1(n2241), .A2(n1538), .B1(n2287), .B2(n1537), .ZN(n1247)
         );
  XNOR2_X1 U1930 ( .A(n1000), .B(n2152), .ZN(n975) );
  XNOR2_X1 U1931 ( .A(n1393), .B(n1415), .ZN(n2152) );
  NAND2_X1 U1932 ( .A1(n2028), .A2(n2364), .ZN(n1781) );
  INV_X1 U1933 ( .A(n1732), .ZN(n2366) );
  INV_X1 U1934 ( .A(n1582), .ZN(n2372) );
  INV_X1 U1935 ( .A(n1657), .ZN(n2369) );
  INV_X1 U1936 ( .A(n1482), .ZN(n2376) );
  XNOR2_X1 U1937 ( .A(n2335), .B(b[0]), .ZN(n1655) );
  XNOR2_X1 U1938 ( .A(n2358), .B(b[0]), .ZN(n1755) );
  XNOR2_X1 U1939 ( .A(n2329), .B(b[0]), .ZN(n1630) );
  XNOR2_X1 U1940 ( .A(n2353), .B(b[0]), .ZN(n1730) );
  XNOR2_X1 U1941 ( .A(n2318), .B(b[0]), .ZN(n1580) );
  XNOR2_X1 U1942 ( .A(n2315), .B(b[22]), .ZN(n1533) );
  XNOR2_X1 U1943 ( .A(n2314), .B(b[18]), .ZN(n1537) );
  XNOR2_X1 U1944 ( .A(a[22]), .B(n2312), .ZN(n2244) );
  XNOR2_X1 U1945 ( .A(n2361), .B(b[22]), .ZN(n1758) );
  XNOR2_X1 U1946 ( .A(n2029), .B(b[16]), .ZN(n1764) );
  XNOR2_X1 U1947 ( .A(n2361), .B(b[20]), .ZN(n1760) );
  XNOR2_X1 U1948 ( .A(n2029), .B(b[12]), .ZN(n1768) );
  XNOR2_X1 U1949 ( .A(n2360), .B(b[8]), .ZN(n1772) );
  XNOR2_X1 U1950 ( .A(n2028), .B(b[14]), .ZN(n1766) );
  XNOR2_X1 U1951 ( .A(n2356), .B(b[22]), .ZN(n1733) );
  XNOR2_X1 U1952 ( .A(n2335), .B(b[12]), .ZN(n1643) );
  XNOR2_X1 U1953 ( .A(n2336), .B(b[14]), .ZN(n1641) );
  XNOR2_X1 U1954 ( .A(n2340), .B(b[14]), .ZN(n1666) );
  XNOR2_X1 U1955 ( .A(n2317), .B(b[8]), .ZN(n1572) );
  XNOR2_X1 U1956 ( .A(n2346), .B(b[12]), .ZN(n1693) );
  XNOR2_X1 U1957 ( .A(n2340), .B(b[12]), .ZN(n1668) );
  XNOR2_X1 U1958 ( .A(n2020), .B(b[8]), .ZN(n1597) );
  XNOR2_X1 U1959 ( .A(n2044), .B(b[8]), .ZN(n1622) );
  XNOR2_X1 U1960 ( .A(n2353), .B(b[16]), .ZN(n1714) );
  XNOR2_X1 U1961 ( .A(n2358), .B(b[20]), .ZN(n1735) );
  XNOR2_X1 U1962 ( .A(n2353), .B(b[20]), .ZN(n1710) );
  XNOR2_X1 U1963 ( .A(n2347), .B(b[16]), .ZN(n1689) );
  XNOR2_X1 U1964 ( .A(n2045), .B(b[12]), .ZN(n1618) );
  XNOR2_X1 U1965 ( .A(n2347), .B(b[22]), .ZN(n1683) );
  XNOR2_X1 U1966 ( .A(n2318), .B(b[22]), .ZN(n1558) );
  XNOR2_X1 U1967 ( .A(n2328), .B(b[14]), .ZN(n1616) );
  XNOR2_X1 U1968 ( .A(n2357), .B(b[14]), .ZN(n1741) );
  XNOR2_X1 U1969 ( .A(n2341), .B(b[22]), .ZN(n1658) );
  XNOR2_X1 U1970 ( .A(n2357), .B(b[12]), .ZN(n1743) );
  XNOR2_X1 U1971 ( .A(n2346), .B(b[14]), .ZN(n1691) );
  XNOR2_X1 U1972 ( .A(n2347), .B(b[20]), .ZN(n1685) );
  XNOR2_X1 U1973 ( .A(n2045), .B(b[22]), .ZN(n1608) );
  XNOR2_X1 U1974 ( .A(n2341), .B(b[16]), .ZN(n1664) );
  XNOR2_X1 U1975 ( .A(n2315), .B(b[8]), .ZN(n1547) );
  XNOR2_X1 U1976 ( .A(n2323), .B(b[12]), .ZN(n1593) );
  XNOR2_X1 U1977 ( .A(n2045), .B(b[16]), .ZN(n1614) );
  XNOR2_X1 U1978 ( .A(n2317), .B(b[12]), .ZN(n1568) );
  XNOR2_X1 U1979 ( .A(n2353), .B(b[22]), .ZN(n1708) );
  XNOR2_X1 U1980 ( .A(n2336), .B(b[8]), .ZN(n1647) );
  XNOR2_X1 U1981 ( .A(n2336), .B(b[22]), .ZN(n1633) );
  XNOR2_X1 U1982 ( .A(n2340), .B(b[8]), .ZN(n1672) );
  XNOR2_X1 U1983 ( .A(n2336), .B(b[16]), .ZN(n1639) );
  XNOR2_X1 U1984 ( .A(n2358), .B(b[16]), .ZN(n1739) );
  XNOR2_X1 U1985 ( .A(n2021), .B(b[14]), .ZN(n1591) );
  XNOR2_X1 U1986 ( .A(n2346), .B(b[8]), .ZN(n1697) );
  XNOR2_X1 U1987 ( .A(n2315), .B(b[16]), .ZN(n1539) );
  XNOR2_X1 U1988 ( .A(n2323), .B(b[20]), .ZN(n1585) );
  XNOR2_X1 U1989 ( .A(n2352), .B(b[14]), .ZN(n1716) );
  XNOR2_X1 U1990 ( .A(n2310), .B(b[8]), .ZN(n1522) );
  XNOR2_X1 U1991 ( .A(n2357), .B(b[8]), .ZN(n1747) );
  XNOR2_X1 U1992 ( .A(n2045), .B(b[20]), .ZN(n1610) );
  XNOR2_X1 U1993 ( .A(n2352), .B(b[8]), .ZN(n1722) );
  XNOR2_X1 U1994 ( .A(n2310), .B(b[14]), .ZN(n1516) );
  XNOR2_X1 U1995 ( .A(n2352), .B(b[12]), .ZN(n1718) );
  XNOR2_X1 U1996 ( .A(n2315), .B(b[14]), .ZN(n1541) );
  XNOR2_X1 U1997 ( .A(n2323), .B(b[22]), .ZN(n1583) );
  XNOR2_X1 U1998 ( .A(n2318), .B(b[16]), .ZN(n1564) );
  XNOR2_X1 U1999 ( .A(n2095), .B(b[12]), .ZN(n1543) );
  XNOR2_X1 U2000 ( .A(n2020), .B(b[16]), .ZN(n1589) );
  XNOR2_X1 U2001 ( .A(n2311), .B(b[22]), .ZN(n1508) );
  XNOR2_X1 U2002 ( .A(n2336), .B(b[20]), .ZN(n1635) );
  XNOR2_X1 U2003 ( .A(n2311), .B(b[20]), .ZN(n1510) );
  XNOR2_X1 U2004 ( .A(n2310), .B(b[12]), .ZN(n1518) );
  XNOR2_X1 U2005 ( .A(n2317), .B(b[14]), .ZN(n1566) );
  XNOR2_X1 U2006 ( .A(n2311), .B(b[16]), .ZN(n1514) );
  XNOR2_X1 U2007 ( .A(n2318), .B(b[20]), .ZN(n1560) );
  XNOR2_X1 U2008 ( .A(n2341), .B(b[20]), .ZN(n1660) );
  XNOR2_X1 U2009 ( .A(n2315), .B(b[20]), .ZN(n1535) );
  XNOR2_X1 U2010 ( .A(n2361), .B(b[18]), .ZN(n1762) );
  XNOR2_X1 U2011 ( .A(n2028), .B(b[10]), .ZN(n1770) );
  XNOR2_X1 U2012 ( .A(n2360), .B(b[2]), .ZN(n1778) );
  XNOR2_X1 U2013 ( .A(n2029), .B(b[4]), .ZN(n1776) );
  XNOR2_X1 U2014 ( .A(n2310), .B(b[4]), .ZN(n1526) );
  XNOR2_X1 U2015 ( .A(n2356), .B(b[18]), .ZN(n1737) );
  XNOR2_X1 U2016 ( .A(n2310), .B(b[2]), .ZN(n1528) );
  XNOR2_X1 U2017 ( .A(n2095), .B(b[4]), .ZN(n1551) );
  XNOR2_X1 U2018 ( .A(n2352), .B(b[18]), .ZN(n1712) );
  XNOR2_X1 U2019 ( .A(n2324), .B(b[10]), .ZN(n1595) );
  XNOR2_X1 U2020 ( .A(n2317), .B(b[2]), .ZN(n1578) );
  XNOR2_X1 U2021 ( .A(n2330), .B(b[2]), .ZN(n1628) );
  XNOR2_X1 U2022 ( .A(n2346), .B(b[2]), .ZN(n1703) );
  XNOR2_X1 U2023 ( .A(n2340), .B(b[18]), .ZN(n1662) );
  XNOR2_X1 U2024 ( .A(n2021), .B(b[2]), .ZN(n1603) );
  XNOR2_X1 U2025 ( .A(n2324), .B(b[4]), .ZN(n1601) );
  XNOR2_X1 U2026 ( .A(n2335), .B(b[4]), .ZN(n1651) );
  XNOR2_X1 U2027 ( .A(n2335), .B(b[18]), .ZN(n1637) );
  XNOR2_X1 U2028 ( .A(n2095), .B(b[10]), .ZN(n1545) );
  XNOR2_X1 U2029 ( .A(n2336), .B(b[2]), .ZN(n1653) );
  XNOR2_X1 U2030 ( .A(n2310), .B(b[18]), .ZN(n1512) );
  XNOR2_X1 U2031 ( .A(n2329), .B(b[4]), .ZN(n1626) );
  XNOR2_X1 U2032 ( .A(n2340), .B(b[10]), .ZN(n1670) );
  XNOR2_X1 U2033 ( .A(n2317), .B(b[10]), .ZN(n1570) );
  XNOR2_X1 U2034 ( .A(n2330), .B(b[10]), .ZN(n1620) );
  XNOR2_X1 U2035 ( .A(n2357), .B(b[10]), .ZN(n1745) );
  XNOR2_X1 U2036 ( .A(n2340), .B(b[4]), .ZN(n1676) );
  XNOR2_X1 U2037 ( .A(n2340), .B(b[2]), .ZN(n1678) );
  XNOR2_X1 U2038 ( .A(n2324), .B(b[18]), .ZN(n1587) );
  XNOR2_X1 U2039 ( .A(n2358), .B(b[4]), .ZN(n1751) );
  XNOR2_X1 U2040 ( .A(n2346), .B(b[10]), .ZN(n1695) );
  XNOR2_X1 U2041 ( .A(n2346), .B(b[4]), .ZN(n1701) );
  XNOR2_X1 U2042 ( .A(n2352), .B(b[4]), .ZN(n1726) );
  XNOR2_X1 U2043 ( .A(n2317), .B(b[18]), .ZN(n1562) );
  XNOR2_X1 U2044 ( .A(n2330), .B(b[18]), .ZN(n1612) );
  XNOR2_X1 U2045 ( .A(n2352), .B(b[2]), .ZN(n1728) );
  XNOR2_X1 U2046 ( .A(n2357), .B(b[2]), .ZN(n1753) );
  XNOR2_X1 U2047 ( .A(n2310), .B(b[10]), .ZN(n1520) );
  XNOR2_X1 U2048 ( .A(n2352), .B(b[10]), .ZN(n1720) );
  XNOR2_X1 U2049 ( .A(n2347), .B(b[0]), .ZN(n1705) );
  XNOR2_X1 U2050 ( .A(n2028), .B(b[6]), .ZN(n1774) );
  XNOR2_X1 U2051 ( .A(n2317), .B(b[6]), .ZN(n1574) );
  XNOR2_X1 U2052 ( .A(n2352), .B(b[6]), .ZN(n1724) );
  XNOR2_X1 U2053 ( .A(n2045), .B(b[6]), .ZN(n1624) );
  XNOR2_X1 U2054 ( .A(n2335), .B(b[6]), .ZN(n1649) );
  XNOR2_X1 U2055 ( .A(n2310), .B(b[6]), .ZN(n1524) );
  XNOR2_X1 U2056 ( .A(n2346), .B(b[6]), .ZN(n1699) );
  XNOR2_X1 U2057 ( .A(n2358), .B(b[6]), .ZN(n1749) );
  XNOR2_X1 U2058 ( .A(n2340), .B(b[6]), .ZN(n1674) );
  XOR2_X1 U2059 ( .A(a[18]), .B(a[17]), .Z(n2154) );
  XNOR2_X1 U2060 ( .A(b[23]), .B(n2052), .ZN(n1557) );
  XNOR2_X1 U2061 ( .A(b[23]), .B(n2328), .ZN(n1607) );
  XNOR2_X1 U2062 ( .A(b[23]), .B(n2008), .ZN(n1707) );
  XNOR2_X1 U2063 ( .A(b[23]), .B(n2334), .ZN(n1632) );
  XNOR2_X1 U2064 ( .A(b[23]), .B(n2339), .ZN(n1657) );
  XNOR2_X1 U2065 ( .A(n2311), .B(b[0]), .ZN(n1530) );
  XNOR2_X1 U2066 ( .A(b[1]), .B(n2305), .ZN(n1504) );
  XNOR2_X1 U2067 ( .A(b[7]), .B(n2052), .ZN(n1573) );
  XNOR2_X1 U2068 ( .A(b[3]), .B(n2052), .ZN(n1577) );
  XNOR2_X1 U2069 ( .A(b[3]), .B(n2001), .ZN(n1502) );
  XNOR2_X1 U2070 ( .A(b[1]), .B(n2052), .ZN(n1579) );
  XNOR2_X1 U2071 ( .A(b[7]), .B(n2008), .ZN(n1723) );
  XNOR2_X1 U2072 ( .A(b[3]), .B(n2329), .ZN(n1627) );
  XNOR2_X1 U2073 ( .A(b[7]), .B(n2330), .ZN(n1623) );
  XNOR2_X1 U2074 ( .A(b[1]), .B(n2339), .ZN(n1679) );
  XNOR2_X1 U2075 ( .A(b[7]), .B(n2334), .ZN(n1648) );
  XNOR2_X1 U2076 ( .A(b[7]), .B(n2339), .ZN(n1673) );
  XNOR2_X1 U2077 ( .A(b[7]), .B(n2002), .ZN(n1498) );
  XNOR2_X1 U2078 ( .A(b[1]), .B(n2334), .ZN(n1654) );
  XNOR2_X1 U2079 ( .A(b[3]), .B(n2339), .ZN(n1677) );
  XNOR2_X1 U2080 ( .A(b[3]), .B(n2005), .ZN(n1652) );
  XNOR2_X1 U2081 ( .A(b[1]), .B(n2044), .ZN(n1629) );
  XNOR2_X1 U2082 ( .A(b[1]), .B(n2008), .ZN(n1729) );
  XNOR2_X1 U2083 ( .A(b[3]), .B(n2008), .ZN(n1727) );
  XNOR2_X1 U2084 ( .A(b[9]), .B(n2052), .ZN(n1571) );
  XNOR2_X1 U2085 ( .A(b[9]), .B(n2329), .ZN(n1621) );
  XNOR2_X1 U2086 ( .A(b[5]), .B(n2002), .ZN(n1500) );
  XNOR2_X1 U2087 ( .A(b[9]), .B(n2339), .ZN(n1671) );
  XNOR2_X1 U2088 ( .A(b[5]), .B(n2334), .ZN(n1650) );
  XNOR2_X1 U2089 ( .A(b[5]), .B(n2328), .ZN(n1625) );
  XNOR2_X1 U2090 ( .A(b[5]), .B(n2339), .ZN(n1675) );
  XNOR2_X1 U2091 ( .A(b[5]), .B(n2008), .ZN(n1725) );
  XNOR2_X1 U2092 ( .A(b[9]), .B(n2002), .ZN(n1496) );
  XNOR2_X1 U2093 ( .A(b[9]), .B(n2008), .ZN(n1721) );
  XNOR2_X1 U2094 ( .A(b[17]), .B(n2001), .ZN(n1488) );
  XNOR2_X1 U2095 ( .A(b[13]), .B(n2001), .ZN(n1492) );
  XNOR2_X1 U2096 ( .A(b[11]), .B(n2001), .ZN(n1494) );
  XNOR2_X1 U2097 ( .A(b[15]), .B(n2002), .ZN(n1490) );
  XNOR2_X1 U2098 ( .A(b[19]), .B(n2001), .ZN(n1486) );
  XNOR2_X1 U2099 ( .A(b[21]), .B(n2002), .ZN(n1484) );
  INV_X1 U2100 ( .A(n1757), .ZN(n2365) );
  XNOR2_X1 U2101 ( .A(n2029), .B(b[0]), .ZN(n1780) );
  XNOR2_X1 U2102 ( .A(a[2]), .B(a[3]), .ZN(n2160) );
  XNOR2_X1 U2103 ( .A(n2020), .B(b[0]), .ZN(n1605) );
  XNOR2_X1 U2104 ( .A(a[4]), .B(n2350), .ZN(n2163) );
  XNOR2_X1 U2105 ( .A(a[10]), .B(n2333), .ZN(n2165) );
  XOR2_X1 U2106 ( .A(a[22]), .B(n2307), .Z(n2167) );
  INV_X1 U2107 ( .A(a[5]), .ZN(n2354) );
  INV_X1 U2108 ( .A(a[11]), .ZN(n2337) );
  XNOR2_X1 U2109 ( .A(n2315), .B(b[0]), .ZN(n1555) );
  XNOR2_X1 U2110 ( .A(a[12]), .B(n2327), .ZN(n2171) );
  XNOR2_X1 U2111 ( .A(n2341), .B(b[0]), .ZN(n1680) );
  XNOR2_X1 U2112 ( .A(a[16]), .B(a[17]), .ZN(n2174) );
  XNOR2_X1 U2113 ( .A(b[23]), .B(n2001), .ZN(n1482) );
  INV_X1 U2114 ( .A(n2161), .ZN(n2277) );
  NOR2_X1 U2115 ( .A1(n821), .A2(n838), .ZN(n502) );
  NAND2_X1 U2116 ( .A1(n963), .A2(n982), .ZN(n559) );
  INV_X1 U2117 ( .A(n2162), .ZN(n2279) );
  AOI21_X1 U2118 ( .B1(n2086), .B2(n670), .A(n519), .ZN(n517) );
  INV_X1 U2119 ( .A(n2086), .ZN(n524) );
  OAI21_X1 U2120 ( .B1(n531), .B2(n535), .A(n532), .ZN(n526) );
  NAND2_X1 U2121 ( .A1(n883), .A2(n885), .ZN(n2181) );
  NAND2_X1 U2122 ( .A1(n883), .A2(n900), .ZN(n2182) );
  NAND2_X1 U2123 ( .A1(n885), .A2(n900), .ZN(n2183) );
  NAND3_X1 U2124 ( .A1(n2181), .A2(n2182), .A3(n2183), .ZN(n878) );
  NAND2_X1 U2125 ( .A1(n898), .A2(n881), .ZN(n2184) );
  NAND2_X1 U2126 ( .A1(n898), .A2(n879), .ZN(n2185) );
  NAND2_X1 U2127 ( .A1(n881), .A2(n879), .ZN(n2186) );
  NAND3_X1 U2128 ( .A1(n2184), .A2(n2185), .A3(n2186), .ZN(n876) );
  INV_X1 U2129 ( .A(n2158), .ZN(n2294) );
  XOR2_X1 U2130 ( .A(n979), .B(n998), .Z(n2187) );
  XOR2_X1 U2131 ( .A(n2187), .B(n2069), .Z(n971) );
  NAND2_X1 U2132 ( .A1(n1305), .A2(n1437), .ZN(n2188) );
  NAND2_X1 U2133 ( .A1(n1305), .A2(n1327), .ZN(n2189) );
  NAND2_X1 U2134 ( .A1(n1437), .A2(n1327), .ZN(n2190) );
  NAND3_X1 U2135 ( .A1(n2188), .A2(n2189), .A3(n2190), .ZN(n976) );
  NAND2_X1 U2136 ( .A1(n998), .A2(n979), .ZN(n2191) );
  NAND2_X1 U2137 ( .A1(n998), .A2(n977), .ZN(n2192) );
  NAND2_X1 U2138 ( .A1(n979), .A2(n977), .ZN(n2193) );
  NAND3_X1 U2139 ( .A1(n2191), .A2(n2192), .A3(n2193), .ZN(n970) );
  AOI21_X1 U2140 ( .B1(n589), .B2(n2134), .A(n1975), .ZN(n583) );
  NAND2_X1 U2141 ( .A1(n588), .A2(n2134), .ZN(n582) );
  NAND2_X1 U2142 ( .A1(n2128), .A2(n2130), .ZN(n402) );
  NAND2_X1 U2143 ( .A1(n1351), .A2(n1263), .ZN(n2195) );
  NAND2_X1 U2144 ( .A1(n1351), .A2(n1285), .ZN(n2196) );
  NAND2_X1 U2145 ( .A1(n1263), .A2(n1285), .ZN(n2197) );
  NAND3_X1 U2146 ( .A1(n2195), .A2(n2196), .A3(n2197), .ZN(n1018) );
  XNOR2_X1 U2147 ( .A(b[9]), .B(n2334), .ZN(n1646) );
  XNOR2_X1 U2148 ( .A(n2335), .B(b[10]), .ZN(n1645) );
  OAI21_X1 U2149 ( .B1(a[0]), .B2(n2172), .A(n2365), .ZN(n1458) );
  INV_X1 U2150 ( .A(a[0]), .ZN(n251) );
  XNOR2_X1 U2151 ( .A(b[23]), .B(n2309), .ZN(n1507) );
  XNOR2_X1 U2152 ( .A(b[9]), .B(n2309), .ZN(n1521) );
  XNOR2_X1 U2153 ( .A(b[1]), .B(n2309), .ZN(n1529) );
  XNOR2_X1 U2154 ( .A(b[7]), .B(n2309), .ZN(n1523) );
  XNOR2_X1 U2155 ( .A(b[5]), .B(n2309), .ZN(n1525) );
  XNOR2_X1 U2156 ( .A(b[3]), .B(n2309), .ZN(n1527) );
  XNOR2_X1 U2157 ( .A(b[23]), .B(n2095), .ZN(n1532) );
  XNOR2_X1 U2158 ( .A(b[9]), .B(n2095), .ZN(n1546) );
  XNOR2_X1 U2159 ( .A(b[7]), .B(n2096), .ZN(n1548) );
  XNOR2_X1 U2160 ( .A(b[1]), .B(n2095), .ZN(n1554) );
  INV_X1 U2161 ( .A(a[23]), .ZN(n2307) );
  NAND2_X1 U2162 ( .A1(n950), .A2(n935), .ZN(n2200) );
  NAND2_X1 U2163 ( .A1(n950), .A2(n931), .ZN(n2201) );
  NAND2_X1 U2164 ( .A1(n935), .A2(n931), .ZN(n2202) );
  NAND3_X1 U2165 ( .A1(n2200), .A2(n2201), .A3(n2202), .ZN(n924) );
  AOI21_X1 U2166 ( .B1(n359), .B2(n2141), .A(n350), .ZN(n348) );
  NOR2_X1 U2167 ( .A1(n1936), .A2(n1550), .ZN(n2206) );
  NOR2_X1 U2168 ( .A1(n2288), .A2(n1549), .ZN(n2207) );
  OR2_X1 U2169 ( .A1(n2206), .A2(n2207), .ZN(n1259) );
  XNOR2_X1 U2170 ( .A(b[5]), .B(n2096), .ZN(n1550) );
  XNOR2_X1 U2171 ( .A(n2315), .B(b[6]), .ZN(n1549) );
  OAI22_X1 U2172 ( .A1(n2241), .A2(n1536), .B1(n2287), .B2(n1535), .ZN(n1245)
         );
  OAI22_X1 U2173 ( .A1(n2241), .A2(n1542), .B1(n2287), .B2(n1541), .ZN(n1251)
         );
  OAI22_X1 U2174 ( .A1(n1936), .A2(n1540), .B1(n2287), .B2(n1539), .ZN(n1249)
         );
  NAND2_X1 U2175 ( .A1(n2126), .A2(n461), .ZN(n313) );
  INV_X1 U2176 ( .A(n461), .ZN(n459) );
  INV_X1 U2177 ( .A(n692), .ZN(n693) );
  NAND2_X1 U2178 ( .A1(n685), .A2(n688), .ZN(n369) );
  NOR2_X1 U2179 ( .A1(n597), .A2(n599), .ZN(n595) );
  XNOR2_X1 U2180 ( .A(b[1]), .B(n2345), .ZN(n1704) );
  XNOR2_X1 U2181 ( .A(b[5]), .B(n2345), .ZN(n1700) );
  XNOR2_X1 U2182 ( .A(b[3]), .B(n2345), .ZN(n1702) );
  XNOR2_X1 U2183 ( .A(b[7]), .B(n2345), .ZN(n1698) );
  XNOR2_X1 U2184 ( .A(b[23]), .B(n2345), .ZN(n1682) );
  XNOR2_X1 U2185 ( .A(b[9]), .B(n2345), .ZN(n1696) );
  XNOR2_X1 U2186 ( .A(n2209), .B(n1390), .ZN(n909) );
  XNOR2_X1 U2187 ( .A(n1368), .B(n938), .ZN(n2209) );
  XNOR2_X1 U2188 ( .A(b[3]), .B(n2322), .ZN(n1602) );
  XNOR2_X1 U2189 ( .A(b[23]), .B(n2322), .ZN(n1582) );
  XNOR2_X1 U2190 ( .A(b[5]), .B(n2322), .ZN(n1600) );
  XNOR2_X1 U2191 ( .A(b[1]), .B(n2322), .ZN(n1604) );
  XNOR2_X1 U2192 ( .A(b[9]), .B(n2322), .ZN(n1596) );
  XNOR2_X1 U2193 ( .A(n2210), .B(n834), .ZN(n813) );
  XNOR2_X1 U2194 ( .A(n830), .B(n1386), .ZN(n2210) );
  OAI21_X1 U2195 ( .B1(n2173), .B2(n2043), .A(n2373), .ZN(n1266) );
  OAI21_X1 U2196 ( .B1(n2110), .B2(n1958), .A(n2375), .ZN(n1218) );
  XNOR2_X1 U2197 ( .A(n1949), .B(b[22]), .ZN(n1483) );
  XNOR2_X1 U2198 ( .A(n1949), .B(b[18]), .ZN(n1487) );
  XNOR2_X1 U2199 ( .A(n1949), .B(b[10]), .ZN(n1495) );
  NAND2_X1 U2200 ( .A1(n1949), .A2(n2364), .ZN(n1506) );
  XNOR2_X1 U2201 ( .A(n1949), .B(b[20]), .ZN(n1485) );
  XNOR2_X1 U2202 ( .A(n1949), .B(b[6]), .ZN(n1499) );
  XNOR2_X1 U2203 ( .A(n1949), .B(b[12]), .ZN(n1493) );
  XNOR2_X1 U2204 ( .A(n1949), .B(b[4]), .ZN(n1501) );
  XNOR2_X1 U2205 ( .A(n1949), .B(b[14]), .ZN(n1491) );
  XNOR2_X1 U2206 ( .A(n1949), .B(b[16]), .ZN(n1489) );
  XNOR2_X1 U2207 ( .A(n1949), .B(b[8]), .ZN(n1497) );
  XNOR2_X1 U2208 ( .A(n1949), .B(b[0]), .ZN(n1505) );
  XNOR2_X1 U2209 ( .A(n1948), .B(b[2]), .ZN(n1503) );
  OAI21_X1 U2210 ( .B1(n2166), .B2(n2244), .A(n2376), .ZN(n1194) );
  NOR2_X1 U2211 ( .A1(n435), .A2(n428), .ZN(n426) );
  INV_X1 U2212 ( .A(n2354), .ZN(n2350) );
  INV_X1 U2213 ( .A(n2332), .ZN(n2327) );
  NAND2_X1 U2214 ( .A1(n830), .A2(n1386), .ZN(n2211) );
  NAND2_X1 U2215 ( .A1(n830), .A2(n834), .ZN(n2212) );
  NAND2_X1 U2216 ( .A1(n1386), .A2(n834), .ZN(n2213) );
  NAND3_X1 U2217 ( .A1(n2211), .A2(n2212), .A3(n2213), .ZN(n812) );
  XOR2_X1 U2218 ( .A(n2214), .B(n2073), .Z(n793) );
  NAND2_X1 U2219 ( .A1(n801), .A2(n797), .ZN(n2215) );
  NAND2_X1 U2220 ( .A1(n801), .A2(n2073), .ZN(n2216) );
  NAND2_X1 U2221 ( .A1(n797), .A2(n812), .ZN(n2217) );
  NAND3_X1 U2222 ( .A1(n2215), .A2(n2216), .A3(n2217), .ZN(n792) );
  NAND2_X1 U2223 ( .A1(n749), .A2(n760), .ZN(n439) );
  NOR2_X1 U2224 ( .A1(n749), .A2(n760), .ZN(n438) );
  NAND2_X1 U2225 ( .A1(n1400), .A2(n1467), .ZN(n2218) );
  NAND2_X1 U2226 ( .A1(n1467), .A2(n1186), .ZN(n2219) );
  NAND2_X1 U2227 ( .A1(n1400), .A2(n1186), .ZN(n2220) );
  NAND3_X1 U2228 ( .A1(n2218), .A2(n2219), .A3(n2220), .ZN(n1094) );
  NAND2_X1 U2229 ( .A1(n1092), .A2(n1289), .ZN(n2221) );
  NAND2_X1 U2230 ( .A1(n1092), .A2(n1094), .ZN(n2222) );
  NAND2_X1 U2231 ( .A1(n1289), .A2(n1094), .ZN(n2223) );
  NAND3_X1 U2232 ( .A1(n2221), .A2(n2222), .A3(n2223), .ZN(n1076) );
  AOI21_X1 U2233 ( .B1(n2256), .B2(n1966), .A(n1976), .ZN(n572) );
  NAND2_X1 U2234 ( .A1(n1390), .A2(n938), .ZN(n2224) );
  NAND2_X1 U2235 ( .A1(n1390), .A2(n1368), .ZN(n2225) );
  NAND2_X1 U2236 ( .A1(n938), .A2(n1368), .ZN(n2226) );
  NAND3_X1 U2237 ( .A1(n2224), .A2(n2225), .A3(n2226), .ZN(n908) );
  XNOR2_X1 U2238 ( .A(n2346), .B(b[18]), .ZN(n1687) );
  NAND2_X1 U2239 ( .A1(n906), .A2(n889), .ZN(n2227) );
  NAND2_X1 U2240 ( .A1(n906), .A2(n893), .ZN(n2228) );
  NAND2_X1 U2241 ( .A1(n889), .A2(n893), .ZN(n2229) );
  NAND3_X1 U2242 ( .A1(n2227), .A2(n2228), .A3(n2229), .ZN(n882) );
  INV_X1 U2243 ( .A(n2337), .ZN(n2333) );
  INV_X1 U2244 ( .A(n553), .ZN(n555) );
  NOR2_X1 U2245 ( .A1(n983), .A2(n1002), .ZN(n563) );
  NAND2_X1 U2246 ( .A1(n983), .A2(n1002), .ZN(n564) );
  NAND3_X1 U2247 ( .A1(n2246), .A2(n2247), .A3(n2248), .ZN(n2230) );
  INV_X1 U2248 ( .A(n2348), .ZN(n2344) );
  XOR2_X1 U2249 ( .A(n1304), .B(n1282), .Z(n2232) );
  XOR2_X1 U2250 ( .A(n2232), .B(n1414), .Z(n955) );
  NAND2_X1 U2251 ( .A1(n1414), .A2(n1304), .ZN(n2233) );
  NAND2_X1 U2252 ( .A1(n1414), .A2(n1282), .ZN(n2234) );
  NAND2_X1 U2253 ( .A1(n1304), .A2(n1282), .ZN(n2235) );
  NAND3_X1 U2254 ( .A1(n2233), .A2(n2234), .A3(n2235), .ZN(n954) );
  XNOR2_X1 U2255 ( .A(b[17]), .B(n2344), .ZN(n1688) );
  OAI21_X1 U2256 ( .B1(n2094), .B2(n2017), .A(n2374), .ZN(n1242) );
  OAI21_X1 U2257 ( .B1(n2170), .B2(n2198), .A(n2371), .ZN(n1314) );
  OAI21_X1 U2258 ( .B1(n628), .B2(n626), .A(n627), .ZN(n625) );
  NOR2_X1 U2259 ( .A1(n1159), .A2(n1161), .ZN(n626) );
  AOI21_X1 U2260 ( .B1(n595), .B2(n609), .A(n596), .ZN(n594) );
  OAI21_X1 U2261 ( .B1(n558), .B2(n564), .A(n559), .ZN(n553) );
  NAND2_X1 U2262 ( .A1(n2203), .A2(n2126), .ZN(n456) );
  XNOR2_X1 U2263 ( .A(b[7]), .B(n2357), .ZN(n1748) );
  XNOR2_X1 U2264 ( .A(b[3]), .B(n2358), .ZN(n1752) );
  XNOR2_X1 U2265 ( .A(b[9]), .B(n2358), .ZN(n1746) );
  XNOR2_X1 U2266 ( .A(b[1]), .B(n2357), .ZN(n1754) );
  XNOR2_X1 U2267 ( .A(b[5]), .B(n2357), .ZN(n1750) );
  XNOR2_X1 U2268 ( .A(b[23]), .B(n2356), .ZN(n1732) );
  NOR2_X1 U2269 ( .A1(n839), .A2(n856), .ZN(n2236) );
  NOR2_X1 U2270 ( .A1(n839), .A2(n856), .ZN(n513) );
  INV_X1 U2271 ( .A(n2012), .ZN(n2321) );
  OAI21_X1 U2272 ( .B1(n2034), .B2(n1993), .A(n2368), .ZN(n1386) );
  NOR2_X1 U2273 ( .A1(n520), .A2(n513), .ZN(n511) );
  NOR2_X1 U2274 ( .A1(n857), .A2(n876), .ZN(n520) );
  NAND2_X1 U2275 ( .A1(n1000), .A2(n1393), .ZN(n2238) );
  NAND2_X1 U2276 ( .A1(n1000), .A2(n1415), .ZN(n2239) );
  NAND2_X1 U2277 ( .A1(n1393), .A2(n1415), .ZN(n2240) );
  NAND3_X1 U2278 ( .A1(n2238), .A2(n2239), .A3(n2240), .ZN(n974) );
  INV_X1 U2279 ( .A(n2094), .ZN(n2241) );
  OR2_X1 U2280 ( .A1(n2199), .A2(n1553), .ZN(n2242) );
  OR2_X1 U2281 ( .A1(n1552), .A2(n2287), .ZN(n2243) );
  NAND2_X1 U2282 ( .A1(n2242), .A2(n2243), .ZN(n1262) );
  XNOR2_X1 U2283 ( .A(n2096), .B(b[2]), .ZN(n1553) );
  XNOR2_X1 U2284 ( .A(b[3]), .B(n2096), .ZN(n1552) );
  OAI21_X1 U2285 ( .B1(n2027), .B2(n2018), .A(n2372), .ZN(n1290) );
  INV_X1 U2286 ( .A(n2312), .ZN(n2308) );
  XOR2_X1 U2287 ( .A(n1416), .B(n1328), .Z(n2245) );
  NAND2_X1 U2288 ( .A1(n1416), .A2(n1306), .ZN(n2246) );
  NAND2_X1 U2289 ( .A1(n1306), .A2(n1328), .ZN(n2247) );
  NAND2_X1 U2290 ( .A1(n1416), .A2(n1328), .ZN(n2248) );
  NAND3_X1 U2291 ( .A1(n2246), .A2(n2248), .A3(n2247), .ZN(n994) );
  XNOR2_X1 U2292 ( .A(n2323), .B(b[6]), .ZN(n1599) );
  XNOR2_X1 U2293 ( .A(b[7]), .B(n2322), .ZN(n1598) );
  OAI21_X1 U2294 ( .B1(n2164), .B2(n2049), .A(n2370), .ZN(n1338) );
  XOR2_X1 U2295 ( .A(n1083), .B(n1081), .Z(n2249) );
  XOR2_X1 U2296 ( .A(n2249), .B(n1079), .Z(n1075) );
  NAND2_X1 U2297 ( .A1(n1399), .A2(n1421), .ZN(n2250) );
  NAND2_X1 U2298 ( .A1(n1399), .A2(n1096), .ZN(n2251) );
  NAND2_X1 U2299 ( .A1(n1421), .A2(n1096), .ZN(n2252) );
  NAND3_X1 U2300 ( .A1(n2250), .A2(n2251), .A3(n2252), .ZN(n1078) );
  NAND2_X1 U2301 ( .A1(n1083), .A2(n1081), .ZN(n2253) );
  NAND2_X1 U2302 ( .A1(n1083), .A2(n1079), .ZN(n2254) );
  NAND2_X1 U2303 ( .A1(n1081), .A2(n1079), .ZN(n2255) );
  NAND3_X1 U2304 ( .A1(n2253), .A2(n2254), .A3(n2255), .ZN(n1074) );
  XNOR2_X1 U2305 ( .A(n486), .B(n315), .ZN(product[31]) );
  INV_X1 U2306 ( .A(n2316), .ZN(n2314) );
  OAI22_X1 U2307 ( .A1(n2179), .A2(n1636), .B1(n1986), .B2(n1635), .ZN(n1341)
         );
  OAI22_X1 U2308 ( .A1(n2179), .A2(n1634), .B1(n2295), .B2(n1633), .ZN(n1339)
         );
  OAI22_X1 U2309 ( .A1(n2180), .A2(n1640), .B1(n2295), .B2(n1639), .ZN(n1345)
         );
  OAI21_X1 U2310 ( .B1(n428), .B2(n436), .A(n429), .ZN(n427) );
  INV_X1 U2311 ( .A(n439), .ZN(n445) );
  NAND2_X1 U2312 ( .A1(n839), .A2(n856), .ZN(n514) );
  NOR2_X1 U2313 ( .A1(n389), .A2(n384), .ZN(n382) );
  OAI22_X1 U2314 ( .A1(n2040), .A2(n2362), .B1(n1781), .B2(n2304), .ZN(n1193)
         );
  OAI22_X1 U2315 ( .A1(n2041), .A2(n1767), .B1(n1766), .B2(n2304), .ZN(n1468)
         );
  OAI22_X1 U2316 ( .A1(n2040), .A2(n1760), .B1(n1759), .B2(n2304), .ZN(n1461)
         );
  OAI22_X1 U2317 ( .A1(n2281), .A2(n1764), .B1(n1763), .B2(n2304), .ZN(n1465)
         );
  OAI22_X1 U2318 ( .A1(n2041), .A2(n1759), .B1(n1758), .B2(n2303), .ZN(n1460)
         );
  OAI22_X1 U2319 ( .A1(n2281), .A2(n1763), .B1(n1762), .B2(n2304), .ZN(n1464)
         );
  OAI22_X1 U2320 ( .A1(n2282), .A2(n1761), .B1(n1760), .B2(n2303), .ZN(n1462)
         );
  OAI22_X1 U2321 ( .A1(n2282), .A2(n1762), .B1(n1761), .B2(n2303), .ZN(n1463)
         );
  OAI22_X1 U2322 ( .A1(n2040), .A2(n1765), .B1(n1764), .B2(n2304), .ZN(n1466)
         );
  OAI22_X1 U2323 ( .A1(n2281), .A2(n1766), .B1(n1765), .B2(n2304), .ZN(n1467)
         );
  OAI22_X1 U2324 ( .A1(n2041), .A2(n1768), .B1(n1767), .B2(n2304), .ZN(n1469)
         );
  OAI22_X1 U2325 ( .A1(n2282), .A2(n1758), .B1(n1757), .B2(n2303), .ZN(n1459)
         );
  XNOR2_X1 U2326 ( .A(b[1]), .B(n2028), .ZN(n1779) );
  XNOR2_X1 U2327 ( .A(b[5]), .B(n2029), .ZN(n1775) );
  XNOR2_X1 U2328 ( .A(b[9]), .B(n2360), .ZN(n1771) );
  XNOR2_X1 U2329 ( .A(b[3]), .B(n2028), .ZN(n1777) );
  XNOR2_X1 U2330 ( .A(b[7]), .B(n2360), .ZN(n1773) );
  XNOR2_X1 U2331 ( .A(b[23]), .B(n2361), .ZN(n1757) );
  NAND2_X1 U2332 ( .A1(n668), .A2(n503), .ZN(n317) );
  INV_X1 U2333 ( .A(n503), .ZN(n501) );
  INV_X1 U2334 ( .A(n2109), .ZN(n492) );
  INV_X1 U2335 ( .A(n2173), .ZN(n2274) );
  OAI22_X1 U2336 ( .A1(n2033), .A2(n1642), .B1(n2295), .B2(n1641), .ZN(n1347)
         );
  OAI22_X1 U2337 ( .A1(n1998), .A2(n1513), .B1(n2013), .B2(n1512), .ZN(n1223)
         );
  OAI22_X1 U2338 ( .A1(n1998), .A2(n1515), .B1(n2285), .B2(n1514), .ZN(n1225)
         );
  OAI22_X1 U2339 ( .A1(n1998), .A2(n1511), .B1(n2285), .B2(n1510), .ZN(n1221)
         );
  OAI22_X1 U2340 ( .A1(n1998), .A2(n1509), .B1(n2285), .B2(n1508), .ZN(n1219)
         );
  OAI22_X1 U2341 ( .A1(n1998), .A2(n1517), .B1(n2285), .B2(n1516), .ZN(n1227)
         );
  NOR2_X1 U2342 ( .A1(n2065), .A2(n467), .ZN(n465) );
  OAI21_X1 U2343 ( .B1(n492), .B2(n467), .A(n468), .ZN(n466) );
  OAI21_X1 U2344 ( .B1(n2162), .B2(n2023), .A(n2367), .ZN(n1410) );
  INV_X1 U2345 ( .A(n2157), .ZN(n2299) );
  NAND2_X1 U2346 ( .A1(n877), .A2(n896), .ZN(n532) );
  OAI21_X1 U2347 ( .B1(n2004), .B2(n2077), .A(n2366), .ZN(n1434) );
  OAI21_X1 U2348 ( .B1(n590), .B2(n593), .A(n591), .ZN(n589) );
  NOR2_X1 U2349 ( .A1(n590), .A2(n592), .ZN(n588) );
  OAI22_X1 U2350 ( .A1(n1939), .A2(n1593), .B1(n1592), .B2(n2291), .ZN(n1300)
         );
  OAI22_X1 U2351 ( .A1(n1931), .A2(n1584), .B1(n2291), .B2(n1583), .ZN(n1291)
         );
  OAI22_X1 U2352 ( .A1(n1931), .A2(n1589), .B1(n1588), .B2(n2290), .ZN(n1296)
         );
  OAI22_X1 U2353 ( .A1(n1931), .A2(n1590), .B1(n2291), .B2(n1589), .ZN(n1297)
         );
  OAI22_X1 U2354 ( .A1(n1931), .A2(n1588), .B1(n2290), .B2(n1587), .ZN(n1295)
         );
  OAI22_X1 U2355 ( .A1(n1931), .A2(n1583), .B1(n1582), .B2(n2290), .ZN(n724)
         );
  OAI22_X1 U2356 ( .A1(n1939), .A2(n1585), .B1(n1584), .B2(n2291), .ZN(n1292)
         );
  OAI22_X1 U2357 ( .A1(n1931), .A2(n1591), .B1(n1590), .B2(n2291), .ZN(n1298)
         );
  OAI22_X1 U2358 ( .A1(n1931), .A2(n1592), .B1(n2291), .B2(n1591), .ZN(n1299)
         );
  OAI22_X1 U2359 ( .A1(n1939), .A2(n1587), .B1(n1586), .B2(n2291), .ZN(n1294)
         );
  OAI22_X1 U2360 ( .A1(n1939), .A2(n1586), .B1(n2290), .B2(n1585), .ZN(n1293)
         );
  OAI22_X1 U2361 ( .A1(n1931), .A2(n2326), .B1(n1606), .B2(n2290), .ZN(n1186)
         );
  NAND2_X1 U2362 ( .A1(n956), .A2(n958), .ZN(n2258) );
  NAND2_X1 U2363 ( .A1(n956), .A2(n954), .ZN(n2259) );
  NAND2_X1 U2364 ( .A1(n958), .A2(n954), .ZN(n2260) );
  NAND3_X1 U2365 ( .A1(n2258), .A2(n2259), .A3(n2260), .ZN(n928) );
  AND2_X1 U2366 ( .A1(n2273), .A2(n2272), .ZN(n2265) );
  AND2_X1 U2367 ( .A1(n2273), .A2(n2272), .ZN(n301) );
  AOI21_X1 U2368 ( .B1(n629), .B2(n635), .A(n630), .ZN(n628) );
  AOI21_X1 U2369 ( .B1(n565), .B2(n2006), .A(n2098), .ZN(n551) );
  INV_X1 U2370 ( .A(n552), .ZN(n554) );
  INV_X1 U2371 ( .A(n2097), .ZN(n667) );
  INV_X1 U2372 ( .A(n2068), .ZN(n673) );
  OAI21_X1 U2373 ( .B1(n2087), .B2(n550), .A(n543), .ZN(n541) );
  NAND2_X1 U2374 ( .A1(n2128), .A2(n418), .ZN(n309) );
  OAI21_X1 U2375 ( .B1(n337), .B2(n334), .A(n335), .ZN(n333) );
  INV_X1 U2376 ( .A(n418), .ZN(n416) );
  AOI21_X1 U2377 ( .B1(n2126), .B2(n1938), .A(n459), .ZN(n457) );
  INV_X1 U2378 ( .A(n505), .ZN(n507) );
  OAI21_X1 U2379 ( .B1(n2161), .B2(n2231), .A(n2369), .ZN(n1362) );
  NAND2_X1 U2380 ( .A1(n2056), .A2(n2091), .ZN(n321) );
  NAND2_X1 U2381 ( .A1(n1085), .A2(n1098), .ZN(n593) );
  NOR2_X1 U2382 ( .A1(n1085), .A2(n1098), .ZN(n592) );
  NOR2_X1 U2383 ( .A1(n1165), .A2(n1170), .ZN(n631) );
  OAI21_X1 U2384 ( .B1(n631), .B2(n634), .A(n632), .ZN(n630) );
  NOR2_X1 U2385 ( .A1(n633), .A2(n631), .ZN(n629) );
  NOR2_X1 U2386 ( .A1(n456), .A2(n480), .ZN(n454) );
  XOR2_X1 U2387 ( .A(n1062), .B(n1053), .Z(n2261) );
  XOR2_X1 U2388 ( .A(n1060), .B(n2261), .Z(n1043) );
  NAND2_X1 U2389 ( .A1(n1060), .A2(n1062), .ZN(n2262) );
  NAND2_X1 U2390 ( .A1(n1060), .A2(n1053), .ZN(n2263) );
  NAND2_X1 U2391 ( .A1(n1062), .A2(n1053), .ZN(n2264) );
  NAND3_X1 U2392 ( .A1(n2262), .A2(n2263), .A3(n2264), .ZN(n1042) );
  XNOR2_X1 U2393 ( .A(n533), .B(n320), .ZN(product[26]) );
  NOR2_X1 U2394 ( .A1(n918), .A2(n897), .ZN(n534) );
  NAND2_X1 U2395 ( .A1(n897), .A2(n918), .ZN(n535) );
  XNOR2_X1 U2396 ( .A(b[17]), .B(n2308), .ZN(n1513) );
  NOR2_X1 U2397 ( .A1(n571), .A2(n1983), .ZN(n567) );
  NAND2_X1 U2398 ( .A1(n821), .A2(n838), .ZN(n503) );
  INV_X1 U2399 ( .A(n874), .ZN(n875) );
  INV_X1 U2400 ( .A(n2003), .ZN(n671) );
  INV_X1 U2401 ( .A(n2107), .ZN(n565) );
  INV_X1 U2402 ( .A(n400), .ZN(n398) );
  NAND2_X1 U2403 ( .A1(n400), .A2(n2132), .ZN(n389) );
  NOR2_X1 U2404 ( .A1(n420), .A2(n402), .ZN(n400) );
  OAI21_X1 U2405 ( .B1(n456), .B2(n481), .A(n457), .ZN(n455) );
  OAI21_X1 U2406 ( .B1(n2097), .B2(n503), .A(n496), .ZN(n490) );
  INV_X1 U2407 ( .A(n2042), .ZN(n508) );
  OAI21_X1 U2408 ( .B1(n2236), .B2(n521), .A(n514), .ZN(n512) );
  OAI21_X1 U2409 ( .B1(n572), .B2(n569), .A(n570), .ZN(n568) );
  INV_X1 U2410 ( .A(n547), .ZN(n674) );
  NOR2_X1 U2411 ( .A1(n554), .A2(n547), .ZN(n545) );
  OAI21_X1 U2412 ( .B1(n555), .B2(n547), .A(n550), .ZN(n546) );
  NOR2_X1 U2413 ( .A1(n542), .A2(n547), .ZN(n540) );
  OAI21_X1 U2414 ( .B1(n594), .B2(n582), .A(n583), .ZN(n581) );
  XNOR2_X1 U2415 ( .A(n475), .B(n314), .ZN(product[32]) );
  INV_X1 U2416 ( .A(n401), .ZN(n399) );
  INV_X1 U2417 ( .A(n383), .ZN(n381) );
  AOI21_X1 U2418 ( .B1(n383), .B2(n2129), .A(n376), .ZN(n372) );
  OAI22_X1 U2419 ( .A1(n1984), .A2(n1683), .B1(n1682), .B2(n2036), .ZN(n2266)
         );
  NAND2_X1 U2420 ( .A1(n1171), .A2(n1174), .ZN(n634) );
  NOR2_X1 U2421 ( .A1(n1171), .A2(n1174), .ZN(n633) );
  NAND2_X1 U2422 ( .A1(n1071), .A2(n1084), .ZN(n591) );
  XNOR2_X1 U2423 ( .A(b[21]), .B(n2052), .ZN(n1559) );
  XNOR2_X1 U2424 ( .A(b[15]), .B(n2052), .ZN(n1565) );
  XNOR2_X1 U2425 ( .A(b[19]), .B(n2052), .ZN(n1561) );
  XNOR2_X1 U2426 ( .A(b[11]), .B(n2052), .ZN(n1569) );
  XNOR2_X1 U2427 ( .A(b[17]), .B(n2052), .ZN(n1563) );
  XNOR2_X1 U2428 ( .A(b[13]), .B(n2052), .ZN(n1567) );
  NAND2_X1 U2429 ( .A1(n382), .A2(n2129), .ZN(n371) );
  NAND2_X1 U2430 ( .A1(n426), .A2(n663), .ZN(n420) );
  NAND2_X1 U2431 ( .A1(n465), .A2(n507), .ZN(n463) );
  NAND2_X1 U2432 ( .A1(n507), .A2(n2115), .ZN(n487) );
  NAND2_X1 U2433 ( .A1(n507), .A2(n668), .ZN(n498) );
  NAND2_X1 U2434 ( .A1(n478), .A2(n507), .ZN(n476) );
  INV_X1 U2435 ( .A(n345), .ZN(n343) );
  NAND2_X1 U2436 ( .A1(n345), .A2(n2142), .ZN(n336) );
  NAND2_X1 U2437 ( .A1(n709), .A2(n716), .ZN(n409) );
  INV_X1 U2438 ( .A(n746), .ZN(n747) );
  AOI21_X1 U2439 ( .B1(n1935), .B2(n465), .A(n466), .ZN(n464) );
  AOI21_X1 U2440 ( .B1(n1935), .B2(n668), .A(n501), .ZN(n499) );
  AOI21_X1 U2441 ( .B1(n508), .B2(n478), .A(n479), .ZN(n477) );
  AOI21_X1 U2442 ( .B1(n508), .B2(n2115), .A(n2109), .ZN(n488) );
  XNOR2_X1 U2443 ( .A(n462), .B(n313), .ZN(product[33]) );
  NAND2_X1 U2444 ( .A1(n805), .A2(n820), .ZN(n496) );
  NAND2_X1 U2445 ( .A1(n996), .A2(n2230), .ZN(n2267) );
  NAND2_X1 U2446 ( .A1(n996), .A2(n1217), .ZN(n2268) );
  NAND2_X1 U2447 ( .A1(n994), .A2(n1217), .ZN(n2269) );
  NAND3_X1 U2448 ( .A1(n2267), .A2(n2268), .A3(n2269), .ZN(n972) );
  OR2_X1 U2449 ( .A1(n2032), .A2(n1576), .ZN(n2270) );
  OR2_X1 U2450 ( .A1(n1575), .A2(n2057), .ZN(n2271) );
  NAND2_X1 U2451 ( .A1(n2270), .A2(n2271), .ZN(n1284) );
  NAND2_X1 U2452 ( .A1(n450), .A2(n537), .ZN(n2272) );
  INV_X1 U2453 ( .A(n451), .ZN(n2273) );
  NOR2_X1 U2454 ( .A1(n2283), .A2(n2364), .ZN(n1217) );
  XNOR2_X1 U2455 ( .A(n2317), .B(b[4]), .ZN(n1576) );
  XNOR2_X1 U2456 ( .A(b[5]), .B(n2052), .ZN(n1575) );
  NOR2_X1 U2457 ( .A1(n505), .A2(n452), .ZN(n450) );
  INV_X1 U2458 ( .A(n420), .ZN(n422) );
  NOR2_X1 U2459 ( .A1(n420), .A2(n347), .ZN(n345) );
  OAI21_X1 U2460 ( .B1(n421), .B2(n402), .A(n405), .ZN(n401) );
  OAI21_X1 U2461 ( .B1(n390), .B2(n384), .A(n387), .ZN(n383) );
  AOI21_X1 U2462 ( .B1(n401), .B2(n2132), .A(n394), .ZN(n390) );
  XNOR2_X1 U2463 ( .A(n437), .B(n311), .ZN(product[35]) );
  OAI22_X1 U2464 ( .A1(n2041), .A2(n1772), .B1(n1771), .B2(n2304), .ZN(n1473)
         );
  OAI22_X1 U2465 ( .A1(n2281), .A2(n1773), .B1(n1772), .B2(n2304), .ZN(n1474)
         );
  OAI22_X1 U2466 ( .A1(n2041), .A2(n1780), .B1(n1779), .B2(n2304), .ZN(n1481)
         );
  OAI22_X1 U2467 ( .A1(n2040), .A2(n1776), .B1(n1775), .B2(n2304), .ZN(n1477)
         );
  OAI22_X1 U2468 ( .A1(n2040), .A2(n1771), .B1(n1770), .B2(n2304), .ZN(n1472)
         );
  OAI22_X1 U2469 ( .A1(n2040), .A2(n1779), .B1(n1778), .B2(n2304), .ZN(n1480)
         );
  OAI22_X1 U2470 ( .A1(n2281), .A2(n1769), .B1(n1768), .B2(n2304), .ZN(n1470)
         );
  OAI22_X1 U2471 ( .A1(n2281), .A2(n1777), .B1(n1776), .B2(n2304), .ZN(n1478)
         );
  OAI22_X1 U2472 ( .A1(n2281), .A2(n1775), .B1(n1774), .B2(n2304), .ZN(n1476)
         );
  OAI22_X1 U2473 ( .A1(n2041), .A2(n1774), .B1(n1773), .B2(n2304), .ZN(n1475)
         );
  OAI22_X1 U2474 ( .A1(n2281), .A2(n1770), .B1(n1769), .B2(n2304), .ZN(n1471)
         );
  OAI22_X1 U2475 ( .A1(n2041), .A2(n1778), .B1(n1777), .B2(n2304), .ZN(n1479)
         );
  XNOR2_X1 U2476 ( .A(n430), .B(n310), .ZN(product[36]) );
  OAI22_X1 U2477 ( .A1(n2179), .A2(n1637), .B1(n1636), .B2(n1985), .ZN(n1342)
         );
  OAI22_X1 U2478 ( .A1(n2179), .A2(n1635), .B1(n1634), .B2(n1986), .ZN(n1340)
         );
  OAI22_X1 U2479 ( .A1(n2180), .A2(n1639), .B1(n1638), .B2(n1986), .ZN(n1344)
         );
  NAND2_X1 U2480 ( .A1(n1165), .A2(n1170), .ZN(n632) );
  XNOR2_X1 U2481 ( .A(n419), .B(n309), .ZN(product[37]) );
  NAND2_X1 U2482 ( .A1(n694), .A2(n689), .ZN(n378) );
  INV_X1 U2483 ( .A(n706), .ZN(n707) );
  OAI21_X1 U2484 ( .B1(n538), .B2(n566), .A(n539), .ZN(n537) );
  XNOR2_X1 U2485 ( .A(n410), .B(n308), .ZN(product[38]) );
  XNOR2_X1 U2486 ( .A(n397), .B(n307), .ZN(product[39]) );
  OAI22_X1 U2487 ( .A1(n2108), .A2(n1695), .B1(n1694), .B2(n2036), .ZN(n1398)
         );
  OAI22_X1 U2488 ( .A1(n2108), .A2(n1704), .B1(n2036), .B2(n1703), .ZN(n1407)
         );
  OAI22_X1 U2489 ( .A1(n2108), .A2(n1701), .B1(n1700), .B2(n2036), .ZN(n1404)
         );
  OAI22_X1 U2490 ( .A1(n1984), .A2(n1702), .B1(n2297), .B2(n1701), .ZN(n1405)
         );
  OAI22_X1 U2491 ( .A1(n2108), .A2(n1698), .B1(n2036), .B2(n1697), .ZN(n1401)
         );
  OAI22_X1 U2492 ( .A1(n2278), .A2(n1694), .B1(n2297), .B2(n1693), .ZN(n1397)
         );
  OAI22_X1 U2493 ( .A1(n2108), .A2(n1696), .B1(n2297), .B2(n1695), .ZN(n1399)
         );
  OAI22_X1 U2494 ( .A1(n2108), .A2(n1700), .B1(n2297), .B2(n1699), .ZN(n1403)
         );
  OAI22_X1 U2495 ( .A1(n2108), .A2(n1699), .B1(n1698), .B2(n2297), .ZN(n1402)
         );
  OAI22_X1 U2496 ( .A1(n2108), .A2(n1705), .B1(n1704), .B2(n2297), .ZN(n1408)
         );
  OAI22_X1 U2497 ( .A1(n2108), .A2(n1703), .B1(n1702), .B2(n2036), .ZN(n1406)
         );
  OAI22_X1 U2498 ( .A1(n1984), .A2(n1697), .B1(n1696), .B2(n2297), .ZN(n1400)
         );
  NOR2_X1 U2499 ( .A1(n402), .A2(n360), .ZN(n356) );
  NAND2_X1 U2500 ( .A1(n362), .A2(n2132), .ZN(n360) );
  NAND2_X1 U2501 ( .A1(n761), .A2(n774), .ZN(n461) );
  NAND2_X1 U2502 ( .A1(n663), .A2(n662), .ZN(n431) );
  XNOR2_X1 U2503 ( .A(b[11]), .B(n2339), .ZN(n1669) );
  XNOR2_X1 U2504 ( .A(b[17]), .B(n2339), .ZN(n1663) );
  XNOR2_X1 U2505 ( .A(b[19]), .B(n2339), .ZN(n1661) );
  XNOR2_X1 U2506 ( .A(b[15]), .B(n2339), .ZN(n1665) );
  XNOR2_X1 U2507 ( .A(b[21]), .B(n2339), .ZN(n1659) );
  XNOR2_X1 U2508 ( .A(b[13]), .B(n2339), .ZN(n1667) );
  OAI22_X1 U2509 ( .A1(n2010), .A2(n1613), .B1(n2015), .B2(n1612), .ZN(n1319)
         );
  OAI22_X1 U2510 ( .A1(n2059), .A2(n1612), .B1(n1611), .B2(n2015), .ZN(n1318)
         );
  OAI22_X1 U2511 ( .A1(n2059), .A2(n1617), .B1(n2292), .B2(n1616), .ZN(n1323)
         );
  OAI22_X1 U2512 ( .A1(n2010), .A2(n1610), .B1(n1609), .B2(n2015), .ZN(n1316)
         );
  OAI22_X1 U2513 ( .A1(n2059), .A2(n1609), .B1(n2016), .B2(n1608), .ZN(n1315)
         );
  OAI22_X1 U2514 ( .A1(n2059), .A2(n2331), .B1(n1631), .B2(n2014), .ZN(n1187)
         );
  OAI22_X1 U2515 ( .A1(n2059), .A2(n1611), .B1(n2292), .B2(n1610), .ZN(n1317)
         );
  OAI22_X1 U2516 ( .A1(n2010), .A2(n1615), .B1(n2015), .B2(n1614), .ZN(n1321)
         );
  OAI22_X1 U2517 ( .A1(n2010), .A2(n1618), .B1(n1617), .B2(n2014), .ZN(n1324)
         );
  OAI22_X1 U2518 ( .A1(n2081), .A2(n1614), .B1(n1613), .B2(n2292), .ZN(n1320)
         );
  XNOR2_X1 U2519 ( .A(b[19]), .B(n2005), .ZN(n1636) );
  OAI22_X1 U2520 ( .A1(n2081), .A2(n1616), .B1(n1615), .B2(n2292), .ZN(n1322)
         );
  XNOR2_X1 U2521 ( .A(b[21]), .B(n2334), .ZN(n1634) );
  XNOR2_X1 U2522 ( .A(b[11]), .B(n2334), .ZN(n1644) );
  XNOR2_X1 U2523 ( .A(b[17]), .B(n2334), .ZN(n1638) );
  XNOR2_X1 U2524 ( .A(b[15]), .B(n2334), .ZN(n1640) );
  XNOR2_X1 U2525 ( .A(b[13]), .B(n2334), .ZN(n1642) );
  XNOR2_X1 U2526 ( .A(n388), .B(n306), .ZN(product[40]) );
  OAI22_X1 U2527 ( .A1(n2275), .A2(n1570), .B1(n1569), .B2(n2057), .ZN(n1278)
         );
  OAI22_X1 U2528 ( .A1(n2275), .A2(n1571), .B1(n2289), .B2(n1570), .ZN(n1279)
         );
  OAI22_X1 U2529 ( .A1(n2275), .A2(n1575), .B1(n2057), .B2(n1574), .ZN(n1283)
         );
  OAI22_X1 U2530 ( .A1(n2275), .A2(n1580), .B1(n1579), .B2(n2289), .ZN(n1288)
         );
  OAI22_X1 U2531 ( .A1(n2275), .A2(n1579), .B1(n2057), .B2(n1578), .ZN(n1287)
         );
  OAI22_X1 U2532 ( .A1(n2275), .A2(n1578), .B1(n1577), .B2(n2289), .ZN(n1286)
         );
  OAI22_X1 U2533 ( .A1(n2275), .A2(n1573), .B1(n2057), .B2(n1572), .ZN(n1281)
         );
  OAI22_X1 U2534 ( .A1(n2274), .A2(n1569), .B1(n2057), .B2(n1568), .ZN(n1277)
         );
  OAI22_X1 U2535 ( .A1(n2274), .A2(n1577), .B1(n2057), .B2(n1576), .ZN(n1285)
         );
  OAI22_X1 U2536 ( .A1(n1572), .A2(n2274), .B1(n1571), .B2(n2289), .ZN(n1280)
         );
  OAI22_X1 U2537 ( .A1(n2274), .A2(n1574), .B1(n1573), .B2(n2057), .ZN(n1282)
         );
  OAI22_X1 U2538 ( .A1(n1998), .A2(n1508), .B1(n1507), .B2(n2013), .ZN(n682)
         );
  OAI22_X1 U2539 ( .A1(n1998), .A2(n1518), .B1(n1517), .B2(n2286), .ZN(n1228)
         );
  OAI22_X1 U2540 ( .A1(n1998), .A2(n1514), .B1(n1513), .B2(n2286), .ZN(n1224)
         );
  XNOR2_X1 U2541 ( .A(b[19]), .B(n2314), .ZN(n1536) );
  OAI22_X1 U2542 ( .A1(n1998), .A2(n1510), .B1(n1509), .B2(n2286), .ZN(n1220)
         );
  OAI22_X1 U2543 ( .A1(n1998), .A2(n1516), .B1(n1515), .B2(n2285), .ZN(n1226)
         );
  XNOR2_X1 U2544 ( .A(b[21]), .B(n2314), .ZN(n1534) );
  OAI22_X1 U2545 ( .A1(n1998), .A2(n2037), .B1(n1531), .B2(n2286), .ZN(n1183)
         );
  OAI22_X1 U2546 ( .A1(n1998), .A2(n1512), .B1(n1511), .B2(n2286), .ZN(n1222)
         );
  XNOR2_X1 U2547 ( .A(b[17]), .B(n2314), .ZN(n1538) );
  XNOR2_X1 U2548 ( .A(b[13]), .B(n2314), .ZN(n1542) );
  XNOR2_X1 U2549 ( .A(b[15]), .B(n2314), .ZN(n1540) );
  XNOR2_X1 U2550 ( .A(b[11]), .B(n2314), .ZN(n1544) );
  OAI22_X1 U2551 ( .A1(n2177), .A2(n2354), .B1(n1731), .B2(n2300), .ZN(n1191)
         );
  OAI22_X1 U2552 ( .A1(n2177), .A2(n1718), .B1(n1717), .B2(n2299), .ZN(n1420)
         );
  OAI22_X1 U2553 ( .A1(n2279), .A2(n1716), .B1(n1715), .B2(n2300), .ZN(n1418)
         );
  OAI22_X1 U2554 ( .A1(n2280), .A2(n1715), .B1(n2300), .B2(n1714), .ZN(n1417)
         );
  OAI22_X1 U2555 ( .A1(n1932), .A2(n1713), .B1(n2300), .B2(n1712), .ZN(n1415)
         );
  OAI22_X1 U2556 ( .A1(n1932), .A2(n1717), .B1(n2300), .B2(n1716), .ZN(n1419)
         );
  OAI22_X1 U2557 ( .A1(n1932), .A2(n1708), .B1(n1707), .B2(n2299), .ZN(n874)
         );
  OAI22_X1 U2558 ( .A1(n2279), .A2(n1711), .B1(n2299), .B2(n1710), .ZN(n1413)
         );
  OAI22_X1 U2559 ( .A1(n2279), .A2(n1709), .B1(n2299), .B2(n1708), .ZN(n1411)
         );
  OAI22_X1 U2560 ( .A1(n2031), .A2(n1710), .B1(n1709), .B2(n2299), .ZN(n1412)
         );
  OAI22_X1 U2561 ( .A1(n1932), .A2(n1712), .B1(n1711), .B2(n2299), .ZN(n1414)
         );
  OAI22_X1 U2562 ( .A1(n2279), .A2(n1714), .B1(n1713), .B2(n2300), .ZN(n1416)
         );
  INV_X1 U2563 ( .A(n2266), .ZN(n837) );
  XNOR2_X1 U2564 ( .A(b[17]), .B(n2360), .ZN(n1763) );
  XNOR2_X1 U2565 ( .A(b[21]), .B(n2029), .ZN(n1759) );
  XNOR2_X1 U2566 ( .A(b[13]), .B(n2360), .ZN(n1767) );
  XNOR2_X1 U2567 ( .A(b[19]), .B(n2361), .ZN(n1761) );
  XNOR2_X1 U2568 ( .A(b[15]), .B(n2360), .ZN(n1765) );
  XNOR2_X1 U2569 ( .A(b[11]), .B(n2360), .ZN(n1769) );
  OAI22_X1 U2570 ( .A1(n2179), .A2(n1652), .B1(n2295), .B2(n1651), .ZN(n1357)
         );
  OAI22_X1 U2571 ( .A1(n2179), .A2(n1645), .B1(n1644), .B2(n1986), .ZN(n1350)
         );
  OAI22_X1 U2572 ( .A1(n2179), .A2(n1649), .B1(n1648), .B2(n1986), .ZN(n1354)
         );
  OAI22_X1 U2573 ( .A1(n2179), .A2(n1653), .B1(n1652), .B2(n2295), .ZN(n1358)
         );
  OAI22_X1 U2574 ( .A1(n2180), .A2(n1648), .B1(n1985), .B2(n1647), .ZN(n1353)
         );
  OAI22_X1 U2575 ( .A1(n2033), .A2(n1644), .B1(n1985), .B2(n1643), .ZN(n1349)
         );
  OAI22_X1 U2576 ( .A1(n2179), .A2(n1654), .B1(n1985), .B2(n1653), .ZN(n1359)
         );
  OAI22_X1 U2577 ( .A1(n2179), .A2(n1655), .B1(n1654), .B2(n1985), .ZN(n1360)
         );
  OAI22_X1 U2578 ( .A1(n2180), .A2(n1647), .B1(n1646), .B2(n2295), .ZN(n1352)
         );
  OAI22_X1 U2579 ( .A1(n2180), .A2(n1651), .B1(n1650), .B2(n2295), .ZN(n1356)
         );
  OAI22_X1 U2580 ( .A1(n2180), .A2(n1650), .B1(n2295), .B2(n1649), .ZN(n1355)
         );
  INV_X1 U2581 ( .A(n421), .ZN(n423) );
  OAI21_X1 U2582 ( .B1(n421), .B2(n347), .A(n348), .ZN(n346) );
  INV_X1 U2583 ( .A(n772), .ZN(n773) );
  OAI22_X1 U2584 ( .A1(n1936), .A2(n1535), .B1(n1534), .B2(n2287), .ZN(n1244)
         );
  OAI22_X1 U2585 ( .A1(n2241), .A2(n1537), .B1(n1536), .B2(n2288), .ZN(n1246)
         );
  OAI22_X1 U2586 ( .A1(n1936), .A2(n1544), .B1(n2288), .B2(n1543), .ZN(n1253)
         );
  OAI22_X1 U2587 ( .A1(n2241), .A2(n2316), .B1(n1556), .B2(n2288), .ZN(n1184)
         );
  OAI22_X1 U2588 ( .A1(n1936), .A2(n1539), .B1(n1538), .B2(n2287), .ZN(n1248)
         );
  OAI22_X1 U2589 ( .A1(n1936), .A2(n1543), .B1(n1542), .B2(n2288), .ZN(n1252)
         );
  OAI22_X1 U2590 ( .A1(n1936), .A2(n1552), .B1(n2288), .B2(n1551), .ZN(n1261)
         );
  OAI22_X1 U2591 ( .A1(n1936), .A2(n1555), .B1(n1554), .B2(n2288), .ZN(n1264)
         );
  OAI22_X1 U2592 ( .A1(n1936), .A2(n1546), .B1(n2288), .B2(n1545), .ZN(n1255)
         );
  OAI22_X1 U2593 ( .A1(n1936), .A2(n1549), .B1(n1548), .B2(n2288), .ZN(n1258)
         );
  OAI22_X1 U2594 ( .A1(n2199), .A2(n1548), .B1(n2288), .B2(n1547), .ZN(n1257)
         );
  OAI22_X1 U2595 ( .A1(n1936), .A2(n1533), .B1(n1532), .B2(n2287), .ZN(n692)
         );
  OAI22_X1 U2596 ( .A1(n2199), .A2(n1547), .B1(n1546), .B2(n2287), .ZN(n1256)
         );
  OAI22_X1 U2597 ( .A1(n2241), .A2(n1541), .B1(n1540), .B2(n2288), .ZN(n1250)
         );
  OAI22_X1 U2598 ( .A1(n2199), .A2(n1545), .B1(n1544), .B2(n2288), .ZN(n1254)
         );
  OAI22_X1 U2599 ( .A1(n2199), .A2(n1554), .B1(n2287), .B2(n1553), .ZN(n1263)
         );
  OAI22_X1 U2600 ( .A1(n2199), .A2(n1551), .B1(n1550), .B2(n2287), .ZN(n1260)
         );
  XNOR2_X1 U2601 ( .A(b[13]), .B(n2344), .ZN(n1692) );
  XNOR2_X1 U2602 ( .A(b[11]), .B(n2344), .ZN(n1694) );
  XNOR2_X1 U2603 ( .A(b[21]), .B(n2344), .ZN(n1684) );
  XNOR2_X1 U2604 ( .A(b[19]), .B(n2344), .ZN(n1686) );
  XNOR2_X1 U2605 ( .A(b[15]), .B(n2344), .ZN(n1690) );
  OAI22_X1 U2606 ( .A1(n2047), .A2(n1747), .B1(n1746), .B2(n2301), .ZN(n1448)
         );
  OAI22_X1 U2607 ( .A1(n2048), .A2(n1749), .B1(n1748), .B2(n2301), .ZN(n1450)
         );
  OAI22_X1 U2608 ( .A1(n2047), .A2(n1748), .B1(n2301), .B2(n1747), .ZN(n1449)
         );
  OAI22_X1 U2609 ( .A1(n2048), .A2(n1744), .B1(n2301), .B2(n1743), .ZN(n1445)
         );
  OAI22_X1 U2610 ( .A1(n2046), .A2(n1753), .B1(n1752), .B2(n2301), .ZN(n1454)
         );
  OAI22_X1 U2611 ( .A1(n2048), .A2(n1750), .B1(n2301), .B2(n1749), .ZN(n1451)
         );
  OAI22_X1 U2612 ( .A1(n2047), .A2(n1745), .B1(n1744), .B2(n2301), .ZN(n1446)
         );
  XNOR2_X1 U2613 ( .A(b[15]), .B(n2308), .ZN(n1515) );
  XNOR2_X1 U2614 ( .A(b[19]), .B(n2308), .ZN(n1511) );
  XNOR2_X1 U2615 ( .A(b[13]), .B(n2308), .ZN(n1517) );
  XNOR2_X1 U2616 ( .A(b[21]), .B(n2308), .ZN(n1509) );
  XNOR2_X1 U2617 ( .A(b[11]), .B(n2308), .ZN(n1519) );
  OAI22_X1 U2618 ( .A1(n2059), .A2(n1623), .B1(n2016), .B2(n1622), .ZN(n1329)
         );
  OAI22_X1 U2619 ( .A1(n2059), .A2(n1626), .B1(n1625), .B2(n2015), .ZN(n1332)
         );
  OAI22_X1 U2620 ( .A1(n2010), .A2(n1630), .B1(n1629), .B2(n2024), .ZN(n1336)
         );
  OAI22_X1 U2621 ( .A1(n2010), .A2(n1620), .B1(n1619), .B2(n2016), .ZN(n1326)
         );
  OAI22_X1 U2622 ( .A1(n2010), .A2(n1625), .B1(n2016), .B2(n1624), .ZN(n1331)
         );
  OAI22_X1 U2623 ( .A1(n2010), .A2(n1621), .B1(n2015), .B2(n1620), .ZN(n1327)
         );
  OAI22_X1 U2624 ( .A1(n2059), .A2(n1629), .B1(n2016), .B2(n1628), .ZN(n1335)
         );
  OAI22_X1 U2625 ( .A1(n2048), .A2(n1755), .B1(n1754), .B2(n2301), .ZN(n1456)
         );
  OAI22_X1 U2626 ( .A1(n2048), .A2(n1751), .B1(n1750), .B2(n2301), .ZN(n1452)
         );
  OAI22_X1 U2627 ( .A1(n2047), .A2(n1752), .B1(n2301), .B2(n1751), .ZN(n1453)
         );
  OAI22_X1 U2628 ( .A1(n2047), .A2(n1754), .B1(n2301), .B2(n1753), .ZN(n1455)
         );
  OAI22_X1 U2629 ( .A1(n2048), .A2(n1746), .B1(n2301), .B2(n1745), .ZN(n1447)
         );
  OAI22_X1 U2630 ( .A1(n2176), .A2(n1669), .B1(n2296), .B2(n1668), .ZN(n1373)
         );
  OAI22_X1 U2631 ( .A1(n2176), .A2(n1670), .B1(n1669), .B2(n2296), .ZN(n1374)
         );
  OAI22_X1 U2632 ( .A1(n2176), .A2(n1671), .B1(n2296), .B2(n1670), .ZN(n1375)
         );
  OAI22_X1 U2633 ( .A1(n2175), .A2(n1672), .B1(n1671), .B2(n2296), .ZN(n1376)
         );
  OAI22_X1 U2634 ( .A1(n2276), .A2(n1679), .B1(n2296), .B2(n1678), .ZN(n1383)
         );
  OAI22_X1 U2635 ( .A1(n2276), .A2(n1677), .B1(n2296), .B2(n1676), .ZN(n1381)
         );
  OAI22_X1 U2636 ( .A1(n2176), .A2(n1675), .B1(n2296), .B2(n1674), .ZN(n1379)
         );
  OAI22_X1 U2637 ( .A1(n2175), .A2(n1676), .B1(n1675), .B2(n2296), .ZN(n1380)
         );
  OAI22_X1 U2638 ( .A1(n2276), .A2(n1680), .B1(n1679), .B2(n2178), .ZN(n1384)
         );
  OAI22_X1 U2639 ( .A1(n2276), .A2(n1674), .B1(n1673), .B2(n2296), .ZN(n1378)
         );
  OAI22_X1 U2640 ( .A1(n2175), .A2(n1673), .B1(n2296), .B2(n1672), .ZN(n1377)
         );
  OAI22_X1 U2641 ( .A1(n2175), .A2(n1678), .B1(n1677), .B2(n2178), .ZN(n1382)
         );
  NAND2_X1 U2642 ( .A1(n332), .A2(n2143), .ZN(n326) );
  AOI21_X1 U2643 ( .B1(n333), .B2(n2143), .A(n2144), .ZN(n327) );
  NAND2_X1 U2644 ( .A1(n356), .A2(n2141), .ZN(n347) );
  OAI22_X1 U2645 ( .A1(n2010), .A2(n1608), .B1(n1607), .B2(n2016), .ZN(n746)
         );
  AOI21_X1 U2646 ( .B1(n490), .B2(n454), .A(n455), .ZN(n453) );
  XNOR2_X1 U2647 ( .A(n379), .B(n305), .ZN(product[41]) );
  NAND2_X1 U2648 ( .A1(n454), .A2(n489), .ZN(n452) );
  NAND2_X1 U2649 ( .A1(n525), .A2(n511), .ZN(n505) );
  OAI22_X1 U2650 ( .A1(n2081), .A2(n1628), .B1(n1627), .B2(n2292), .ZN(n1334)
         );
  OAI22_X1 U2651 ( .A1(n2059), .A2(n1622), .B1(n1621), .B2(n2292), .ZN(n1328)
         );
  OAI22_X1 U2652 ( .A1(n2010), .A2(n1627), .B1(n2292), .B2(n1626), .ZN(n1333)
         );
  OAI22_X1 U2653 ( .A1(n2010), .A2(n1619), .B1(n2292), .B2(n1618), .ZN(n1325)
         );
  OAI22_X1 U2654 ( .A1(n2081), .A2(n1624), .B1(n1623), .B2(n2292), .ZN(n1330)
         );
  INV_X1 U2655 ( .A(n346), .ZN(n344) );
  AOI21_X1 U2656 ( .B1(n346), .B2(n2142), .A(n339), .ZN(n337) );
  OAI22_X1 U2657 ( .A1(n1940), .A2(n1483), .B1(n1482), .B2(n2000), .ZN(n676)
         );
  OAI22_X1 U2658 ( .A1(n1941), .A2(n1484), .B1(n2284), .B2(n1483), .ZN(n1195)
         );
  NAND2_X1 U2659 ( .A1(n717), .A2(n726), .ZN(n418) );
  OAI22_X1 U2660 ( .A1(n1940), .A2(n1485), .B1(n1484), .B2(n2000), .ZN(n1196)
         );
  OAI22_X1 U2661 ( .A1(n1941), .A2(n1491), .B1(n1490), .B2(n2000), .ZN(n1202)
         );
  OAI22_X1 U2662 ( .A1(n1940), .A2(n1486), .B1(n2284), .B2(n1485), .ZN(n1197)
         );
  OAI22_X1 U2663 ( .A1(n1941), .A2(n1488), .B1(n2284), .B2(n1487), .ZN(n1199)
         );
  OAI22_X1 U2664 ( .A1(n1940), .A2(n1487), .B1(n1486), .B2(n2000), .ZN(n1198)
         );
  OAI22_X1 U2665 ( .A1(n1941), .A2(n1492), .B1(n2284), .B2(n1491), .ZN(n1203)
         );
  OAI22_X1 U2666 ( .A1(n1941), .A2(n1490), .B1(n2284), .B2(n1489), .ZN(n1201)
         );
  OAI22_X1 U2667 ( .A1(n2070), .A2(n2307), .B1(n1506), .B2(n2284), .ZN(n1182)
         );
  OAI22_X1 U2668 ( .A1(n1940), .A2(n1493), .B1(n1492), .B2(n2284), .ZN(n1204)
         );
  OAI22_X1 U2669 ( .A1(n1940), .A2(n1489), .B1(n1488), .B2(n2283), .ZN(n1200)
         );
  XNOR2_X1 U2670 ( .A(n1237), .B(n1215), .ZN(n939) );
  OAI21_X1 U2671 ( .B1(n506), .B2(n452), .A(n453), .ZN(n451) );
  XNOR2_X1 U2672 ( .A(n370), .B(n304), .ZN(product[42]) );
  OAI22_X1 U2673 ( .A1(n2205), .A2(n1497), .B1(n1496), .B2(n2284), .ZN(n1208)
         );
  OAI22_X1 U2674 ( .A1(n1941), .A2(n1496), .B1(n2283), .B2(n1495), .ZN(n1207)
         );
  OAI22_X1 U2675 ( .A1(n2205), .A2(n1495), .B1(n1494), .B2(n2283), .ZN(n1206)
         );
  OAI22_X1 U2676 ( .A1(n2204), .A2(n1954), .B1(n2283), .B2(n1501), .ZN(n1213)
         );
  OAI22_X1 U2677 ( .A1(n2204), .A2(n1501), .B1(n1500), .B2(n2283), .ZN(n1212)
         );
  OAI22_X1 U2678 ( .A1(n1940), .A2(n1494), .B1(n2284), .B2(n1493), .ZN(n1205)
         );
  OAI22_X1 U2679 ( .A1(n2205), .A2(n1500), .B1(n2284), .B2(n1499), .ZN(n1211)
         );
  OAI22_X1 U2680 ( .A1(n2070), .A2(n1504), .B1(n2284), .B2(n1503), .ZN(n1215)
         );
  OAI22_X1 U2681 ( .A1(n2070), .A2(n1503), .B1(n1502), .B2(n2283), .ZN(n1214)
         );
  OAI22_X1 U2682 ( .A1(n2205), .A2(n1498), .B1(n2284), .B2(n1497), .ZN(n1209)
         );
  OAI22_X1 U2683 ( .A1(n1941), .A2(n1499), .B1(n1498), .B2(n2283), .ZN(n1210)
         );
  OAI22_X1 U2684 ( .A1(n2337), .A2(n2033), .B1(n1656), .B2(n2295), .ZN(n1188)
         );
  OAI22_X1 U2685 ( .A1(n2033), .A2(n1641), .B1(n1640), .B2(n1985), .ZN(n1346)
         );
  OAI22_X1 U2686 ( .A1(n2033), .A2(n1643), .B1(n1642), .B2(n2295), .ZN(n1348)
         );
  OAI22_X1 U2687 ( .A1(n2180), .A2(n1633), .B1(n1632), .B2(n1986), .ZN(n772)
         );
  OAI22_X1 U2688 ( .A1(n2180), .A2(n1638), .B1(n2295), .B2(n1637), .ZN(n1343)
         );
  XNOR2_X1 U2689 ( .A(n353), .B(n303), .ZN(product[43]) );
  OAI22_X1 U2690 ( .A1(n2175), .A2(n1661), .B1(n2296), .B2(n1660), .ZN(n1365)
         );
  OAI22_X1 U2691 ( .A1(n2175), .A2(n1660), .B1(n1659), .B2(n2178), .ZN(n1364)
         );
  OAI22_X1 U2692 ( .A1(n2175), .A2(n2342), .B1(n1681), .B2(n2178), .ZN(n1189)
         );
  OAI22_X1 U2693 ( .A1(n2175), .A2(n1663), .B1(n2296), .B2(n1662), .ZN(n1367)
         );
  OAI22_X1 U2694 ( .A1(n2176), .A2(n1667), .B1(n2296), .B2(n1666), .ZN(n1371)
         );
  OAI22_X1 U2695 ( .A1(n2176), .A2(n1664), .B1(n1663), .B2(n2178), .ZN(n1368)
         );
  OAI22_X1 U2696 ( .A1(n2175), .A2(n1665), .B1(n2296), .B2(n1664), .ZN(n1369)
         );
  OAI22_X1 U2697 ( .A1(n2176), .A2(n1662), .B1(n1661), .B2(n2178), .ZN(n1366)
         );
  OAI22_X1 U2698 ( .A1(n2176), .A2(n1658), .B1(n1657), .B2(n2178), .ZN(n802)
         );
  OAI22_X1 U2699 ( .A1(n2276), .A2(n1666), .B1(n1665), .B2(n2178), .ZN(n1370)
         );
  OAI22_X1 U2700 ( .A1(n2276), .A2(n1659), .B1(n2296), .B2(n1658), .ZN(n1363)
         );
  OAI22_X1 U2701 ( .A1(n2276), .A2(n1668), .B1(n1667), .B2(n2178), .ZN(n1372)
         );
  NAND2_X1 U2702 ( .A1(n1937), .A2(n552), .ZN(n538) );
  AOI21_X1 U2703 ( .B1(n553), .B2(n540), .A(n541), .ZN(n539) );
  OAI22_X1 U2704 ( .A1(n2070), .A2(n1505), .B1(n1504), .B2(n2283), .ZN(n1216)
         );
  XNOR2_X1 U2705 ( .A(n342), .B(n302), .ZN(product[44]) );
  OAI22_X1 U2706 ( .A1(n2047), .A2(n2359), .B1(n1756), .B2(n2301), .ZN(n1192)
         );
  OAI22_X1 U2707 ( .A1(n2047), .A2(n1738), .B1(n2301), .B2(n1737), .ZN(n1439)
         );
  OAI22_X1 U2708 ( .A1(n2048), .A2(n1741), .B1(n1740), .B2(n2301), .ZN(n1442)
         );
  OAI22_X1 U2709 ( .A1(n2047), .A2(n1740), .B1(n2301), .B2(n1739), .ZN(n1441)
         );
  OAI22_X1 U2710 ( .A1(n2046), .A2(n1735), .B1(n1734), .B2(n2301), .ZN(n1436)
         );
  OAI22_X1 U2711 ( .A1(n2046), .A2(n1739), .B1(n1738), .B2(n2302), .ZN(n1440)
         );
  INV_X1 U2712 ( .A(n916), .ZN(n917) );
  OAI22_X1 U2713 ( .A1(n2047), .A2(n1736), .B1(n2302), .B2(n1735), .ZN(n1437)
         );
  OAI22_X1 U2714 ( .A1(n2047), .A2(n1734), .B1(n2301), .B2(n1733), .ZN(n1435)
         );
  OAI22_X1 U2715 ( .A1(n2046), .A2(n1743), .B1(n1742), .B2(n2301), .ZN(n1444)
         );
  OAI22_X1 U2716 ( .A1(n1970), .A2(n1737), .B1(n1736), .B2(n2302), .ZN(n1438)
         );
  OAI22_X1 U2717 ( .A1(n1998), .A2(n1522), .B1(n1521), .B2(n2286), .ZN(n1232)
         );
  OAI22_X1 U2718 ( .A1(n1998), .A2(n1521), .B1(n2285), .B2(n1520), .ZN(n1231)
         );
  OAI22_X1 U2719 ( .A1(n1998), .A2(n1519), .B1(n2285), .B2(n1518), .ZN(n1229)
         );
  OAI22_X1 U2720 ( .A1(n1998), .A2(n1520), .B1(n1519), .B2(n2286), .ZN(n1230)
         );
  OAI22_X1 U2721 ( .A1(n1998), .A2(n1525), .B1(n2285), .B2(n1524), .ZN(n1235)
         );
  OAI22_X1 U2722 ( .A1(n2089), .A2(n1524), .B1(n1523), .B2(n2286), .ZN(n1234)
         );
  OAI22_X1 U2723 ( .A1(n1998), .A2(n1523), .B1(n2285), .B2(n1522), .ZN(n1233)
         );
  OAI22_X1 U2724 ( .A1(n1943), .A2(n1529), .B1(n2285), .B2(n1997), .ZN(n1239)
         );
  OAI22_X1 U2725 ( .A1(n2089), .A2(n1526), .B1(n1525), .B2(n2285), .ZN(n1236)
         );
  OAI22_X1 U2726 ( .A1(n1943), .A2(n1530), .B1(n1529), .B2(n2285), .ZN(n1240)
         );
  OAI22_X1 U2727 ( .A1(n2089), .A2(n1527), .B1(n2286), .B2(n1526), .ZN(n1237)
         );
  OAI22_X1 U2728 ( .A1(n1939), .A2(n1602), .B1(n2290), .B2(n1601), .ZN(n1309)
         );
  OAI22_X1 U2729 ( .A1(n1931), .A2(n1600), .B1(n2291), .B2(n1599), .ZN(n1307)
         );
  OAI22_X1 U2730 ( .A1(n1939), .A2(n1601), .B1(n1600), .B2(n2291), .ZN(n1308)
         );
  OAI22_X1 U2731 ( .A1(n1931), .A2(n1594), .B1(n2290), .B2(n1593), .ZN(n1301)
         );
  OAI22_X1 U2732 ( .A1(n1939), .A2(n1596), .B1(n2290), .B2(n1595), .ZN(n1303)
         );
  OAI22_X1 U2733 ( .A1(n1931), .A2(n1598), .B1(n2291), .B2(n1597), .ZN(n1305)
         );
  OAI22_X1 U2734 ( .A1(n1931), .A2(n1603), .B1(n1602), .B2(n2291), .ZN(n1310)
         );
  OAI22_X1 U2735 ( .A1(n1931), .A2(n1597), .B1(n1596), .B2(n2290), .ZN(n1304)
         );
  OAI22_X1 U2736 ( .A1(n1939), .A2(n1604), .B1(n2290), .B2(n1603), .ZN(n1311)
         );
  OAI22_X1 U2737 ( .A1(n1939), .A2(n1595), .B1(n1594), .B2(n2291), .ZN(n1302)
         );
  OAI22_X1 U2738 ( .A1(n1939), .A2(n1605), .B1(n1604), .B2(n2290), .ZN(n1312)
         );
  XNOR2_X1 U2739 ( .A(b[19]), .B(n2044), .ZN(n1611) );
  XNOR2_X1 U2740 ( .A(b[21]), .B(n2330), .ZN(n1609) );
  XNOR2_X1 U2741 ( .A(b[11]), .B(n2329), .ZN(n1619) );
  XNOR2_X1 U2742 ( .A(b[13]), .B(n2044), .ZN(n1617) );
  XNOR2_X1 U2743 ( .A(b[15]), .B(n2044), .ZN(n1615) );
  XNOR2_X1 U2744 ( .A(b[17]), .B(n2328), .ZN(n1613) );
  XOR2_X1 U2745 ( .A(n1988), .B(n321), .Z(product[25]) );
  OAI21_X1 U2746 ( .B1(n1989), .B2(n1999), .A(n2056), .ZN(n533) );
  OAI21_X1 U2747 ( .B1(n1988), .B2(n487), .A(n488), .ZN(n486) );
  OAI21_X1 U2748 ( .B1(n1988), .B2(n463), .A(n464), .ZN(n462) );
  OAI21_X1 U2749 ( .B1(n1987), .B2(n2090), .A(n524), .ZN(n522) );
  OAI21_X1 U2750 ( .B1(n1987), .B2(n476), .A(n477), .ZN(n475) );
  OAI21_X1 U2751 ( .B1(n1989), .B2(n516), .A(n517), .ZN(n515) );
  OAI21_X1 U2752 ( .B1(n1987), .B2(n2064), .A(n1990), .ZN(n504) );
  OAI21_X1 U2753 ( .B1(n1989), .B2(n498), .A(n499), .ZN(n497) );
  OAI22_X1 U2754 ( .A1(n2177), .A2(n1727), .B1(n2299), .B2(n1726), .ZN(n1429)
         );
  OAI22_X1 U2755 ( .A1(n2177), .A2(n1720), .B1(n1719), .B2(n2299), .ZN(n1422)
         );
  OAI22_X1 U2756 ( .A1(n2177), .A2(n1721), .B1(n2300), .B2(n1720), .ZN(n1423)
         );
  OAI22_X1 U2757 ( .A1(n2177), .A2(n1726), .B1(n1725), .B2(n2299), .ZN(n1428)
         );
  OAI22_X1 U2758 ( .A1(n2177), .A2(n1730), .B1(n1729), .B2(n2300), .ZN(n1432)
         );
  OAI22_X1 U2759 ( .A1(n2177), .A2(n1725), .B1(n2299), .B2(n1724), .ZN(n1427)
         );
  OAI22_X1 U2760 ( .A1(n2177), .A2(n1723), .B1(n2300), .B2(n1722), .ZN(n1425)
         );
  OAI22_X1 U2761 ( .A1(n2177), .A2(n1728), .B1(n1727), .B2(n2299), .ZN(n1430)
         );
  OAI22_X1 U2762 ( .A1(n2280), .A2(n1722), .B1(n1721), .B2(n2299), .ZN(n1424)
         );
  OAI22_X1 U2763 ( .A1(n2177), .A2(n1729), .B1(n2300), .B2(n1728), .ZN(n1431)
         );
  OAI22_X1 U2764 ( .A1(n2280), .A2(n1719), .B1(n2300), .B2(n1718), .ZN(n1421)
         );
  OAI22_X1 U2765 ( .A1(n2280), .A2(n1724), .B1(n1723), .B2(n2299), .ZN(n1426)
         );
  XNOR2_X1 U2766 ( .A(b[15]), .B(n2357), .ZN(n1740) );
  XNOR2_X1 U2767 ( .A(b[21]), .B(n2358), .ZN(n1734) );
  XNOR2_X1 U2768 ( .A(b[19]), .B(n2357), .ZN(n1736) );
  XNOR2_X1 U2769 ( .A(b[11]), .B(n2358), .ZN(n1744) );
  XNOR2_X1 U2770 ( .A(b[17]), .B(n2358), .ZN(n1738) );
  XNOR2_X1 U2771 ( .A(b[13]), .B(n2357), .ZN(n1742) );
  INV_X1 U2772 ( .A(n325), .ZN(product[47]) );
  AOI21_X1 U2773 ( .B1(n423), .B2(n356), .A(n359), .ZN(n355) );
  NAND2_X1 U2774 ( .A1(n422), .A2(n356), .ZN(n354) );
  OAI22_X1 U2775 ( .A1(n2038), .A2(n1563), .B1(n2289), .B2(n1562), .ZN(n1271)
         );
  OAI22_X1 U2776 ( .A1(n2038), .A2(n1567), .B1(n2289), .B2(n1566), .ZN(n1275)
         );
  OAI22_X1 U2777 ( .A1(n2275), .A2(n1566), .B1(n1565), .B2(n2057), .ZN(n1274)
         );
  OAI22_X1 U2778 ( .A1(n2038), .A2(n1561), .B1(n2057), .B2(n1560), .ZN(n1269)
         );
  OAI22_X1 U2779 ( .A1(n2038), .A2(n1564), .B1(n1563), .B2(n2289), .ZN(n1272)
         );
  OAI22_X1 U2780 ( .A1(n2038), .A2(n1560), .B1(n1559), .B2(n2057), .ZN(n1268)
         );
  OAI22_X1 U2781 ( .A1(n2275), .A2(n1565), .B1(n2057), .B2(n1564), .ZN(n1273)
         );
  OAI22_X1 U2782 ( .A1(n2275), .A2(n2319), .B1(n1581), .B2(n2289), .ZN(n1185)
         );
  OAI22_X1 U2783 ( .A1(n2038), .A2(n1559), .B1(n2057), .B2(n1558), .ZN(n1267)
         );
  OAI22_X1 U2784 ( .A1(n2275), .A2(n1562), .B1(n1561), .B2(n2057), .ZN(n1270)
         );
  OAI22_X1 U2785 ( .A1(n2275), .A2(n1568), .B1(n1567), .B2(n2057), .ZN(n1276)
         );
  XNOR2_X1 U2786 ( .A(b[17]), .B(n2321), .ZN(n1588) );
  XNOR2_X1 U2787 ( .A(b[15]), .B(n2321), .ZN(n1590) );
  XNOR2_X1 U2788 ( .A(b[13]), .B(n2321), .ZN(n1592) );
  OAI22_X1 U2789 ( .A1(n2038), .A2(n1558), .B1(n1557), .B2(n2289), .ZN(n706)
         );
  XNOR2_X1 U2790 ( .A(b[19]), .B(n2321), .ZN(n1586) );
  XNOR2_X1 U2791 ( .A(b[21]), .B(n2321), .ZN(n1584) );
  XNOR2_X1 U2792 ( .A(b[11]), .B(n2321), .ZN(n1594) );
  OAI21_X1 U2793 ( .B1(n2265), .B2(n326), .A(n327), .ZN(n325) );
  NAND2_X1 U2794 ( .A1(n2071), .A2(n474), .ZN(n314) );
  OAI21_X1 U2795 ( .B1(n1933), .B2(n431), .A(n432), .ZN(n430) );
  OAI21_X1 U2796 ( .B1(n2051), .B2(n420), .A(n421), .ZN(n419) );
  OAI21_X1 U2797 ( .B1(n301), .B2(n438), .A(n439), .ZN(n437) );
  OAI21_X1 U2798 ( .B1(n2051), .B2(n411), .A(n412), .ZN(n410) );
  OAI21_X1 U2799 ( .B1(n301), .B2(n354), .A(n355), .ZN(n353) );
  OAI21_X1 U2800 ( .B1(n301), .B2(n371), .A(n372), .ZN(n370) );
  OAI21_X1 U2801 ( .B1(n1933), .B2(n380), .A(n381), .ZN(n379) );
  OAI21_X1 U2802 ( .B1(n2051), .B2(n343), .A(n344), .ZN(n342) );
  OAI21_X1 U2803 ( .B1(n1933), .B2(n398), .A(n399), .ZN(n397) );
  OAI21_X1 U2804 ( .B1(n2265), .B2(n389), .A(n390), .ZN(n388) );
  AOI21_X1 U2805 ( .B1(n2071), .B2(n483), .A(n1938), .ZN(n468) );
  NAND2_X1 U2806 ( .A1(n2071), .A2(n666), .ZN(n467) );
  OAI22_X1 U2807 ( .A1(n1984), .A2(n1691), .B1(n1690), .B2(n2036), .ZN(n1394)
         );
  OAI22_X1 U2808 ( .A1(n1984), .A2(n1686), .B1(n2036), .B2(n1685), .ZN(n1389)
         );
  OAI22_X1 U2809 ( .A1(n2108), .A2(n1689), .B1(n1688), .B2(n2297), .ZN(n1392)
         );
  OAI22_X1 U2810 ( .A1(n1984), .A2(n1690), .B1(n2297), .B2(n1689), .ZN(n1393)
         );
  OAI22_X1 U2811 ( .A1(n1984), .A2(n1692), .B1(n2036), .B2(n1691), .ZN(n1395)
         );
  OAI22_X1 U2812 ( .A1(n1984), .A2(n1685), .B1(n1684), .B2(n2036), .ZN(n1388)
         );
  OAI22_X1 U2813 ( .A1(n2108), .A2(n1688), .B1(n2297), .B2(n1687), .ZN(n1391)
         );
  OAI22_X1 U2814 ( .A1(n2278), .A2(n1684), .B1(n2035), .B2(n1683), .ZN(n1387)
         );
  OAI22_X1 U2815 ( .A1(n1984), .A2(n2348), .B1(n1706), .B2(n2297), .ZN(n1190)
         );
  OAI22_X1 U2816 ( .A1(n2278), .A2(n1693), .B1(n1692), .B2(n2035), .ZN(n1396)
         );
  XNOR2_X1 U2817 ( .A(b[13]), .B(n2008), .ZN(n1717) );
  XNOR2_X1 U2818 ( .A(b[21]), .B(n2007), .ZN(n1709) );
  XNOR2_X1 U2819 ( .A(b[15]), .B(n2008), .ZN(n1715) );
  XNOR2_X1 U2820 ( .A(b[11]), .B(n2008), .ZN(n1719) );
  XNOR2_X1 U2821 ( .A(b[19]), .B(n2008), .ZN(n1711) );
  XNOR2_X1 U2822 ( .A(b[17]), .B(n2007), .ZN(n1713) );
  INV_X2 U2823 ( .A(n2061), .ZN(n2275) );
  INV_X1 U2824 ( .A(n2158), .ZN(n2295) );
  INV_X1 U2825 ( .A(n2157), .ZN(n2300) );
  INV_X1 U2826 ( .A(n2037), .ZN(n2311) );
  INV_X1 U2827 ( .A(a[21]), .ZN(n2312) );
  INV_X1 U2828 ( .A(a[21]), .ZN(n2313) );
  INV_X1 U2829 ( .A(n2316), .ZN(n2315) );
  INV_X1 U2830 ( .A(a[19]), .ZN(n2316) );
  INV_X1 U2831 ( .A(n2320), .ZN(n2318) );
  INV_X1 U2832 ( .A(a[17]), .ZN(n2319) );
  INV_X1 U2833 ( .A(a[17]), .ZN(n2320) );
  INV_X1 U2834 ( .A(n2326), .ZN(n2324) );
  INV_X1 U2835 ( .A(a[15]), .ZN(n2325) );
  INV_X1 U2836 ( .A(a[15]), .ZN(n2326) );
  INV_X1 U2837 ( .A(n2331), .ZN(n2330) );
  INV_X1 U2838 ( .A(a[13]), .ZN(n2331) );
  INV_X1 U2839 ( .A(a[13]), .ZN(n2332) );
  INV_X1 U2840 ( .A(n2338), .ZN(n2336) );
  INV_X1 U2841 ( .A(a[11]), .ZN(n2338) );
  INV_X1 U2842 ( .A(n2343), .ZN(n2341) );
  INV_X1 U2843 ( .A(a[9]), .ZN(n2342) );
  INV_X1 U2844 ( .A(a[9]), .ZN(n2343) );
  INV_X1 U2845 ( .A(n2349), .ZN(n2347) );
  INV_X1 U2846 ( .A(a[7]), .ZN(n2348) );
  INV_X1 U2847 ( .A(a[7]), .ZN(n2349) );
  INV_X1 U2848 ( .A(n2355), .ZN(n2353) );
  INV_X1 U2849 ( .A(a[5]), .ZN(n2355) );
  INV_X1 U2850 ( .A(n2359), .ZN(n2358) );
  INV_X1 U2851 ( .A(a[3]), .ZN(n2359) );
  INV_X1 U2852 ( .A(n2363), .ZN(n2361) );
  INV_X1 U2853 ( .A(a[1]), .ZN(n2362) );
  INV_X1 U2854 ( .A(a[1]), .ZN(n2363) );
  INV_X2 U2855 ( .A(b[0]), .ZN(n2364) );
endmodule


module iir_filter_DW_mult_tc_4 ( a, b, product );
  input [23:0] a;
  input [23:0] b;
  output [47:0] product;
  wire   n251, n277, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n325, n326, n327, n332, n333, n334, n335, n336, n337,
         n339, n341, n342, n343, n344, n345, n346, n347, n348, n350, n352,
         n353, n354, n355, n356, n359, n360, n361, n362, n363, n364, n365,
         n367, n369, n370, n371, n372, n376, n378, n379, n380, n381, n382,
         n383, n384, n387, n388, n389, n390, n394, n396, n397, n398, n399,
         n400, n401, n402, n405, n407, n409, n410, n411, n412, n416, n418,
         n419, n420, n421, n422, n423, n426, n427, n428, n429, n430, n431,
         n432, n434, n435, n436, n437, n438, n439, n445, n450, n451, n452,
         n453, n454, n455, n456, n457, n459, n461, n462, n463, n464, n465,
         n466, n467, n468, n472, n474, n475, n476, n477, n478, n479, n480,
         n481, n483, n486, n487, n488, n489, n490, n491, n492, n495, n496,
         n497, n498, n499, n501, n502, n503, n504, n505, n506, n508, n511,
         n512, n513, n514, n515, n516, n517, n520, n521, n522, n524, n525,
         n526, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n543, n544, n545, n546, n547, n550, n551, n552, n553, n555,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n581, n582, n583, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n609, n610,
         n611, n620, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n643, n644, n645, n646, n657, n661,
         n662, n663, n666, n668, n672, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1809, n1812, n1814, n1817, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317;

  FA_X1 U546 ( .A(n1195), .B(n682), .CI(n1218), .CO(n678), .S(n679) );
  FA_X1 U547 ( .A(n683), .B(n1196), .CI(n686), .CO(n680), .S(n681) );
  FA_X1 U549 ( .A(n690), .B(n1242), .CI(n687), .CO(n684), .S(n685) );
  FA_X1 U550 ( .A(n1219), .B(n692), .CI(n1197), .CO(n686), .S(n687) );
  FA_X1 U551 ( .A(n691), .B(n698), .CI(n696), .CO(n688), .S(n689) );
  FA_X1 U552 ( .A(n1198), .B(n1220), .CI(n693), .CO(n690), .S(n691) );
  FA_X1 U554 ( .A(n702), .B(n699), .CI(n697), .CO(n694), .S(n695) );
  FA_X1 U555 ( .A(n1266), .B(n1243), .CI(n704), .CO(n696), .S(n697) );
  FA_X1 U556 ( .A(n1221), .B(n1199), .CI(n706), .CO(n698), .S(n699) );
  FA_X1 U557 ( .A(n710), .B(n712), .CI(n703), .CO(n700), .S(n701) );
  FA_X1 U558 ( .A(n714), .B(n1244), .CI(n705), .CO(n702), .S(n703) );
  FA_X1 U559 ( .A(n1222), .B(n1200), .CI(n707), .CO(n704), .S(n705) );
  FA_X1 U561 ( .A(n718), .B(n713), .CI(n711), .CO(n708), .S(n709) );
  FA_X1 U562 ( .A(n715), .B(n722), .CI(n720), .CO(n710), .S(n711) );
  FA_X1 U563 ( .A(n1245), .B(n1223), .CI(n1290), .CO(n712), .S(n713) );
  FA_X1 U564 ( .A(n1267), .B(n1201), .CI(n724), .CO(n714), .S(n715) );
  FA_X1 U565 ( .A(n728), .B(n721), .CI(n719), .CO(n716), .S(n717) );
  FA_X1 U566 ( .A(n723), .B(n732), .CI(n730), .CO(n718), .S(n719) );
  FA_X1 U567 ( .A(n1202), .B(n1246), .CI(n734), .CO(n720), .S(n721) );
  FA_X1 U568 ( .A(n1268), .B(n1224), .CI(n725), .CO(n722), .S(n723) );
  FA_X1 U570 ( .A(n738), .B(n731), .CI(n729), .CO(n726), .S(n727) );
  FA_X1 U571 ( .A(n735), .B(n733), .CI(n740), .CO(n728), .S(n729) );
  FA_X1 U572 ( .A(n744), .B(n1314), .CI(n742), .CO(n730), .S(n731) );
  FA_X1 U573 ( .A(n1225), .B(n1291), .CI(n1269), .CO(n732), .S(n733) );
  FA_X1 U574 ( .A(n746), .B(n1203), .CI(n1247), .CO(n734), .S(n735) );
  FA_X1 U575 ( .A(n750), .B(n741), .CI(n739), .CO(n736), .S(n737) );
  FA_X1 U576 ( .A(n754), .B(n745), .CI(n752), .CO(n738), .S(n739) );
  FA_X1 U577 ( .A(n756), .B(n758), .CI(n743), .CO(n740), .S(n741) );
  FA_X1 U578 ( .A(n1226), .B(n1204), .CI(n1270), .CO(n742), .S(n743) );
  FA_X1 U579 ( .A(n1292), .B(n1248), .CI(n747), .CO(n744), .S(n745) );
  FA_X1 U581 ( .A(n762), .B(n753), .CI(n751), .CO(n748), .S(n749) );
  FA_X1 U582 ( .A(n755), .B(n766), .CI(n764), .CO(n750), .S(n751) );
  FA_X1 U583 ( .A(n757), .B(n768), .CI(n759), .CO(n752), .S(n753) );
  FA_X1 U584 ( .A(n1338), .B(n1271), .CI(n770), .CO(n754), .S(n755) );
  FA_X1 U585 ( .A(n1249), .B(n1293), .CI(n1315), .CO(n756), .S(n757) );
  FA_X1 U586 ( .A(n772), .B(n1205), .CI(n1227), .CO(n758), .S(n759) );
  FA_X1 U587 ( .A(n776), .B(n765), .CI(n763), .CO(n760), .S(n761) );
  FA_X1 U589 ( .A(n771), .B(n769), .CI(n782), .CO(n764), .S(n765) );
  FA_X1 U590 ( .A(n786), .B(n1228), .CI(n784), .CO(n766), .S(n767) );
  FA_X1 U591 ( .A(n1294), .B(n1206), .CI(n1272), .CO(n768), .S(n769) );
  FA_X1 U592 ( .A(n1316), .B(n1250), .CI(n773), .CO(n770), .S(n771) );
  FA_X1 U594 ( .A(n790), .B(n779), .CI(n777), .CO(n774), .S(n775) );
  FA_X1 U596 ( .A(n796), .B(n787), .CI(n783), .CO(n778), .S(n779) );
  FA_X1 U597 ( .A(n798), .B(n800), .CI(n785), .CO(n780), .S(n781) );
  FA_X1 U598 ( .A(n1339), .B(n1229), .CI(n1362), .CO(n782), .S(n783) );
  FA_X1 U599 ( .A(n1273), .B(n1317), .CI(n1295), .CO(n784), .S(n785) );
  FA_X1 U600 ( .A(n1996), .B(n1207), .CI(n1251), .CO(n786), .S(n787) );
  FA_X1 U601 ( .A(n806), .B(n793), .CI(n791), .CO(n788), .S(n789) );
  FA_X1 U603 ( .A(n797), .B(n801), .CI(n812), .CO(n792), .S(n793) );
  FA_X1 U604 ( .A(n814), .B(n816), .CI(n799), .CO(n794), .S(n795) );
  FA_X1 U606 ( .A(n1208), .B(n1318), .CI(n1230), .CO(n798), .S(n799) );
  FA_X1 U607 ( .A(n1340), .B(n1252), .CI(n803), .CO(n800), .S(n801) );
  FA_X1 U609 ( .A(n822), .B(n809), .CI(n807), .CO(n804), .S(n805) );
  FA_X1 U610 ( .A(n811), .B(n826), .CI(n824), .CO(n806), .S(n807) );
  FA_X1 U612 ( .A(n815), .B(n832), .CI(n817), .CO(n810), .S(n811) );
  FA_X1 U613 ( .A(n830), .B(n1386), .CI(n834), .CO(n812), .S(n813) );
  FA_X1 U614 ( .A(n1319), .B(n1253), .CI(n1341), .CO(n814), .S(n815) );
  FA_X1 U615 ( .A(n1231), .B(n1297), .CI(n1275), .CO(n816), .S(n817) );
  FA_X1 U616 ( .A(n1363), .B(n1209), .CI(n2032), .CO(n818), .S(n819) );
  FA_X1 U617 ( .A(n840), .B(n825), .CI(n823), .CO(n820), .S(n821) );
  FA_X1 U619 ( .A(n846), .B(n848), .CI(n829), .CO(n824), .S(n825) );
  FA_X1 U620 ( .A(n835), .B(n831), .CI(n833), .CO(n826), .S(n827) );
  FA_X1 U621 ( .A(n850), .B(n854), .CI(n852), .CO(n828), .S(n829) );
  FA_X1 U622 ( .A(n1254), .B(n1320), .CI(n1298), .CO(n830), .S(n831) );
  FA_X1 U623 ( .A(n1232), .B(n1364), .CI(n1342), .CO(n832), .S(n833) );
  FA_X1 U624 ( .A(n1210), .B(n1276), .CI(n837), .CO(n834), .S(n835) );
  FA_X1 U626 ( .A(n858), .B(n843), .CI(n841), .CO(n838), .S(n839) );
  FA_X1 U627 ( .A(n845), .B(n847), .CI(n860), .CO(n840), .S(n841) );
  FA_X1 U629 ( .A(n855), .B(n853), .CI(n866), .CO(n844), .S(n845) );
  FA_X1 U630 ( .A(n868), .B(n870), .CI(n851), .CO(n846), .S(n847) );
  FA_X1 U631 ( .A(n1410), .B(n1365), .CI(n872), .CO(n848), .S(n849) );
  FA_X1 U632 ( .A(n1299), .B(n1277), .CI(n1343), .CO(n850), .S(n851) );
  FA_X1 U633 ( .A(n1255), .B(n1321), .CI(n1962), .CO(n852), .S(n853) );
  FA_X1 U634 ( .A(n1233), .B(n1211), .CI(n1387), .CO(n854), .S(n855) );
  FA_X1 U637 ( .A(n884), .B(n867), .CI(n865), .CO(n860), .S(n861) );
  FA_X1 U638 ( .A(n888), .B(n873), .CI(n886), .CO(n862), .S(n863) );
  FA_X1 U639 ( .A(n869), .B(n890), .CI(n871), .CO(n864), .S(n865) );
  FA_X1 U640 ( .A(n894), .B(n1300), .CI(n892), .CO(n866), .S(n867) );
  FA_X1 U641 ( .A(n1234), .B(n1322), .CI(n1256), .CO(n868), .S(n869) );
  FA_X1 U642 ( .A(n1366), .B(n1212), .CI(n1344), .CO(n870), .S(n871) );
  FA_X1 U643 ( .A(n1388), .B(n1278), .CI(n875), .CO(n872), .S(n873) );
  FA_X1 U645 ( .A(n898), .B(n881), .CI(n879), .CO(n876), .S(n877) );
  FA_X1 U646 ( .A(n883), .B(n885), .CI(n900), .CO(n878), .S(n879) );
  FA_X1 U647 ( .A(n887), .B(n904), .CI(n902), .CO(n880), .S(n881) );
  FA_X1 U648 ( .A(n889), .B(n893), .CI(n906), .CO(n882), .S(n883) );
  FA_X1 U649 ( .A(n891), .B(n908), .CI(n895), .CO(n884), .S(n885) );
  FA_X1 U650 ( .A(n912), .B(n910), .CI(n914), .CO(n886), .S(n887) );
  FA_X1 U651 ( .A(n1367), .B(n1389), .CI(n1434), .CO(n888), .S(n889) );
  FA_X1 U652 ( .A(n1257), .B(n1301), .CI(n1345), .CO(n890), .S(n891) );
  FA_X1 U653 ( .A(n2204), .B(n1323), .CI(n1279), .CO(n892), .S(n893) );
  FA_X1 U654 ( .A(n1235), .B(n1213), .CI(n1411), .CO(n894), .S(n895) );
  FA_X1 U656 ( .A(n903), .B(n924), .CI(n922), .CO(n898), .S(n899) );
  FA_X1 U657 ( .A(n907), .B(n926), .CI(n905), .CO(n900), .S(n901) );
  FA_X1 U658 ( .A(n909), .B(n930), .CI(n928), .CO(n902), .S(n903) );
  FA_X1 U659 ( .A(n911), .B(n913), .CI(n915), .CO(n904), .S(n905) );
  FA_X1 U660 ( .A(n934), .B(n936), .CI(n932), .CO(n906), .S(n907) );
  FA_X1 U661 ( .A(n1368), .B(n1390), .CI(n938), .CO(n908), .S(n909) );
  FA_X1 U662 ( .A(n1280), .B(n1346), .CI(n1324), .CO(n910), .S(n911) );
  FA_X1 U663 ( .A(n1258), .B(n1236), .CI(n1412), .CO(n912), .S(n913) );
  FA_X1 U664 ( .A(n1214), .B(n1302), .CI(n917), .CO(n914), .S(n915) );
  FA_X1 U667 ( .A(n925), .B(n927), .CI(n944), .CO(n920), .S(n921) );
  FA_X1 U668 ( .A(n929), .B(n948), .CI(n946), .CO(n922), .S(n923) );
  FA_X1 U669 ( .A(n950), .B(n935), .CI(n931), .CO(n924), .S(n925) );
  FA_X1 U670 ( .A(n937), .B(n933), .CI(n952), .CO(n926), .S(n927) );
  FA_X1 U671 ( .A(n956), .B(n958), .CI(n954), .CO(n928), .S(n929) );
  FA_X1 U672 ( .A(n939), .B(n1939), .CI(n1458), .CO(n930), .S(n931) );
  FA_X1 U673 ( .A(n1325), .B(n1435), .CI(n1413), .CO(n932), .S(n933) );
  FA_X1 U674 ( .A(n1281), .B(n1369), .CI(n1391), .CO(n934), .S(n935) );
  FA_X1 U675 ( .A(n1259), .B(n1303), .CI(n1347), .CO(n936), .S(n937) );
  FA_X1 U678 ( .A(n964), .B(n945), .CI(n943), .CO(n940), .S(n941) );
  FA_X1 U680 ( .A(n951), .B(n970), .CI(n968), .CO(n944), .S(n945) );
  FA_X1 U681 ( .A(n972), .B(n959), .CI(n953), .CO(n946), .S(n947) );
  FA_X1 U682 ( .A(n955), .B(n974), .CI(n957), .CO(n948), .S(n949) );
  FA_X1 U683 ( .A(n976), .B(n980), .CI(n978), .CO(n950), .S(n951) );
  FA_X1 U684 ( .A(n1326), .B(n1392), .CI(n961), .CO(n952), .S(n953) );
  FA_X1 U685 ( .A(n1282), .B(n1304), .CI(n1414), .CO(n954), .S(n955) );
  FA_X1 U689 ( .A(n984), .B(n967), .CI(n965), .CO(n962), .S(n963) );
  FA_X1 U690 ( .A(n969), .B(n971), .CI(n986), .CO(n964), .S(n965) );
  FA_X1 U691 ( .A(n973), .B(n990), .CI(n988), .CO(n966), .S(n967) );
  FA_X1 U692 ( .A(n975), .B(n981), .CI(n992), .CO(n968), .S(n969) );
  FA_X1 U693 ( .A(n977), .B(n998), .CI(n979), .CO(n970), .S(n971) );
  FA_X1 U696 ( .A(n1305), .B(n1437), .CI(n1327), .CO(n976), .S(n977) );
  FA_X1 U697 ( .A(n1460), .B(n1371), .CI(n1283), .CO(n978), .S(n979) );
  FA_X1 U698 ( .A(n1239), .B(n1349), .CI(n1261), .CO(n980), .S(n981) );
  FA_X1 U699 ( .A(n1004), .B(n987), .CI(n985), .CO(n982), .S(n983) );
  FA_X1 U700 ( .A(n989), .B(n991), .CI(n1006), .CO(n984), .S(n985) );
  FA_X1 U701 ( .A(n993), .B(n1010), .CI(n1008), .CO(n986), .S(n987) );
  FA_X1 U702 ( .A(n999), .B(n997), .CI(n1012), .CO(n988), .S(n989) );
  FA_X1 U703 ( .A(n1014), .B(n1016), .CI(n995), .CO(n990), .S(n991) );
  FA_X1 U704 ( .A(n1018), .B(n1394), .CI(n1001), .CO(n992), .S(n993) );
  FA_X1 U705 ( .A(n1306), .B(n1328), .CI(n1416), .CO(n994), .S(n995) );
  FA_X1 U707 ( .A(n1461), .B(n1350), .CI(n1183), .CO(n998), .S(n999) );
  HA_X1 U708 ( .A(n1240), .B(n1262), .CO(n1000), .S(n1001) );
  FA_X1 U709 ( .A(n1022), .B(n1007), .CI(n1005), .CO(n1002), .S(n1003) );
  FA_X1 U710 ( .A(n1009), .B(n1011), .CI(n1024), .CO(n1004), .S(n1005) );
  FA_X1 U711 ( .A(n1013), .B(n1028), .CI(n1026), .CO(n1006), .S(n1007) );
  FA_X1 U712 ( .A(n1015), .B(n1019), .CI(n1017), .CO(n1008), .S(n1009) );
  FA_X1 U713 ( .A(n1030), .B(n1034), .CI(n1241), .CO(n1010), .S(n1011) );
  FA_X1 U714 ( .A(n1036), .B(n1439), .CI(n1032), .CO(n1012), .S(n1013) );
  FA_X1 U715 ( .A(n1395), .B(n1462), .CI(n1417), .CO(n1014), .S(n1015) );
  FA_X1 U716 ( .A(n1307), .B(n1373), .CI(n1329), .CO(n1016), .S(n1017) );
  FA_X1 U717 ( .A(n1351), .B(n1285), .CI(n1263), .CO(n1018), .S(n1019) );
  FA_X1 U718 ( .A(n1040), .B(n1025), .CI(n1023), .CO(n1020), .S(n1021) );
  FA_X1 U719 ( .A(n1027), .B(n1044), .CI(n1042), .CO(n1022), .S(n1023) );
  FA_X1 U720 ( .A(n1046), .B(n1035), .CI(n1029), .CO(n1024), .S(n1025) );
  FA_X1 U721 ( .A(n1031), .B(n1048), .CI(n1033), .CO(n1026), .S(n1027) );
  FA_X1 U722 ( .A(n1052), .B(n1037), .CI(n1050), .CO(n1028), .S(n1029) );
  FA_X1 U723 ( .A(n1352), .B(n1440), .CI(n1418), .CO(n1030), .S(n1031) );
  FA_X1 U724 ( .A(n1396), .B(n1330), .CI(n1463), .CO(n1032), .S(n1033) );
  FA_X1 U725 ( .A(n1308), .B(n1374), .CI(n1184), .CO(n1034), .S(n1035) );
  HA_X1 U726 ( .A(n1264), .B(n1286), .CO(n1036), .S(n1037) );
  FA_X1 U727 ( .A(n1056), .B(n1043), .CI(n1041), .CO(n1038), .S(n1039) );
  FA_X1 U729 ( .A(n1062), .B(n1053), .CI(n1060), .CO(n1042), .S(n1043) );
  FA_X1 U730 ( .A(n1049), .B(n1265), .CI(n1051), .CO(n1044), .S(n1045) );
  FA_X1 U731 ( .A(n1064), .B(n1068), .CI(n1066), .CO(n1046), .S(n1047) );
  FA_X1 U732 ( .A(n1397), .B(n1441), .CI(n1419), .CO(n1048), .S(n1049) );
  FA_X1 U733 ( .A(n1331), .B(n1353), .CI(n1375), .CO(n1050), .S(n1051) );
  FA_X1 U734 ( .A(n1309), .B(n1287), .CI(n1464), .CO(n1052), .S(n1053) );
  FA_X1 U735 ( .A(n1072), .B(n1059), .CI(n1057), .CO(n1054), .S(n1055) );
  FA_X1 U736 ( .A(n1074), .B(n1063), .CI(n1061), .CO(n1056), .S(n1057) );
  FA_X1 U738 ( .A(n1080), .B(n1082), .CI(n1078), .CO(n1060), .S(n1061) );
  FA_X1 U739 ( .A(n1398), .B(n1420), .CI(n1069), .CO(n1062), .S(n1063) );
  FA_X1 U740 ( .A(n1442), .B(n1354), .CI(n1332), .CO(n1064), .S(n1065) );
  FA_X1 U741 ( .A(n1465), .B(n1376), .CI(n1185), .CO(n1066), .S(n1067) );
  HA_X1 U742 ( .A(n1288), .B(n1310), .CO(n1068), .S(n1069) );
  FA_X1 U743 ( .A(n1086), .B(n1075), .CI(n1073), .CO(n1070), .S(n1071) );
  FA_X1 U744 ( .A(n1088), .B(n1090), .CI(n1077), .CO(n1072), .S(n1073) );
  FA_X1 U745 ( .A(n1083), .B(n1081), .CI(n1079), .CO(n1074), .S(n1075) );
  FA_X1 U746 ( .A(n1092), .B(n1094), .CI(n1289), .CO(n1076), .S(n1077) );
  FA_X1 U747 ( .A(n1399), .B(n1421), .CI(n1096), .CO(n1078), .S(n1079) );
  FA_X1 U748 ( .A(n1377), .B(n1443), .CI(n1355), .CO(n1080), .S(n1081) );
  FA_X1 U749 ( .A(n1311), .B(n1333), .CI(n1466), .CO(n1082), .S(n1083) );
  FA_X1 U750 ( .A(n1100), .B(n1089), .CI(n1087), .CO(n1084), .S(n1085) );
  FA_X1 U751 ( .A(n1102), .B(n1104), .CI(n1091), .CO(n1086), .S(n1087) );
  FA_X1 U752 ( .A(n1093), .B(n1106), .CI(n1095), .CO(n1088), .S(n1089) );
  FA_X1 U753 ( .A(n1097), .B(n1422), .CI(n1108), .CO(n1090), .S(n1091) );
  FA_X1 U754 ( .A(n1356), .B(n1444), .CI(n1378), .CO(n1092), .S(n1093) );
  FA_X1 U755 ( .A(n1467), .B(n1186), .CI(n1400), .CO(n1094), .S(n1095) );
  HA_X1 U756 ( .A(n1312), .B(n1334), .CO(n1096), .S(n1097) );
  FA_X1 U757 ( .A(n1103), .B(n1112), .CI(n1101), .CO(n1098), .S(n1099) );
  FA_X1 U758 ( .A(n1114), .B(n1109), .CI(n1105), .CO(n1100), .S(n1101) );
  FA_X1 U759 ( .A(n1313), .B(n1116), .CI(n1107), .CO(n1102), .S(n1103) );
  FA_X1 U760 ( .A(n1120), .B(n1423), .CI(n1118), .CO(n1104), .S(n1105) );
  FA_X1 U761 ( .A(n1379), .B(n1445), .CI(n1401), .CO(n1106), .S(n1107) );
  FA_X1 U762 ( .A(n1335), .B(n1468), .CI(n1357), .CO(n1108), .S(n1109) );
  FA_X1 U763 ( .A(n1124), .B(n1115), .CI(n1113), .CO(n1110), .S(n1111) );
  FA_X1 U764 ( .A(n1119), .B(n1117), .CI(n1126), .CO(n1112), .S(n1113) );
  FA_X1 U765 ( .A(n1130), .B(n1121), .CI(n1128), .CO(n1114), .S(n1115) );
  FA_X1 U766 ( .A(n1380), .B(n1446), .CI(n1424), .CO(n1116), .S(n1117) );
  FA_X1 U767 ( .A(n1469), .B(n1402), .CI(n1187), .CO(n1118), .S(n1119) );
  HA_X1 U768 ( .A(n1336), .B(n1358), .CO(n1120), .S(n1121) );
  FA_X1 U769 ( .A(n1127), .B(n1134), .CI(n1125), .CO(n1122), .S(n1123) );
  FA_X1 U770 ( .A(n1131), .B(n1129), .CI(n1136), .CO(n1124), .S(n1125) );
  FA_X1 U771 ( .A(n1138), .B(n1140), .CI(n1337), .CO(n1126), .S(n1127) );
  FA_X1 U772 ( .A(n1403), .B(n1447), .CI(n1425), .CO(n1128), .S(n1129) );
  FA_X1 U773 ( .A(n1359), .B(n1470), .CI(n1381), .CO(n1130), .S(n1131) );
  FA_X1 U774 ( .A(n1144), .B(n1137), .CI(n1135), .CO(n1132), .S(n1133) );
  FA_X1 U775 ( .A(n1146), .B(n1148), .CI(n1139), .CO(n1134), .S(n1135) );
  FA_X1 U776 ( .A(n1404), .B(n1448), .CI(n1141), .CO(n1136), .S(n1137) );
  FA_X1 U777 ( .A(n1188), .B(n1426), .CI(n1471), .CO(n1138), .S(n1139) );
  HA_X1 U778 ( .A(n1360), .B(n1382), .CO(n1140), .S(n1141) );
  FA_X1 U779 ( .A(n1152), .B(n1147), .CI(n1145), .CO(n1142), .S(n1143) );
  FA_X1 U780 ( .A(n1361), .B(n1154), .CI(n1149), .CO(n1144), .S(n1145) );
  FA_X1 U781 ( .A(n1427), .B(n1449), .CI(n1156), .CO(n1146), .S(n1147) );
  FA_X1 U782 ( .A(n1383), .B(n1472), .CI(n1405), .CO(n1148), .S(n1149) );
  FA_X1 U783 ( .A(n1160), .B(n1155), .CI(n1153), .CO(n1150), .S(n1151) );
  FA_X1 U784 ( .A(n1157), .B(n1473), .CI(n1162), .CO(n1152), .S(n1153) );
  FA_X1 U785 ( .A(n1450), .B(n1428), .CI(n1189), .CO(n1154), .S(n1155) );
  HA_X1 U786 ( .A(n1384), .B(n1406), .CO(n1156), .S(n1157) );
  FA_X1 U787 ( .A(n1163), .B(n1385), .CI(n1164), .CO(n1158), .S(n1159) );
  FA_X1 U788 ( .A(n1168), .B(n1429), .CI(n1166), .CO(n1160), .S(n1161) );
  FA_X1 U789 ( .A(n1451), .B(n1474), .CI(n1407), .CO(n1162), .S(n1163) );
  FA_X1 U790 ( .A(n1172), .B(n1169), .CI(n1167), .CO(n1164), .S(n1165) );
  FA_X1 U791 ( .A(n1452), .B(n1475), .CI(n1190), .CO(n1166), .S(n1167) );
  HA_X1 U792 ( .A(n1408), .B(n1430), .CO(n1168), .S(n1169) );
  FA_X1 U793 ( .A(n1409), .B(n1176), .CI(n1173), .CO(n1170), .S(n1171) );
  FA_X1 U794 ( .A(n1476), .B(n1453), .CI(n1431), .CO(n1172), .S(n1173) );
  FA_X1 U795 ( .A(n1191), .B(n1454), .CI(n1177), .CO(n1174), .S(n1175) );
  HA_X1 U796 ( .A(n1432), .B(n1477), .CO(n1176), .S(n1177) );
  FA_X1 U797 ( .A(n1455), .B(n1478), .CI(n1180), .CO(n1178), .S(n1179) );
  HA_X1 U798 ( .A(n1456), .B(n1479), .CO(n1180), .S(n1181) );
  OR2_X1 U1448 ( .A1(n1021), .A2(n1038), .ZN(n1929) );
  INV_X2 U1449 ( .A(n2294), .ZN(n2291) );
  INV_X1 U1450 ( .A(n2059), .ZN(n2061) );
  XOR2_X1 U1451 ( .A(b[3]), .B(n2270), .Z(n1627) );
  INV_X1 U1452 ( .A(n2270), .ZN(n2267) );
  INV_X1 U1453 ( .A(n2139), .ZN(n1931) );
  INV_X1 U1454 ( .A(n2139), .ZN(n1930) );
  INV_X1 U1455 ( .A(n2139), .ZN(n2072) );
  NOR2_X1 U1456 ( .A1(n531), .A2(n534), .ZN(n1932) );
  NOR2_X1 U1457 ( .A1(n919), .A2(n940), .ZN(n1933) );
  CLKBUF_X3 U1458 ( .A(n1957), .Z(n2149) );
  INV_X1 U1459 ( .A(n2170), .ZN(n1934) );
  INV_X2 U1460 ( .A(n1985), .ZN(n2230) );
  OR2_X1 U1461 ( .A1(n558), .A2(n563), .ZN(n1935) );
  CLKBUF_X1 U1462 ( .A(n511), .Z(n1936) );
  INV_X2 U1463 ( .A(n2261), .ZN(n2258) );
  INV_X1 U1464 ( .A(n1966), .ZN(n2238) );
  INV_X2 U1465 ( .A(n1966), .ZN(n2239) );
  NAND3_X1 U1466 ( .A1(n2018), .A2(n2019), .A3(n2020), .ZN(n1938) );
  NAND3_X1 U1467 ( .A1(n2018), .A2(n2019), .A3(n2020), .ZN(n1937) );
  INV_X1 U1468 ( .A(n2014), .ZN(n2175) );
  INV_X1 U1469 ( .A(n2149), .ZN(n2142) );
  INV_X1 U1470 ( .A(n2169), .ZN(n2237) );
  INV_X1 U1471 ( .A(n2141), .ZN(n2095) );
  AND2_X1 U1472 ( .A1(n1967), .A2(n1216), .ZN(n1939) );
  AND2_X1 U1473 ( .A1(n1111), .A2(n1122), .ZN(n1940) );
  AND2_X1 U1474 ( .A1(n1021), .A2(n1038), .ZN(n1941) );
  OR2_X1 U1475 ( .A1(n1945), .A2(n982), .ZN(n1942) );
  XNOR2_X1 U1476 ( .A(n560), .B(n1943), .ZN(product[22]) );
  AND2_X1 U1477 ( .A1(n1942), .A2(n559), .ZN(n1943) );
  XNOR2_X1 U1478 ( .A(n301), .B(n1944), .ZN(product[34]) );
  AND2_X1 U1479 ( .A1(n663), .A2(n439), .ZN(n1944) );
  INV_X2 U1480 ( .A(n2139), .ZN(n2215) );
  CLKBUF_X1 U1481 ( .A(n963), .Z(n1945) );
  INV_X2 U1482 ( .A(n2135), .ZN(n2213) );
  INV_X1 U1483 ( .A(n2270), .ZN(n1988) );
  INV_X1 U1484 ( .A(n2270), .ZN(n1989) );
  BUF_X1 U1485 ( .A(n536), .Z(n1946) );
  BUF_X1 U1486 ( .A(n536), .Z(n1948) );
  BUF_X1 U1487 ( .A(n536), .Z(n1947) );
  INV_X1 U1488 ( .A(a[23]), .ZN(n1949) );
  BUF_X2 U1489 ( .A(n2070), .Z(n2146) );
  INV_X1 U1490 ( .A(n2070), .ZN(n2170) );
  INV_X1 U1491 ( .A(n2062), .ZN(n2167) );
  BUF_X2 U1492 ( .A(a[5]), .Z(n1978) );
  XOR2_X1 U1493 ( .A(a[20]), .B(a[19]), .Z(n1950) );
  NOR2_X1 U1494 ( .A1(n1003), .A2(n1020), .ZN(n1951) );
  CLKBUF_X1 U1495 ( .A(n581), .Z(n1952) );
  XNOR2_X1 U1496 ( .A(n966), .B(n1953), .ZN(n943) );
  XNOR2_X1 U1497 ( .A(n947), .B(n949), .ZN(n1953) );
  OR2_X1 U1498 ( .A1(n941), .A2(n962), .ZN(n1954) );
  XNOR2_X1 U1499 ( .A(a[18]), .B(n2254), .ZN(n2098) );
  CLKBUF_X1 U1500 ( .A(n781), .Z(n1955) );
  XNOR2_X1 U1501 ( .A(b[3]), .B(n2246), .ZN(n1956) );
  XNOR2_X1 U1502 ( .A(a[10]), .B(n2275), .ZN(n1812) );
  OR2_X2 U1503 ( .A1(n1958), .A2(n2059), .ZN(n1957) );
  XNOR2_X1 U1504 ( .A(a[4]), .B(n2290), .ZN(n1958) );
  CLKBUF_X1 U1505 ( .A(n1957), .Z(n1959) );
  INV_X1 U1506 ( .A(n2265), .ZN(n1961) );
  INV_X1 U1507 ( .A(n2265), .ZN(n1960) );
  OAI22_X1 U1508 ( .A1(n1959), .A2(n1708), .B1(n1707), .B2(n2237), .ZN(n1962)
         );
  CLKBUF_X1 U1509 ( .A(n839), .Z(n1963) );
  INV_X1 U1510 ( .A(n2040), .ZN(n1964) );
  NOR2_X1 U1511 ( .A1(n963), .A2(n982), .ZN(n1965) );
  NOR2_X1 U1512 ( .A1(n963), .A2(n982), .ZN(n558) );
  BUF_X1 U1513 ( .A(n2165), .Z(n1966) );
  OAI22_X1 U1514 ( .A1(n2077), .A2(n1528), .B1(n1956), .B2(n2225), .ZN(n1967)
         );
  INV_X2 U1515 ( .A(n2298), .ZN(n1968) );
  INV_X2 U1516 ( .A(n2169), .ZN(n1969) );
  INV_X1 U1517 ( .A(n2136), .ZN(n1970) );
  OAI22_X1 U1518 ( .A1(n2205), .A2(n1505), .B1(n1504), .B2(n2147), .ZN(n1971)
         );
  INV_X1 U1519 ( .A(n2250), .ZN(n1973) );
  INV_X1 U1520 ( .A(n2250), .ZN(n1972) );
  AND2_X1 U1521 ( .A1(n1817), .A2(n2240), .ZN(n1974) );
  INV_X1 U1522 ( .A(n672), .ZN(n1975) );
  XNOR2_X1 U1523 ( .A(a[2]), .B(a[3]), .ZN(n2140) );
  INV_X2 U1524 ( .A(n2134), .ZN(n1977) );
  INV_X1 U1525 ( .A(n2134), .ZN(n1976) );
  INV_X1 U1526 ( .A(n2134), .ZN(n2210) );
  INV_X1 U1527 ( .A(n2139), .ZN(n2073) );
  INV_X1 U1528 ( .A(n492), .ZN(n1979) );
  XOR2_X1 U1529 ( .A(a[22]), .B(a[21]), .Z(n1980) );
  XOR2_X1 U1530 ( .A(a[10]), .B(n2282), .Z(n1981) );
  CLKBUF_X1 U1531 ( .A(n489), .Z(n1982) );
  CLKBUF_X1 U1532 ( .A(a[3]), .Z(n1983) );
  BUF_X1 U1533 ( .A(n2056), .Z(n1984) );
  XOR2_X1 U1534 ( .A(a[14]), .B(a[13]), .Z(n1985) );
  XOR2_X1 U1535 ( .A(a[14]), .B(a[13]), .Z(n2133) );
  XNOR2_X1 U1536 ( .A(a[6]), .B(n1978), .ZN(n1986) );
  INV_X1 U1537 ( .A(n2279), .ZN(n1987) );
  INV_X2 U1538 ( .A(n2281), .ZN(n2279) );
  XNOR2_X1 U1539 ( .A(a[18]), .B(a[17]), .ZN(n2079) );
  INV_X1 U1540 ( .A(n2131), .ZN(n1990) );
  INV_X1 U1541 ( .A(n2271), .ZN(n1992) );
  INV_X1 U1542 ( .A(n2271), .ZN(n1991) );
  CLKBUF_X1 U1543 ( .A(n877), .Z(n1993) );
  INV_X1 U1544 ( .A(n2154), .ZN(n1994) );
  CLKBUF_X3 U1545 ( .A(n1981), .Z(n2154) );
  XNOR2_X1 U1546 ( .A(a[10]), .B(n2281), .ZN(n2194) );
  XNOR2_X1 U1547 ( .A(n2033), .B(n921), .ZN(n1995) );
  OAI22_X1 U1548 ( .A1(n2217), .A2(n1658), .B1(n1657), .B2(n2150), .ZN(n1996)
         );
  OAI21_X1 U1549 ( .B1(n535), .B2(n2042), .A(n532), .ZN(n1997) );
  XNOR2_X1 U1550 ( .A(a[6]), .B(n2288), .ZN(n1814) );
  XOR2_X1 U1551 ( .A(a[2]), .B(a[1]), .Z(n2165) );
  INV_X1 U1552 ( .A(n2132), .ZN(n1999) );
  INV_X1 U1553 ( .A(n1974), .ZN(n1998) );
  XOR2_X1 U1554 ( .A(n781), .B(n794), .Z(n2000) );
  XOR2_X1 U1555 ( .A(n792), .B(n2000), .Z(n777) );
  NAND2_X1 U1556 ( .A1(n792), .A2(n1955), .ZN(n2001) );
  NAND2_X1 U1557 ( .A1(n792), .A2(n794), .ZN(n2002) );
  NAND2_X1 U1558 ( .A1(n1955), .A2(n794), .ZN(n2003) );
  NAND3_X1 U1559 ( .A1(n2001), .A2(n2002), .A3(n2003), .ZN(n776) );
  INV_X1 U1560 ( .A(n2141), .ZN(n2004) );
  OR2_X2 U1561 ( .A1(n775), .A2(n788), .ZN(n2102) );
  INV_X1 U1562 ( .A(n2239), .ZN(n2005) );
  XOR2_X1 U1563 ( .A(a[20]), .B(a[19]), .Z(n2161) );
  INV_X1 U1564 ( .A(n2141), .ZN(n2218) );
  INV_X2 U1565 ( .A(n1949), .ZN(n2242) );
  XOR2_X1 U1566 ( .A(n813), .B(n819), .Z(n2006) );
  XOR2_X1 U1567 ( .A(n828), .B(n2006), .Z(n809) );
  NAND2_X1 U1568 ( .A1(n828), .A2(n813), .ZN(n2007) );
  NAND2_X1 U1569 ( .A1(n828), .A2(n819), .ZN(n2008) );
  NAND2_X1 U1570 ( .A1(n813), .A2(n819), .ZN(n2009) );
  NAND3_X1 U1571 ( .A1(n2007), .A2(n2008), .A3(n2009), .ZN(n808) );
  NOR2_X1 U1572 ( .A1(n456), .A2(n480), .ZN(n2010) );
  BUF_X2 U1573 ( .A(n277), .Z(n2012) );
  CLKBUF_X2 U1574 ( .A(n277), .Z(n2011) );
  CLKBUF_X1 U1575 ( .A(n277), .Z(n2155) );
  XNOR2_X1 U1576 ( .A(n2013), .B(n1058), .ZN(n1041) );
  XNOR2_X1 U1577 ( .A(n1047), .B(n1045), .ZN(n2013) );
  XNOR2_X1 U1578 ( .A(a[8]), .B(a[7]), .ZN(n2014) );
  INV_X2 U1579 ( .A(n2175), .ZN(n2234) );
  OR2_X2 U1580 ( .A1(n2133), .A2(n2138), .ZN(n2015) );
  CLKBUF_X1 U1581 ( .A(n805), .Z(n2016) );
  XOR2_X1 U1582 ( .A(n849), .B(n864), .Z(n2017) );
  XOR2_X1 U1583 ( .A(n862), .B(n2017), .Z(n843) );
  NAND2_X1 U1584 ( .A1(n862), .A2(n849), .ZN(n2018) );
  NAND2_X1 U1585 ( .A1(n862), .A2(n864), .ZN(n2019) );
  NAND2_X1 U1586 ( .A1(n849), .A2(n864), .ZN(n2020) );
  NAND3_X1 U1587 ( .A1(n2018), .A2(n2019), .A3(n2020), .ZN(n842) );
  AND2_X2 U1588 ( .A1(n2098), .A2(n2079), .ZN(n2131) );
  INV_X1 U1589 ( .A(n2131), .ZN(n2208) );
  NAND2_X1 U1590 ( .A1(n966), .A2(n947), .ZN(n2021) );
  NAND2_X1 U1591 ( .A1(n966), .A2(n949), .ZN(n2022) );
  NAND2_X1 U1592 ( .A1(n947), .A2(n949), .ZN(n2023) );
  NAND3_X1 U1593 ( .A1(n2021), .A2(n2022), .A3(n2023), .ZN(n942) );
  XNOR2_X1 U1594 ( .A(n2024), .B(n859), .ZN(n857) );
  XNOR2_X1 U1595 ( .A(n878), .B(n861), .ZN(n2024) );
  XNOR2_X1 U1596 ( .A(a[21]), .B(a[20]), .ZN(n2145) );
  XOR2_X1 U1597 ( .A(n1067), .B(n1065), .Z(n2025) );
  XOR2_X1 U1598 ( .A(n2025), .B(n1076), .Z(n1059) );
  NAND2_X1 U1599 ( .A1(n1067), .A2(n1065), .ZN(n2026) );
  NAND2_X1 U1600 ( .A1(n1067), .A2(n1076), .ZN(n2027) );
  NAND2_X1 U1601 ( .A1(n1065), .A2(n1076), .ZN(n2028) );
  NAND3_X1 U1602 ( .A1(n2026), .A2(n2027), .A3(n2028), .ZN(n1058) );
  NAND2_X1 U1603 ( .A1(n1047), .A2(n1045), .ZN(n2029) );
  NAND2_X1 U1604 ( .A1(n1047), .A2(n1058), .ZN(n2030) );
  NAND2_X1 U1605 ( .A1(n1045), .A2(n1058), .ZN(n2031) );
  NAND3_X1 U1606 ( .A1(n2029), .A2(n2030), .A3(n2031), .ZN(n1040) );
  INV_X2 U1607 ( .A(n2143), .ZN(n2216) );
  NOR2_X2 U1608 ( .A1(n789), .A2(n804), .ZN(n480) );
  OAI22_X1 U1609 ( .A1(n2095), .A2(n1683), .B1(n1682), .B2(n2236), .ZN(n2032)
         );
  XNOR2_X1 U1610 ( .A(n921), .B(n2033), .ZN(n919) );
  XNOR2_X1 U1611 ( .A(n942), .B(n923), .ZN(n2033) );
  BUF_X4 U1612 ( .A(n2243), .Z(n2152) );
  OAI22_X1 U1613 ( .A1(n2205), .A2(n1504), .B1(n2224), .B2(n1503), .ZN(n2034)
         );
  BUF_X1 U1614 ( .A(n553), .Z(n2041) );
  BUF_X4 U1615 ( .A(n251), .Z(n2240) );
  OR2_X1 U1616 ( .A1(n1964), .A2(n534), .ZN(n2035) );
  NAND2_X1 U1617 ( .A1(n921), .A2(n942), .ZN(n2036) );
  NAND2_X1 U1618 ( .A1(n921), .A2(n923), .ZN(n2037) );
  NAND2_X1 U1619 ( .A1(n942), .A2(n923), .ZN(n2038) );
  NAND3_X1 U1620 ( .A1(n2036), .A2(n2037), .A3(n2038), .ZN(n918) );
  BUF_X2 U1621 ( .A(n2079), .Z(n2151) );
  CLKBUF_X1 U1622 ( .A(a[8]), .Z(n2039) );
  OR2_X1 U1623 ( .A1(n896), .A2(n1993), .ZN(n2040) );
  XNOR2_X1 U1624 ( .A(a[4]), .B(a[3]), .ZN(n2078) );
  NOR2_X1 U1625 ( .A1(n877), .A2(n896), .ZN(n2042) );
  INV_X1 U1626 ( .A(n1935), .ZN(n2043) );
  XOR2_X1 U1627 ( .A(n863), .B(n882), .Z(n2044) );
  XOR2_X1 U1628 ( .A(n2044), .B(n880), .Z(n859) );
  NAND2_X1 U1629 ( .A1(n863), .A2(n882), .ZN(n2045) );
  NAND2_X1 U1630 ( .A1(n863), .A2(n880), .ZN(n2046) );
  NAND2_X1 U1631 ( .A1(n882), .A2(n880), .ZN(n2047) );
  NAND3_X1 U1632 ( .A1(n2045), .A2(n2046), .A3(n2047), .ZN(n858) );
  NAND2_X1 U1633 ( .A1(n878), .A2(n861), .ZN(n2048) );
  NAND2_X1 U1634 ( .A1(n878), .A2(n859), .ZN(n2049) );
  NAND2_X1 U1635 ( .A1(n861), .A2(n859), .ZN(n2050) );
  NAND3_X1 U1636 ( .A1(n2048), .A2(n2049), .A3(n2050), .ZN(n856) );
  INV_X1 U1637 ( .A(n1954), .ZN(n2051) );
  NOR2_X1 U1638 ( .A1(n941), .A2(n962), .ZN(n547) );
  XOR2_X1 U1639 ( .A(n1348), .B(n1182), .Z(n2052) );
  XOR2_X1 U1640 ( .A(n2052), .B(n1260), .Z(n959) );
  NAND2_X1 U1641 ( .A1(n1260), .A2(n1348), .ZN(n2053) );
  NAND2_X1 U1642 ( .A1(n1260), .A2(n1182), .ZN(n2054) );
  NAND2_X1 U1643 ( .A1(n1348), .A2(n1182), .ZN(n2055) );
  NAND3_X1 U1644 ( .A1(n2053), .A2(n2054), .A3(n2055), .ZN(n958) );
  INV_X2 U1645 ( .A(n2254), .ZN(n2251) );
  NOR2_X1 U1646 ( .A1(n839), .A2(n856), .ZN(n2056) );
  OAI22_X1 U1647 ( .A1(n2077), .A2(n1527), .B1(n2225), .B2(n1526), .ZN(n2057)
         );
  INV_X1 U1648 ( .A(n2226), .ZN(n2058) );
  NOR2_X1 U1649 ( .A1(n839), .A2(n856), .ZN(n513) );
  INV_X1 U1650 ( .A(n2078), .ZN(n2059) );
  INV_X1 U1651 ( .A(n2059), .ZN(n2060) );
  INV_X1 U1652 ( .A(n2139), .ZN(n2214) );
  XNOR2_X1 U1653 ( .A(a[16]), .B(a[15]), .ZN(n2062) );
  INV_X2 U1654 ( .A(n2167), .ZN(n2228) );
  BUF_X2 U1655 ( .A(n2062), .Z(n2153) );
  NOR2_X1 U1656 ( .A1(n919), .A2(n940), .ZN(n2063) );
  XNOR2_X1 U1657 ( .A(n1372), .B(n2064), .ZN(n997) );
  XNOR2_X1 U1658 ( .A(n1284), .B(n1438), .ZN(n2064) );
  XOR2_X1 U1659 ( .A(n1274), .B(n1296), .Z(n2065) );
  XOR2_X1 U1660 ( .A(n818), .B(n2065), .Z(n797) );
  NAND2_X1 U1661 ( .A1(n818), .A2(n1274), .ZN(n2066) );
  NAND2_X1 U1662 ( .A1(n818), .A2(n1296), .ZN(n2067) );
  NAND2_X1 U1663 ( .A1(n1274), .A2(n1296), .ZN(n2068) );
  NAND3_X1 U1664 ( .A1(n2066), .A2(n2067), .A3(n2068), .ZN(n796) );
  XNOR2_X1 U1665 ( .A(a[22]), .B(n2244), .ZN(n2101) );
  INV_X1 U1666 ( .A(n2079), .ZN(n2176) );
  CLKBUF_X1 U1667 ( .A(n568), .Z(n2069) );
  INV_X1 U1668 ( .A(n2060), .ZN(n2169) );
  INV_X2 U1669 ( .A(n2134), .ZN(n2209) );
  XNOR2_X1 U1670 ( .A(a[12]), .B(a[11]), .ZN(n2070) );
  INV_X2 U1671 ( .A(n2170), .ZN(n2231) );
  XNOR2_X1 U1672 ( .A(a[21]), .B(a[22]), .ZN(n2071) );
  BUF_X2 U1673 ( .A(n2071), .Z(n2147) );
  INV_X1 U1674 ( .A(n2293), .ZN(n2290) );
  INV_X2 U1675 ( .A(n2293), .ZN(n2289) );
  XNOR2_X1 U1676 ( .A(n2039), .B(n2282), .ZN(n2099) );
  XOR2_X1 U1677 ( .A(n1971), .B(n1238), .Z(n961) );
  INV_X1 U1678 ( .A(n2077), .ZN(n2144) );
  INV_X2 U1679 ( .A(n2275), .ZN(n2272) );
  XNOR2_X1 U1680 ( .A(a[16]), .B(n2261), .ZN(n1809) );
  NAND2_X1 U1681 ( .A1(n1372), .A2(n1284), .ZN(n2074) );
  NAND2_X1 U1682 ( .A1(n1372), .A2(n1438), .ZN(n2075) );
  NAND2_X1 U1683 ( .A1(n1284), .A2(n1438), .ZN(n2076) );
  NAND3_X1 U1684 ( .A1(n2074), .A2(n2075), .A3(n2076), .ZN(n996) );
  OR2_X4 U1685 ( .A1(n1950), .A2(n2145), .ZN(n2077) );
  INV_X1 U1686 ( .A(n2303), .ZN(n2300) );
  INV_X2 U1687 ( .A(n2303), .ZN(n2299) );
  AND2_X2 U1688 ( .A1(n1814), .A2(n1986), .ZN(n2141) );
  XOR2_X1 U1689 ( .A(a[14]), .B(n2266), .Z(n2138) );
  INV_X1 U1690 ( .A(n2265), .ZN(n2262) );
  INV_X2 U1691 ( .A(n2176), .ZN(n2227) );
  INV_X2 U1692 ( .A(n2281), .ZN(n2278) );
  INV_X2 U1693 ( .A(n2297), .ZN(n2295) );
  OR2_X1 U1694 ( .A1(n1995), .A2(n940), .ZN(n2080) );
  INV_X2 U1695 ( .A(n2136), .ZN(n2206) );
  OR2_X2 U1696 ( .A1(n2140), .A2(n2165), .ZN(n277) );
  OR2_X1 U1697 ( .A1(n1963), .A2(n856), .ZN(n2081) );
  BUF_X1 U1698 ( .A(n1957), .Z(n2148) );
  AND2_X2 U1699 ( .A1(n1809), .A2(n2062), .ZN(n2134) );
  XNOR2_X1 U1700 ( .A(n996), .B(n2082), .ZN(n973) );
  XNOR2_X1 U1701 ( .A(n994), .B(n1217), .ZN(n2082) );
  INV_X2 U1702 ( .A(n2249), .ZN(n2246) );
  CLKBUF_X1 U1703 ( .A(n1997), .Z(n2083) );
  INV_X2 U1704 ( .A(n2136), .ZN(n2205) );
  AND2_X2 U1705 ( .A1(n2101), .A2(n2071), .ZN(n2136) );
  XOR2_X1 U1706 ( .A(n1459), .B(n1370), .Z(n2084) );
  XOR2_X1 U1707 ( .A(n2084), .B(n1436), .Z(n957) );
  NAND2_X1 U1708 ( .A1(n1436), .A2(n1459), .ZN(n2085) );
  NAND2_X1 U1709 ( .A1(n1436), .A2(n1370), .ZN(n2086) );
  NAND2_X1 U1710 ( .A1(n1459), .A2(n1370), .ZN(n2087) );
  NAND3_X1 U1711 ( .A1(n2085), .A2(n2086), .A3(n2087), .ZN(n956) );
  AND2_X1 U1712 ( .A1(n857), .A2(n876), .ZN(n2088) );
  AND2_X2 U1713 ( .A1(n2014), .A2(n2099), .ZN(n2143) );
  INV_X2 U1714 ( .A(n2143), .ZN(n2217) );
  INV_X2 U1715 ( .A(n2135), .ZN(n2212) );
  AND2_X2 U1716 ( .A1(n2100), .A2(n2070), .ZN(n2135) );
  XOR2_X1 U1717 ( .A(n844), .B(n827), .Z(n2089) );
  XOR2_X1 U1718 ( .A(n1938), .B(n2089), .Z(n823) );
  NAND2_X1 U1719 ( .A1(n1937), .A2(n844), .ZN(n2090) );
  NAND2_X1 U1720 ( .A1(n842), .A2(n827), .ZN(n2091) );
  NAND2_X1 U1721 ( .A1(n844), .A2(n827), .ZN(n2092) );
  NAND3_X1 U1722 ( .A1(n2090), .A2(n2091), .A3(n2092), .ZN(n822) );
  INV_X1 U1723 ( .A(n491), .ZN(n2093) );
  NOR2_X1 U1724 ( .A1(n495), .A2(n502), .ZN(n489) );
  INV_X2 U1725 ( .A(n2132), .ZN(n2223) );
  AND2_X2 U1726 ( .A1(n1812), .A2(n1981), .ZN(n2139) );
  INV_X1 U1727 ( .A(n2141), .ZN(n2096) );
  XOR2_X1 U1728 ( .A(a[6]), .B(n1978), .Z(n2094) );
  OR2_X1 U1729 ( .A1(n1123), .A2(n1132), .ZN(n2097) );
  XOR2_X1 U1730 ( .A(a[12]), .B(a[13]), .Z(n2100) );
  NOR2_X1 U1731 ( .A1(n491), .A2(n467), .ZN(n465) );
  INV_X1 U1732 ( .A(n420), .ZN(n422) );
  INV_X1 U1733 ( .A(n400), .ZN(n398) );
  NAND2_X1 U1734 ( .A1(n426), .A2(n663), .ZN(n420) );
  NAND2_X1 U1735 ( .A1(n666), .A2(n481), .ZN(n315) );
  NAND2_X1 U1736 ( .A1(n668), .A2(n503), .ZN(n317) );
  NAND2_X1 U1737 ( .A1(n2081), .A2(n514), .ZN(n318) );
  NAND2_X1 U1738 ( .A1(n2040), .A2(n532), .ZN(n320) );
  OAI21_X1 U1739 ( .B1(n492), .B2(n467), .A(n468), .ZN(n466) );
  INV_X1 U1740 ( .A(n481), .ZN(n483) );
  INV_X1 U1741 ( .A(n503), .ZN(n501) );
  NOR2_X1 U1742 ( .A1(n402), .A2(n360), .ZN(n356) );
  AOI21_X1 U1743 ( .B1(n565), .B2(n561), .A(n562), .ZN(n560) );
  XOR2_X1 U1744 ( .A(n544), .B(n322), .Z(product[24]) );
  NAND2_X1 U1745 ( .A1(n2080), .A2(n543), .ZN(n322) );
  AOI21_X1 U1746 ( .B1(n565), .B2(n545), .A(n546), .ZN(n544) );
  XOR2_X1 U1747 ( .A(n551), .B(n323), .Z(product[23]) );
  NOR2_X1 U1748 ( .A1(n420), .A2(n402), .ZN(n400) );
  INV_X1 U1749 ( .A(n563), .ZN(n561) );
  INV_X1 U1750 ( .A(n564), .ZN(n562) );
  NAND2_X1 U1751 ( .A1(n663), .A2(n662), .ZN(n431) );
  AOI21_X1 U1752 ( .B1(n426), .B2(n445), .A(n427), .ZN(n421) );
  INV_X1 U1753 ( .A(n435), .ZN(n662) );
  NOR2_X1 U1754 ( .A1(n435), .A2(n428), .ZN(n426) );
  NAND2_X1 U1755 ( .A1(n2114), .A2(n461), .ZN(n313) );
  NAND2_X1 U1756 ( .A1(n2163), .A2(n496), .ZN(n316) );
  NOR2_X1 U1757 ( .A1(n384), .A2(n364), .ZN(n362) );
  NAND2_X1 U1758 ( .A1(n2108), .A2(n418), .ZN(n309) );
  NAND2_X1 U1759 ( .A1(n789), .A2(n804), .ZN(n481) );
  NAND2_X1 U1760 ( .A1(n657), .A2(n387), .ZN(n306) );
  INV_X1 U1761 ( .A(n384), .ZN(n657) );
  NAND2_X1 U1762 ( .A1(n661), .A2(n429), .ZN(n310) );
  NAND2_X1 U1763 ( .A1(n2111), .A2(n396), .ZN(n307) );
  INV_X1 U1764 ( .A(n438), .ZN(n663) );
  NOR2_X1 U1765 ( .A1(n1071), .A2(n1084), .ZN(n590) );
  AOI21_X1 U1766 ( .B1(n2110), .B2(n416), .A(n407), .ZN(n405) );
  INV_X1 U1767 ( .A(n409), .ZN(n407) );
  NAND2_X1 U1768 ( .A1(n821), .A2(n838), .ZN(n503) );
  INV_X1 U1769 ( .A(n418), .ZN(n416) );
  NOR2_X1 U1770 ( .A1(n420), .A2(n347), .ZN(n345) );
  NAND2_X1 U1771 ( .A1(n662), .A2(n436), .ZN(n311) );
  NAND2_X1 U1772 ( .A1(n2110), .A2(n409), .ZN(n308) );
  NAND2_X1 U1773 ( .A1(n422), .A2(n2108), .ZN(n411) );
  NAND2_X1 U1774 ( .A1(n2164), .A2(n378), .ZN(n305) );
  OR2_X1 U1775 ( .A1(n1021), .A2(n1038), .ZN(n2103) );
  AOI21_X1 U1776 ( .B1(n423), .B2(n2108), .A(n416), .ZN(n412) );
  AOI21_X1 U1777 ( .B1(n662), .B2(n445), .A(n434), .ZN(n432) );
  INV_X1 U1778 ( .A(n436), .ZN(n434) );
  INV_X1 U1779 ( .A(n378), .ZN(n376) );
  NAND2_X1 U1780 ( .A1(n2108), .A2(n2110), .ZN(n402) );
  INV_X1 U1781 ( .A(n396), .ZN(n394) );
  OR2_X1 U1782 ( .A1(n1055), .A2(n1070), .ZN(n2104) );
  OR2_X1 U1783 ( .A1(n1039), .A2(n1054), .ZN(n2105) );
  NAND2_X1 U1784 ( .A1(n362), .A2(n2111), .ZN(n360) );
  AND2_X1 U1785 ( .A1(n1039), .A2(n1054), .ZN(n2106) );
  AND2_X1 U1786 ( .A1(n1055), .A2(n1070), .ZN(n2107) );
  NOR2_X1 U1787 ( .A1(n1099), .A2(n1110), .ZN(n597) );
  OR2_X1 U1788 ( .A1(n717), .A2(n726), .ZN(n2108) );
  XNOR2_X1 U1789 ( .A(n2109), .B(n899), .ZN(n897) );
  XNOR2_X1 U1790 ( .A(n920), .B(n901), .ZN(n2109) );
  INV_X1 U1791 ( .A(n352), .ZN(n350) );
  NOR2_X1 U1792 ( .A1(n727), .A2(n736), .ZN(n428) );
  NOR2_X1 U1793 ( .A1(n695), .A2(n700), .ZN(n384) );
  NOR2_X1 U1794 ( .A1(n737), .A2(n748), .ZN(n435) );
  OR2_X1 U1795 ( .A1(n709), .A2(n716), .ZN(n2110) );
  OR2_X1 U1796 ( .A1(n694), .A2(n689), .ZN(n2164) );
  NAND2_X1 U1797 ( .A1(n2121), .A2(n341), .ZN(n302) );
  OR2_X1 U1798 ( .A1(n701), .A2(n708), .ZN(n2111) );
  NAND2_X1 U1799 ( .A1(n737), .A2(n748), .ZN(n436) );
  OAI21_X1 U1800 ( .B1(n405), .B2(n360), .A(n361), .ZN(n359) );
  AOI21_X1 U1801 ( .B1(n362), .B2(n394), .A(n363), .ZN(n361) );
  OAI21_X1 U1802 ( .B1(n364), .B2(n387), .A(n365), .ZN(n363) );
  AOI21_X1 U1803 ( .B1(n376), .B2(n2119), .A(n367), .ZN(n365) );
  AOI21_X1 U1804 ( .B1(n2112), .B2(n2115), .A(n2116), .ZN(n611) );
  NAND2_X1 U1805 ( .A1(n2117), .A2(n2112), .ZN(n610) );
  AOI21_X1 U1806 ( .B1(n625), .B2(n2124), .A(n2127), .ZN(n620) );
  OR2_X1 U1807 ( .A1(n1133), .A2(n1142), .ZN(n2112) );
  NAND2_X1 U1808 ( .A1(n2119), .A2(n369), .ZN(n304) );
  NAND2_X1 U1809 ( .A1(n2120), .A2(n352), .ZN(n303) );
  NAND2_X1 U1810 ( .A1(n695), .A2(n700), .ZN(n387) );
  NOR2_X1 U1811 ( .A1(n1085), .A2(n1098), .ZN(n592) );
  NAND2_X1 U1812 ( .A1(n727), .A2(n736), .ZN(n429) );
  OAI21_X1 U1813 ( .B1(n590), .B2(n593), .A(n591), .ZN(n589) );
  NAND2_X1 U1814 ( .A1(n1085), .A2(n1098), .ZN(n593) );
  OAI21_X1 U1815 ( .B1(n600), .B2(n597), .A(n598), .ZN(n596) );
  AOI21_X1 U1816 ( .B1(n2113), .B2(n2118), .A(n1940), .ZN(n600) );
  OR2_X1 U1817 ( .A1(n1111), .A2(n1122), .ZN(n2113) );
  OR2_X1 U1818 ( .A1(n761), .A2(n774), .ZN(n2114) );
  NAND2_X1 U1819 ( .A1(n701), .A2(n708), .ZN(n396) );
  NAND2_X1 U1820 ( .A1(n2164), .A2(n2119), .ZN(n364) );
  INV_X1 U1821 ( .A(n369), .ZN(n367) );
  AND2_X1 U1822 ( .A1(n1143), .A2(n1150), .ZN(n2115) );
  AND2_X1 U1823 ( .A1(n1133), .A2(n1142), .ZN(n2116) );
  NOR2_X1 U1824 ( .A1(n597), .A2(n599), .ZN(n595) );
  OR2_X1 U1825 ( .A1(n1143), .A2(n1150), .ZN(n2117) );
  AND2_X1 U1826 ( .A1(n1123), .A2(n1132), .ZN(n2118) );
  NAND2_X1 U1827 ( .A1(n1159), .A2(n1161), .ZN(n627) );
  AOI21_X1 U1828 ( .B1(n629), .B2(n635), .A(n630), .ZN(n628) );
  NOR2_X1 U1829 ( .A1(n1159), .A2(n1161), .ZN(n626) );
  NAND2_X1 U1830 ( .A1(n1175), .A2(n1178), .ZN(n637) );
  NOR2_X1 U1831 ( .A1(n1175), .A2(n1178), .ZN(n636) );
  AOI21_X1 U1832 ( .B1(n643), .B2(n2123), .A(n2126), .ZN(n638) );
  NOR2_X1 U1833 ( .A1(n1165), .A2(n1170), .ZN(n631) );
  OR2_X1 U1834 ( .A1(n685), .A2(n688), .ZN(n2119) );
  BUF_X1 U1835 ( .A(n2014), .Z(n2150) );
  NAND2_X1 U1836 ( .A1(n678), .A2(n677), .ZN(n335) );
  INV_X1 U1837 ( .A(n341), .ZN(n339) );
  OR2_X1 U1838 ( .A1(n681), .A2(n684), .ZN(n2120) );
  OAI21_X1 U1839 ( .B1(n631), .B2(n634), .A(n632), .ZN(n630) );
  OR2_X1 U1840 ( .A1(n679), .A2(n680), .ZN(n2121) );
  NAND2_X1 U1841 ( .A1(n681), .A2(n684), .ZN(n352) );
  NAND2_X1 U1842 ( .A1(n679), .A2(n680), .ZN(n341) );
  OR2_X1 U1843 ( .A1(n1457), .A2(n1480), .ZN(n2122) );
  OR2_X1 U1844 ( .A1(n1179), .A2(n1433), .ZN(n2123) );
  OR2_X1 U1845 ( .A1(n1151), .A2(n1158), .ZN(n2124) );
  AND2_X1 U1846 ( .A1(n1457), .A2(n1480), .ZN(n2125) );
  AND2_X1 U1847 ( .A1(n1179), .A2(n1433), .ZN(n2126) );
  AND2_X1 U1848 ( .A1(n1151), .A2(n1158), .ZN(n2127) );
  INV_X1 U1849 ( .A(n676), .ZN(n677) );
  OR2_X1 U1850 ( .A1(n1194), .A2(n676), .ZN(n2128) );
  AND2_X1 U1851 ( .A1(n1194), .A2(n676), .ZN(n2129) );
  NOR2_X1 U1852 ( .A1(n678), .A2(n677), .ZN(n334) );
  NAND2_X1 U1853 ( .A1(n2296), .A2(n2305), .ZN(n1756) );
  INV_X1 U1854 ( .A(n2271), .ZN(n2268) );
  INV_X1 U1855 ( .A(n2276), .ZN(n2273) );
  INV_X1 U1856 ( .A(n2250), .ZN(n2247) );
  INV_X1 U1857 ( .A(n2304), .ZN(n2301) );
  INV_X1 U1858 ( .A(n2288), .ZN(n2285) );
  INV_X1 U1859 ( .A(n2265), .ZN(n2263) );
  INV_X1 U1860 ( .A(n2255), .ZN(n2252) );
  INV_X1 U1861 ( .A(n2260), .ZN(n2257) );
  NOR2_X1 U1862 ( .A1(n2061), .A2(n2305), .ZN(n1433) );
  NOR2_X1 U1863 ( .A1(n2239), .A2(n2305), .ZN(n1457) );
  OAI22_X1 U1864 ( .A1(n2077), .A2(n1515), .B1(n2226), .B2(n1514), .ZN(n1225)
         );
  INV_X1 U1865 ( .A(n2161), .ZN(n2226) );
  INV_X1 U1866 ( .A(n2161), .ZN(n2225) );
  INV_X1 U1867 ( .A(n1507), .ZN(n2316) );
  INV_X1 U1868 ( .A(n682), .ZN(n683) );
  NAND2_X1 U1869 ( .A1(n2291), .A2(n2305), .ZN(n1731) );
  NOR2_X1 U1870 ( .A1(n2234), .A2(n2305), .ZN(n1385) );
  INV_X1 U1871 ( .A(n2141), .ZN(n2219) );
  INV_X1 U1872 ( .A(n1974), .ZN(n2222) );
  NOR2_X1 U1873 ( .A1(n2224), .A2(n2305), .ZN(n1217) );
  OAI21_X1 U1874 ( .B1(n646), .B2(n644), .A(n645), .ZN(n643) );
  NAND2_X1 U1875 ( .A1(n1181), .A2(n1192), .ZN(n645) );
  NOR2_X1 U1876 ( .A1(n1181), .A2(n1192), .ZN(n644) );
  AOI21_X1 U1877 ( .B1(n2122), .B2(n2130), .A(n2125), .ZN(n646) );
  INV_X1 U1878 ( .A(n1632), .ZN(n2311) );
  INV_X1 U1879 ( .A(n1532), .ZN(n2315) );
  NOR2_X1 U1880 ( .A1(n2235), .A2(n2305), .ZN(n1409) );
  NAND2_X1 U1881 ( .A1(n1960), .A2(n2305), .ZN(n1606) );
  NAND2_X1 U1882 ( .A1(n2273), .A2(n2305), .ZN(n1656) );
  NAND2_X1 U1883 ( .A1(n2252), .A2(n2305), .ZN(n1556) );
  NAND2_X1 U1884 ( .A1(n2268), .A2(n2305), .ZN(n1631) );
  NAND2_X1 U1885 ( .A1(n2285), .A2(n2305), .ZN(n1706) );
  NAND2_X1 U1886 ( .A1(n1972), .A2(n2305), .ZN(n1531) );
  NAND2_X1 U1887 ( .A1(n2279), .A2(n2305), .ZN(n1681) );
  NAND2_X1 U1888 ( .A1(n2258), .A2(n2305), .ZN(n1581) );
  NAND2_X1 U1889 ( .A1(n2301), .A2(n2305), .ZN(n1781) );
  INV_X1 U1890 ( .A(n1707), .ZN(n2308) );
  OAI22_X1 U1891 ( .A1(n2077), .A2(n1511), .B1(n2226), .B2(n1510), .ZN(n1221)
         );
  INV_X1 U1892 ( .A(n1682), .ZN(n2309) );
  OAI21_X1 U1893 ( .B1(n2221), .B2(n2005), .A(n2307), .ZN(n1434) );
  NOR2_X1 U1894 ( .A1(n2229), .A2(n2305), .ZN(n1313) );
  INV_X1 U1895 ( .A(n692), .ZN(n693) );
  OAI22_X1 U1896 ( .A1(n2077), .A2(n1509), .B1(n2225), .B2(n1508), .ZN(n1219)
         );
  OAI22_X1 U1897 ( .A1(n2077), .A2(n1517), .B1(n2225), .B2(n1516), .ZN(n1227)
         );
  NOR2_X1 U1898 ( .A1(n2232), .A2(n2305), .ZN(n1361) );
  NOR2_X1 U1899 ( .A1(n2227), .A2(n2305), .ZN(n1265) );
  NOR2_X1 U1900 ( .A1(n2225), .A2(n2305), .ZN(n1241) );
  OAI22_X1 U1901 ( .A1(n2077), .A2(n1513), .B1(n2226), .B2(n1512), .ZN(n1223)
         );
  INV_X1 U1902 ( .A(n802), .ZN(n803) );
  NOR2_X1 U1903 ( .A1(n1934), .A2(n2305), .ZN(n1337) );
  NOR2_X1 U1904 ( .A1(n2228), .A2(n2305), .ZN(n1289) );
  INV_X1 U1905 ( .A(n1557), .ZN(n2314) );
  INV_X1 U1906 ( .A(n1607), .ZN(n2312) );
  INV_X1 U1907 ( .A(n772), .ZN(n773) );
  INV_X1 U1908 ( .A(n1732), .ZN(n2307) );
  INV_X1 U1909 ( .A(n724), .ZN(n725) );
  CLKBUF_X1 U1910 ( .A(n251), .Z(n2241) );
  AND2_X1 U1911 ( .A1(n1193), .A2(n1481), .ZN(n2130) );
  INV_X1 U1912 ( .A(n1657), .ZN(n2310) );
  INV_X1 U1913 ( .A(n1582), .ZN(n2313) );
  INV_X1 U1914 ( .A(n1482), .ZN(n2317) );
  XNOR2_X1 U1915 ( .A(n2280), .B(b[0]), .ZN(n1680) );
  XNOR2_X1 U1916 ( .A(n2274), .B(b[0]), .ZN(n1655) );
  XNOR2_X1 U1917 ( .A(n2253), .B(b[0]), .ZN(n1555) );
  XNOR2_X1 U1918 ( .A(n2262), .B(b[0]), .ZN(n1605) );
  XNOR2_X1 U1919 ( .A(n2259), .B(b[0]), .ZN(n1580) );
  XNOR2_X1 U1920 ( .A(n2296), .B(b[22]), .ZN(n1733) );
  XNOR2_X1 U1921 ( .A(n1973), .B(b[14]), .ZN(n1516) );
  XNOR2_X1 U1922 ( .A(n1973), .B(b[18]), .ZN(n1512) );
  XNOR2_X1 U1923 ( .A(n2248), .B(b[22]), .ZN(n1508) );
  XNOR2_X1 U1924 ( .A(n2248), .B(b[16]), .ZN(n1514) );
  XNOR2_X1 U1925 ( .A(n1972), .B(b[20]), .ZN(n1510) );
  XNOR2_X1 U1926 ( .A(n2301), .B(b[18]), .ZN(n1762) );
  XNOR2_X1 U1927 ( .A(n2302), .B(b[22]), .ZN(n1758) );
  XNOR2_X1 U1928 ( .A(n2301), .B(b[14]), .ZN(n1766) );
  XNOR2_X1 U1929 ( .A(n2301), .B(b[10]), .ZN(n1770) );
  XNOR2_X1 U1930 ( .A(n2302), .B(b[16]), .ZN(n1764) );
  XNOR2_X1 U1931 ( .A(n2302), .B(b[20]), .ZN(n1760) );
  XNOR2_X1 U1932 ( .A(n2301), .B(b[6]), .ZN(n1774) );
  XNOR2_X1 U1933 ( .A(n2301), .B(b[4]), .ZN(n1776) );
  XNOR2_X1 U1934 ( .A(n2301), .B(b[8]), .ZN(n1772) );
  XNOR2_X1 U1935 ( .A(n2273), .B(b[10]), .ZN(n1645) );
  XNOR2_X1 U1936 ( .A(n2252), .B(b[6]), .ZN(n1549) );
  XNOR2_X1 U1937 ( .A(n2273), .B(b[14]), .ZN(n1641) );
  XNOR2_X1 U1938 ( .A(n2258), .B(b[8]), .ZN(n1572) );
  XNOR2_X1 U1939 ( .A(n2247), .B(b[4]), .ZN(n1526) );
  XNOR2_X1 U1940 ( .A(n2286), .B(b[22]), .ZN(n1683) );
  XNOR2_X1 U1941 ( .A(n2252), .B(b[4]), .ZN(n1551) );
  XNOR2_X1 U1942 ( .A(n2279), .B(b[14]), .ZN(n1666) );
  XNOR2_X1 U1943 ( .A(n2264), .B(b[6]), .ZN(n1599) );
  XNOR2_X1 U1944 ( .A(n2292), .B(b[16]), .ZN(n1714) );
  XNOR2_X1 U1945 ( .A(n2286), .B(b[16]), .ZN(n1689) );
  XNOR2_X1 U1946 ( .A(n2258), .B(b[4]), .ZN(n1576) );
  XNOR2_X1 U1947 ( .A(n1960), .B(b[10]), .ZN(n1595) );
  XNOR2_X1 U1948 ( .A(n2292), .B(b[20]), .ZN(n1710) );
  XNOR2_X1 U1949 ( .A(n2268), .B(b[6]), .ZN(n1624) );
  XNOR2_X1 U1950 ( .A(n2291), .B(b[18]), .ZN(n1712) );
  XNOR2_X1 U1951 ( .A(n2296), .B(b[20]), .ZN(n1735) );
  XNOR2_X1 U1952 ( .A(n2264), .B(b[8]), .ZN(n1597) );
  XNOR2_X1 U1953 ( .A(n2258), .B(b[6]), .ZN(n1574) );
  XNOR2_X1 U1954 ( .A(n2269), .B(b[14]), .ZN(n1616) );
  XNOR2_X1 U1955 ( .A(n2285), .B(b[8]), .ZN(n1697) );
  XNOR2_X1 U1956 ( .A(n2296), .B(b[14]), .ZN(n1741) );
  XNOR2_X1 U1957 ( .A(n1992), .B(b[8]), .ZN(n1622) );
  XNOR2_X1 U1958 ( .A(n2291), .B(b[6]), .ZN(n1724) );
  XNOR2_X1 U1959 ( .A(n2248), .B(b[6]), .ZN(n1524) );
  XNOR2_X1 U1960 ( .A(n2273), .B(b[4]), .ZN(n1651) );
  XNOR2_X1 U1961 ( .A(n2273), .B(b[6]), .ZN(n1649) );
  XNOR2_X1 U1962 ( .A(n2279), .B(b[18]), .ZN(n1662) );
  XNOR2_X1 U1963 ( .A(n2280), .B(b[22]), .ZN(n1658) );
  XNOR2_X1 U1964 ( .A(n1968), .B(b[10]), .ZN(n1745) );
  XNOR2_X1 U1965 ( .A(n2274), .B(b[22]), .ZN(n1633) );
  XNOR2_X1 U1966 ( .A(n2252), .B(b[8]), .ZN(n1547) );
  XNOR2_X1 U1967 ( .A(n2285), .B(b[6]), .ZN(n1699) );
  XNOR2_X1 U1968 ( .A(n2292), .B(b[22]), .ZN(n1708) );
  XNOR2_X1 U1969 ( .A(n2279), .B(b[6]), .ZN(n1674) );
  XNOR2_X1 U1970 ( .A(n1992), .B(b[16]), .ZN(n1614) );
  XNOR2_X1 U1971 ( .A(n2285), .B(b[14]), .ZN(n1691) );
  XNOR2_X1 U1972 ( .A(n2269), .B(b[10]), .ZN(n1620) );
  XNOR2_X1 U1973 ( .A(n2252), .B(b[10]), .ZN(n1545) );
  XNOR2_X1 U1974 ( .A(n2273), .B(b[18]), .ZN(n1637) );
  XNOR2_X1 U1975 ( .A(n1991), .B(b[22]), .ZN(n1608) );
  XNOR2_X1 U1976 ( .A(n2285), .B(b[10]), .ZN(n1695) );
  XNOR2_X1 U1977 ( .A(n2274), .B(b[16]), .ZN(n1639) );
  XNOR2_X1 U1978 ( .A(n2269), .B(b[4]), .ZN(n1626) );
  XNOR2_X1 U1979 ( .A(n1968), .B(b[18]), .ZN(n1737) );
  XNOR2_X1 U1980 ( .A(n2279), .B(b[8]), .ZN(n1672) );
  XNOR2_X1 U1981 ( .A(n2279), .B(b[4]), .ZN(n1676) );
  XNOR2_X1 U1982 ( .A(n2280), .B(b[16]), .ZN(n1664) );
  XNOR2_X1 U1983 ( .A(n2291), .B(b[8]), .ZN(n1722) );
  XNOR2_X1 U1984 ( .A(n1968), .B(b[4]), .ZN(n1751) );
  XNOR2_X1 U1985 ( .A(n1991), .B(b[20]), .ZN(n1610) );
  XNOR2_X1 U1986 ( .A(n2279), .B(b[10]), .ZN(n1670) );
  XNOR2_X1 U1987 ( .A(n1960), .B(b[4]), .ZN(n1601) );
  XNOR2_X1 U1988 ( .A(n2259), .B(b[16]), .ZN(n1564) );
  XNOR2_X1 U1989 ( .A(n2296), .B(b[16]), .ZN(n1739) );
  XNOR2_X1 U1990 ( .A(n2273), .B(b[8]), .ZN(n1647) );
  XNOR2_X1 U1991 ( .A(n1960), .B(b[14]), .ZN(n1591) );
  XNOR2_X1 U1992 ( .A(n1972), .B(b[8]), .ZN(n1522) );
  XNOR2_X1 U1993 ( .A(n2285), .B(b[4]), .ZN(n1701) );
  XNOR2_X1 U1994 ( .A(n2252), .B(b[14]), .ZN(n1541) );
  XNOR2_X1 U1995 ( .A(n2253), .B(b[16]), .ZN(n1539) );
  XNOR2_X1 U1996 ( .A(n2264), .B(b[20]), .ZN(n1585) );
  XNOR2_X1 U1997 ( .A(n2259), .B(b[22]), .ZN(n1558) );
  XNOR2_X1 U1998 ( .A(n2285), .B(b[18]), .ZN(n1687) );
  XNOR2_X1 U1999 ( .A(n2252), .B(b[18]), .ZN(n1537) );
  XNOR2_X1 U2000 ( .A(n2263), .B(b[18]), .ZN(n1587) );
  XNOR2_X1 U2001 ( .A(n2286), .B(b[20]), .ZN(n1685) );
  XNOR2_X1 U2002 ( .A(n2291), .B(b[14]), .ZN(n1716) );
  XNOR2_X1 U2003 ( .A(n2258), .B(b[10]), .ZN(n1570) );
  XNOR2_X1 U2004 ( .A(n1968), .B(b[8]), .ZN(n1747) );
  XNOR2_X1 U2005 ( .A(n2291), .B(b[4]), .ZN(n1726) );
  XNOR2_X1 U2006 ( .A(n2268), .B(b[18]), .ZN(n1612) );
  XNOR2_X1 U2007 ( .A(n2296), .B(b[6]), .ZN(n1749) );
  XNOR2_X1 U2008 ( .A(n2274), .B(b[20]), .ZN(n1635) );
  XNOR2_X1 U2009 ( .A(n2258), .B(b[18]), .ZN(n1562) );
  XNOR2_X1 U2010 ( .A(n1961), .B(b[16]), .ZN(n1589) );
  XNOR2_X1 U2011 ( .A(n2248), .B(b[10]), .ZN(n1520) );
  XNOR2_X1 U2012 ( .A(n1960), .B(b[22]), .ZN(n1583) );
  XNOR2_X1 U2013 ( .A(n2253), .B(b[22]), .ZN(n1533) );
  XNOR2_X1 U2014 ( .A(n2258), .B(b[14]), .ZN(n1566) );
  XNOR2_X1 U2015 ( .A(n2280), .B(b[20]), .ZN(n1660) );
  XNOR2_X1 U2016 ( .A(n2259), .B(b[20]), .ZN(n1560) );
  XNOR2_X1 U2017 ( .A(n2291), .B(b[10]), .ZN(n1720) );
  XNOR2_X1 U2018 ( .A(n2253), .B(b[20]), .ZN(n1535) );
  XNOR2_X1 U2019 ( .A(n1972), .B(b[0]), .ZN(n1530) );
  XNOR2_X1 U2020 ( .A(n2301), .B(b[2]), .ZN(n1778) );
  XNOR2_X1 U2021 ( .A(n2301), .B(b[12]), .ZN(n1768) );
  XNOR2_X1 U2022 ( .A(n2268), .B(b[2]), .ZN(n1628) );
  XNOR2_X1 U2023 ( .A(n2285), .B(b[12]), .ZN(n1693) );
  XNOR2_X1 U2024 ( .A(n2273), .B(b[12]), .ZN(n1643) );
  XNOR2_X1 U2025 ( .A(n1991), .B(b[12]), .ZN(n1618) );
  XNOR2_X1 U2026 ( .A(n2279), .B(b[2]), .ZN(n1678) );
  XNOR2_X1 U2027 ( .A(n2247), .B(b[2]), .ZN(n1528) );
  XNOR2_X1 U2028 ( .A(n2258), .B(b[12]), .ZN(n1568) );
  XNOR2_X1 U2029 ( .A(n2263), .B(b[2]), .ZN(n1603) );
  XNOR2_X1 U2030 ( .A(n1968), .B(b[12]), .ZN(n1743) );
  XNOR2_X1 U2031 ( .A(n2285), .B(b[2]), .ZN(n1703) );
  XNOR2_X1 U2032 ( .A(n1960), .B(b[12]), .ZN(n1593) );
  XNOR2_X1 U2033 ( .A(n2273), .B(b[2]), .ZN(n1653) );
  XNOR2_X1 U2034 ( .A(n2258), .B(b[2]), .ZN(n1578) );
  XNOR2_X1 U2035 ( .A(n2291), .B(b[12]), .ZN(n1718) );
  XNOR2_X1 U2036 ( .A(n2291), .B(b[2]), .ZN(n1728) );
  XNOR2_X1 U2037 ( .A(n2252), .B(b[12]), .ZN(n1543) );
  XNOR2_X1 U2038 ( .A(n1968), .B(b[2]), .ZN(n1753) );
  XNOR2_X1 U2039 ( .A(n1973), .B(b[12]), .ZN(n1518) );
  XNOR2_X1 U2040 ( .A(n1992), .B(b[0]), .ZN(n1630) );
  XNOR2_X1 U2041 ( .A(n2286), .B(b[0]), .ZN(n1705) );
  XNOR2_X1 U2042 ( .A(n2292), .B(b[0]), .ZN(n1730) );
  AND2_X1 U2043 ( .A1(n1817), .A2(n2240), .ZN(n2132) );
  XNOR2_X1 U2044 ( .A(b[23]), .B(n1988), .ZN(n1607) );
  XNOR2_X1 U2045 ( .A(b[23]), .B(n2257), .ZN(n1557) );
  XNOR2_X1 U2046 ( .A(b[23]), .B(n2251), .ZN(n1532) );
  XNOR2_X1 U2047 ( .A(b[7]), .B(n2251), .ZN(n1548) );
  XNOR2_X1 U2048 ( .A(b[1]), .B(n2251), .ZN(n1554) );
  XNOR2_X1 U2049 ( .A(b[5]), .B(n2251), .ZN(n1550) );
  XNOR2_X1 U2050 ( .A(b[7]), .B(n1988), .ZN(n1623) );
  XNOR2_X1 U2051 ( .A(b[9]), .B(n2257), .ZN(n1571) );
  XNOR2_X1 U2052 ( .A(b[1]), .B(n2242), .ZN(n1504) );
  XNOR2_X1 U2053 ( .A(b[3]), .B(n2242), .ZN(n1502) );
  XNOR2_X1 U2054 ( .A(b[9]), .B(n1989), .ZN(n1621) );
  XNOR2_X1 U2055 ( .A(b[9]), .B(n2251), .ZN(n1546) );
  XNOR2_X1 U2056 ( .A(b[7]), .B(n2242), .ZN(n1498) );
  XNOR2_X1 U2057 ( .A(b[3]), .B(n2257), .ZN(n1577) );
  XNOR2_X1 U2058 ( .A(b[1]), .B(n1989), .ZN(n1629) );
  XNOR2_X1 U2059 ( .A(b[5]), .B(n2242), .ZN(n1500) );
  XNOR2_X1 U2060 ( .A(b[7]), .B(n2257), .ZN(n1573) );
  XNOR2_X1 U2061 ( .A(b[5]), .B(n2257), .ZN(n1575) );
  XNOR2_X1 U2062 ( .A(b[9]), .B(n2242), .ZN(n1496) );
  XNOR2_X1 U2063 ( .A(b[5]), .B(n2267), .ZN(n1625) );
  XNOR2_X1 U2064 ( .A(b[1]), .B(n2257), .ZN(n1579) );
  XNOR2_X1 U2065 ( .A(b[3]), .B(n2272), .ZN(n1652) );
  NOR2_X1 U2066 ( .A1(n2138), .A2(n1985), .ZN(n2137) );
  XNOR2_X1 U2067 ( .A(b[13]), .B(n2242), .ZN(n1492) );
  XNOR2_X1 U2068 ( .A(b[11]), .B(n2242), .ZN(n1494) );
  XNOR2_X1 U2069 ( .A(b[17]), .B(n2242), .ZN(n1488) );
  XNOR2_X1 U2070 ( .A(b[15]), .B(n2242), .ZN(n1490) );
  XNOR2_X1 U2071 ( .A(b[19]), .B(n2242), .ZN(n1486) );
  XNOR2_X1 U2072 ( .A(b[21]), .B(n2242), .ZN(n1484) );
  XNOR2_X1 U2073 ( .A(n2302), .B(b[0]), .ZN(n1780) );
  OAI21_X1 U2074 ( .B1(a[0]), .B2(n1974), .A(n2306), .ZN(n1458) );
  INV_X1 U2075 ( .A(n1757), .ZN(n2306) );
  INV_X1 U2076 ( .A(a[23]), .ZN(n2244) );
  XNOR2_X1 U2077 ( .A(n2296), .B(b[0]), .ZN(n1755) );
  INV_X1 U2078 ( .A(a[0]), .ZN(n251) );
  XNOR2_X1 U2079 ( .A(b[23]), .B(n2242), .ZN(n1482) );
  INV_X1 U2080 ( .A(n2244), .ZN(n2243) );
  INV_X1 U2081 ( .A(n2287), .ZN(n2284) );
  INV_X1 U2082 ( .A(n2133), .ZN(n2229) );
  INV_X1 U2083 ( .A(n277), .ZN(n2221) );
  OAI21_X1 U2084 ( .B1(n2142), .B2(n2169), .A(n2308), .ZN(n1410) );
  INV_X1 U2085 ( .A(n2131), .ZN(n2157) );
  INV_X1 U2086 ( .A(n2131), .ZN(n2156) );
  OAI21_X1 U2087 ( .B1(n2136), .B2(n1980), .A(n2317), .ZN(n1194) );
  OAI22_X1 U2088 ( .A1(n2206), .A2(n1484), .B1(n2147), .B2(n1483), .ZN(n1195)
         );
  OAI22_X1 U2089 ( .A1(n2206), .A2(n1488), .B1(n2147), .B2(n1487), .ZN(n1199)
         );
  OAI22_X1 U2090 ( .A1(n2206), .A2(n1486), .B1(n2147), .B2(n1485), .ZN(n1197)
         );
  OAI22_X1 U2091 ( .A1(n2206), .A2(n1490), .B1(n2224), .B2(n1489), .ZN(n1201)
         );
  OAI22_X1 U2092 ( .A1(n2206), .A2(n1492), .B1(n2224), .B2(n1491), .ZN(n1203)
         );
  INV_X1 U2093 ( .A(n1980), .ZN(n2224) );
  CLKBUF_X1 U2094 ( .A(n505), .Z(n2158) );
  INV_X1 U2095 ( .A(n2035), .ZN(n2159) );
  OAI21_X1 U2096 ( .B1(n2135), .B2(n2170), .A(n2312), .ZN(n1314) );
  OR2_X1 U2097 ( .A1(n857), .A2(n876), .ZN(n2160) );
  OAI21_X1 U2098 ( .B1(n2143), .B2(n2175), .A(n2310), .ZN(n1362) );
  AOI21_X1 U2099 ( .B1(n1952), .B2(n567), .A(n2069), .ZN(n2162) );
  OAI21_X1 U2100 ( .B1(n2131), .B2(n2176), .A(n2315), .ZN(n1242) );
  OAI22_X1 U2101 ( .A1(n2157), .A2(n1536), .B1(n2227), .B2(n1535), .ZN(n1245)
         );
  OAI22_X1 U2102 ( .A1(n2208), .A2(n1534), .B1(n2227), .B2(n1533), .ZN(n1243)
         );
  OAI22_X1 U2103 ( .A1(n2156), .A2(n1538), .B1(n2227), .B2(n1537), .ZN(n1247)
         );
  OAI22_X1 U2104 ( .A1(n2156), .A2(n1540), .B1(n2227), .B2(n1539), .ZN(n1249)
         );
  OAI22_X1 U2105 ( .A1(n2208), .A2(n1542), .B1(n2227), .B2(n1541), .ZN(n1251)
         );
  OR2_X1 U2106 ( .A1(n2016), .A2(n820), .ZN(n2163) );
  OAI21_X1 U2107 ( .B1(n628), .B2(n626), .A(n627), .ZN(n625) );
  XNOR2_X1 U2108 ( .A(b[9]), .B(n2278), .ZN(n1671) );
  XNOR2_X1 U2109 ( .A(b[1]), .B(n2278), .ZN(n1679) );
  XNOR2_X1 U2110 ( .A(b[7]), .B(n2278), .ZN(n1673) );
  XNOR2_X1 U2111 ( .A(b[5]), .B(n2278), .ZN(n1675) );
  XNOR2_X1 U2112 ( .A(b[3]), .B(n2278), .ZN(n1677) );
  XNOR2_X1 U2113 ( .A(b[23]), .B(n2278), .ZN(n1657) );
  XNOR2_X1 U2114 ( .A(b[23]), .B(n2272), .ZN(n1632) );
  XNOR2_X1 U2115 ( .A(b[9]), .B(n2272), .ZN(n1646) );
  XNOR2_X1 U2116 ( .A(b[1]), .B(n2272), .ZN(n1654) );
  XNOR2_X1 U2117 ( .A(b[5]), .B(n2272), .ZN(n1650) );
  XNOR2_X1 U2118 ( .A(b[7]), .B(n2272), .ZN(n1648) );
  XNOR2_X1 U2119 ( .A(b[9]), .B(n2289), .ZN(n1721) );
  XNOR2_X1 U2120 ( .A(b[5]), .B(n2289), .ZN(n1725) );
  XNOR2_X1 U2121 ( .A(b[1]), .B(n2289), .ZN(n1729) );
  XNOR2_X1 U2122 ( .A(b[3]), .B(n2289), .ZN(n1727) );
  XNOR2_X1 U2123 ( .A(b[7]), .B(n2289), .ZN(n1723) );
  XNOR2_X1 U2124 ( .A(b[23]), .B(n2289), .ZN(n1707) );
  NAND2_X1 U2125 ( .A1(n1954), .A2(n550), .ZN(n323) );
  INV_X1 U2126 ( .A(n2131), .ZN(n2207) );
  OAI22_X1 U2127 ( .A1(n1998), .A2(n2303), .B1(n1781), .B2(n2240), .ZN(n1193)
         );
  OAI22_X1 U2128 ( .A1(n2223), .A2(n1764), .B1(n1763), .B2(n2240), .ZN(n1465)
         );
  OAI22_X1 U2129 ( .A1(n2222), .A2(n1768), .B1(n1767), .B2(n2240), .ZN(n1469)
         );
  OAI22_X1 U2130 ( .A1(n2222), .A2(n1760), .B1(n1759), .B2(n2241), .ZN(n1461)
         );
  OAI22_X1 U2131 ( .A1(n2223), .A2(n1763), .B1(n1762), .B2(n2240), .ZN(n1464)
         );
  OAI22_X1 U2132 ( .A1(n2223), .A2(n1767), .B1(n1766), .B2(n2240), .ZN(n1468)
         );
  OAI22_X1 U2133 ( .A1(n1999), .A2(n1761), .B1(n1760), .B2(n2241), .ZN(n1462)
         );
  OAI22_X1 U2134 ( .A1(n1998), .A2(n1759), .B1(n1758), .B2(n2241), .ZN(n1460)
         );
  OAI22_X1 U2135 ( .A1(n2223), .A2(n1766), .B1(n1765), .B2(n2240), .ZN(n1467)
         );
  OAI22_X1 U2136 ( .A1(n1999), .A2(n1765), .B1(n1764), .B2(n2240), .ZN(n1466)
         );
  OAI22_X1 U2137 ( .A1(n1999), .A2(n1758), .B1(n1757), .B2(n2241), .ZN(n1459)
         );
  OAI22_X1 U2138 ( .A1(n1999), .A2(n1762), .B1(n1761), .B2(n2241), .ZN(n1463)
         );
  NAND2_X1 U2139 ( .A1(n1099), .A2(n1110), .ZN(n598) );
  OAI21_X1 U2140 ( .B1(n2141), .B2(n2094), .A(n2309), .ZN(n1386) );
  OAI22_X1 U2141 ( .A1(n2004), .A2(n1695), .B1(n1694), .B2(n2235), .ZN(n1398)
         );
  OAI22_X1 U2142 ( .A1(n2004), .A2(n1701), .B1(n1700), .B2(n2235), .ZN(n1404)
         );
  OAI22_X1 U2143 ( .A1(n2218), .A2(n1704), .B1(n2235), .B2(n1703), .ZN(n1407)
         );
  OAI22_X1 U2144 ( .A1(n2096), .A2(n1694), .B1(n2236), .B2(n1693), .ZN(n1397)
         );
  OAI22_X1 U2145 ( .A1(n2096), .A2(n1702), .B1(n2235), .B2(n1701), .ZN(n1405)
         );
  OAI22_X1 U2146 ( .A1(n2096), .A2(n1698), .B1(n2235), .B2(n1697), .ZN(n1401)
         );
  OAI22_X1 U2147 ( .A1(n2004), .A2(n1700), .B1(n2235), .B2(n1699), .ZN(n1403)
         );
  OAI22_X1 U2148 ( .A1(n2095), .A2(n1696), .B1(n1986), .B2(n1695), .ZN(n1399)
         );
  OAI22_X1 U2149 ( .A1(n2095), .A2(n1697), .B1(n1696), .B2(n2235), .ZN(n1400)
         );
  OAI22_X1 U2150 ( .A1(n2218), .A2(n1699), .B1(n1698), .B2(n2235), .ZN(n1402)
         );
  INV_X1 U2151 ( .A(n2094), .ZN(n2235) );
  NOR2_X1 U2152 ( .A1(n531), .A2(n534), .ZN(n525) );
  XNOR2_X1 U2153 ( .A(b[23]), .B(n2263), .ZN(n1582) );
  XNOR2_X1 U2154 ( .A(b[3]), .B(n2263), .ZN(n1602) );
  XNOR2_X1 U2155 ( .A(b[5]), .B(n2262), .ZN(n1600) );
  XNOR2_X1 U2156 ( .A(b[9]), .B(n2263), .ZN(n1596) );
  XNOR2_X1 U2157 ( .A(b[7]), .B(n1961), .ZN(n1598) );
  XNOR2_X1 U2158 ( .A(b[1]), .B(n2262), .ZN(n1604) );
  XNOR2_X1 U2159 ( .A(b[23]), .B(n2246), .ZN(n1507) );
  XNOR2_X1 U2160 ( .A(b[9]), .B(n2246), .ZN(n1521) );
  XNOR2_X1 U2161 ( .A(b[1]), .B(n2246), .ZN(n1529) );
  XNOR2_X1 U2162 ( .A(b[7]), .B(n2246), .ZN(n1523) );
  XNOR2_X1 U2163 ( .A(b[5]), .B(n2246), .ZN(n1525) );
  XNOR2_X1 U2164 ( .A(b[3]), .B(n2246), .ZN(n1527) );
  NOR2_X1 U2165 ( .A1(n896), .A2(n877), .ZN(n531) );
  XNOR2_X1 U2166 ( .A(n2152), .B(b[22]), .ZN(n1483) );
  XNOR2_X1 U2167 ( .A(n2152), .B(b[20]), .ZN(n1485) );
  XNOR2_X1 U2168 ( .A(n2152), .B(b[18]), .ZN(n1487) );
  NAND2_X1 U2169 ( .A1(n2152), .A2(n2305), .ZN(n1506) );
  XNOR2_X1 U2170 ( .A(n2152), .B(b[16]), .ZN(n1489) );
  XNOR2_X1 U2171 ( .A(n2152), .B(b[12]), .ZN(n1493) );
  XNOR2_X1 U2172 ( .A(n2152), .B(b[10]), .ZN(n1495) );
  XNOR2_X1 U2173 ( .A(n2152), .B(b[14]), .ZN(n1491) );
  XNOR2_X1 U2174 ( .A(n2152), .B(b[4]), .ZN(n1501) );
  XNOR2_X1 U2175 ( .A(n2152), .B(b[8]), .ZN(n1497) );
  XNOR2_X1 U2176 ( .A(n2152), .B(b[6]), .ZN(n1499) );
  XNOR2_X1 U2177 ( .A(n2152), .B(b[2]), .ZN(n1503) );
  XNOR2_X1 U2178 ( .A(n2152), .B(b[0]), .ZN(n1505) );
  XNOR2_X1 U2179 ( .A(b[7]), .B(n1968), .ZN(n1748) );
  XNOR2_X1 U2180 ( .A(b[3]), .B(n1968), .ZN(n1752) );
  XNOR2_X1 U2181 ( .A(b[9]), .B(n1968), .ZN(n1746) );
  XNOR2_X1 U2182 ( .A(b[5]), .B(n1968), .ZN(n1750) );
  XNOR2_X1 U2183 ( .A(b[1]), .B(n1968), .ZN(n1754) );
  XNOR2_X1 U2184 ( .A(b[23]), .B(n2295), .ZN(n1732) );
  NOR2_X1 U2185 ( .A1(n983), .A2(n1002), .ZN(n563) );
  NAND2_X1 U2186 ( .A1(n1165), .A2(n1170), .ZN(n632) );
  NAND2_X1 U2187 ( .A1(n2160), .A2(n521), .ZN(n319) );
  NAND2_X1 U2188 ( .A1(n857), .A2(n876), .ZN(n521) );
  OAI21_X1 U2189 ( .B1(n1984), .B2(n521), .A(n514), .ZN(n2166) );
  OAI21_X1 U2190 ( .B1(n2137), .B2(n1985), .A(n2313), .ZN(n1290) );
  NOR2_X1 U2191 ( .A1(n520), .A2(n513), .ZN(n2168) );
  XNOR2_X1 U2192 ( .A(b[3]), .B(n2286), .ZN(n1702) );
  XNOR2_X1 U2193 ( .A(b[1]), .B(n2284), .ZN(n1704) );
  XNOR2_X1 U2194 ( .A(b[5]), .B(n2284), .ZN(n1700) );
  XNOR2_X1 U2195 ( .A(b[9]), .B(n2284), .ZN(n1696) );
  XNOR2_X1 U2196 ( .A(b[7]), .B(n2286), .ZN(n1698) );
  XNOR2_X1 U2197 ( .A(b[23]), .B(n2284), .ZN(n1682) );
  NOR2_X1 U2198 ( .A1(n805), .A2(n820), .ZN(n495) );
  OAI21_X1 U2199 ( .B1(n2134), .B2(n2167), .A(n2314), .ZN(n1266) );
  NAND2_X1 U2200 ( .A1(n899), .A2(n920), .ZN(n2171) );
  NAND2_X1 U2201 ( .A1(n899), .A2(n901), .ZN(n2172) );
  NAND2_X1 U2202 ( .A1(n920), .A2(n901), .ZN(n2173) );
  NAND3_X1 U2203 ( .A1(n2171), .A2(n2172), .A3(n2173), .ZN(n896) );
  AND2_X1 U2204 ( .A1(n1932), .A2(n2168), .ZN(n2174) );
  AOI21_X1 U2205 ( .B1(n359), .B2(n2120), .A(n350), .ZN(n348) );
  INV_X1 U2206 ( .A(n2287), .ZN(n2283) );
  INV_X1 U2207 ( .A(n2260), .ZN(n2256) );
  INV_X1 U2208 ( .A(n502), .ZN(n668) );
  NOR2_X1 U2209 ( .A1(n821), .A2(n838), .ZN(n502) );
  OAI21_X1 U2210 ( .B1(n2144), .B2(n2058), .A(n2316), .ZN(n1218) );
  NAND2_X1 U2211 ( .A1(n877), .A2(n896), .ZN(n532) );
  AOI21_X1 U2212 ( .B1(n581), .B2(n567), .A(n568), .ZN(n566) );
  OAI22_X1 U2213 ( .A1(n2222), .A2(n1772), .B1(n1771), .B2(n2240), .ZN(n1473)
         );
  OAI22_X1 U2214 ( .A1(n2222), .A2(n1780), .B1(n1779), .B2(n2240), .ZN(n1481)
         );
  OAI22_X1 U2215 ( .A1(n1998), .A2(n1776), .B1(n1775), .B2(n2240), .ZN(n1477)
         );
  OAI22_X1 U2216 ( .A1(n2223), .A2(n1773), .B1(n1772), .B2(n2240), .ZN(n1474)
         );
  OAI22_X1 U2217 ( .A1(n1998), .A2(n1779), .B1(n1778), .B2(n2240), .ZN(n1480)
         );
  OAI22_X1 U2218 ( .A1(n2223), .A2(n1777), .B1(n1776), .B2(n2240), .ZN(n1478)
         );
  OAI22_X1 U2219 ( .A1(n2222), .A2(n1771), .B1(n1770), .B2(n2240), .ZN(n1472)
         );
  OAI22_X1 U2220 ( .A1(n1998), .A2(n1775), .B1(n1774), .B2(n2240), .ZN(n1476)
         );
  OAI22_X1 U2221 ( .A1(n2223), .A2(n1770), .B1(n1769), .B2(n2240), .ZN(n1471)
         );
  OAI22_X1 U2222 ( .A1(n1998), .A2(n1769), .B1(n1768), .B2(n2240), .ZN(n1470)
         );
  OAI22_X1 U2223 ( .A1(n2222), .A2(n1778), .B1(n1777), .B2(n2240), .ZN(n1479)
         );
  OAI22_X1 U2224 ( .A1(n2223), .A2(n1774), .B1(n1773), .B2(n2240), .ZN(n1475)
         );
  XNOR2_X1 U2225 ( .A(b[1]), .B(n2299), .ZN(n1779) );
  XNOR2_X1 U2226 ( .A(b[9]), .B(n2299), .ZN(n1771) );
  XNOR2_X1 U2227 ( .A(b[5]), .B(n2299), .ZN(n1775) );
  XNOR2_X1 U2228 ( .A(b[23]), .B(n2299), .ZN(n1757) );
  XNOR2_X1 U2229 ( .A(b[3]), .B(n2299), .ZN(n1777) );
  XNOR2_X1 U2230 ( .A(b[7]), .B(n2299), .ZN(n1773) );
  XOR2_X1 U2231 ( .A(a[0]), .B(n2300), .Z(n1817) );
  XOR2_X1 U2232 ( .A(n1415), .B(n1393), .Z(n2177) );
  XOR2_X1 U2233 ( .A(n1000), .B(n2177), .Z(n975) );
  NAND2_X1 U2234 ( .A1(n1000), .A2(n1415), .ZN(n2178) );
  NAND2_X1 U2235 ( .A1(n1000), .A2(n1393), .ZN(n2179) );
  NAND2_X1 U2236 ( .A1(n1415), .A2(n1393), .ZN(n2180) );
  NAND3_X1 U2237 ( .A1(n2178), .A2(n2179), .A3(n2180), .ZN(n974) );
  AND2_X1 U2238 ( .A1(n2202), .A2(n2203), .ZN(n2181) );
  OR2_X1 U2239 ( .A1(n2207), .A2(n1553), .ZN(n2182) );
  OR2_X1 U2240 ( .A1(n1552), .A2(n2151), .ZN(n2183) );
  NAND2_X1 U2241 ( .A1(n2182), .A2(n2183), .ZN(n1262) );
  XNOR2_X1 U2242 ( .A(n2252), .B(b[2]), .ZN(n1553) );
  XNOR2_X1 U2243 ( .A(b[3]), .B(n2251), .ZN(n1552) );
  XNOR2_X1 U2244 ( .A(n533), .B(n320), .ZN(product[26]) );
  XNOR2_X1 U2245 ( .A(n522), .B(n319), .ZN(product[27]) );
  XNOR2_X1 U2246 ( .A(n515), .B(n318), .ZN(product[28]) );
  XNOR2_X1 U2247 ( .A(n504), .B(n317), .ZN(product[29]) );
  XNOR2_X1 U2248 ( .A(n497), .B(n316), .ZN(product[30]) );
  XNOR2_X1 U2249 ( .A(n486), .B(n315), .ZN(product[31]) );
  XNOR2_X1 U2250 ( .A(n475), .B(n314), .ZN(product[32]) );
  XNOR2_X1 U2251 ( .A(n462), .B(n313), .ZN(product[33]) );
  INV_X1 U2252 ( .A(n461), .ZN(n459) );
  NAND2_X1 U2253 ( .A1(n749), .A2(n760), .ZN(n439) );
  NOR2_X1 U2254 ( .A1(n749), .A2(n760), .ZN(n438) );
  XOR2_X1 U2255 ( .A(n795), .B(n810), .Z(n2184) );
  XOR2_X1 U2256 ( .A(n808), .B(n2184), .Z(n791) );
  NAND2_X1 U2257 ( .A1(n808), .A2(n795), .ZN(n2185) );
  NAND2_X1 U2258 ( .A1(n808), .A2(n810), .ZN(n2186) );
  NAND2_X1 U2259 ( .A1(n795), .A2(n810), .ZN(n2187) );
  NAND3_X1 U2260 ( .A1(n2185), .A2(n2186), .A3(n2187), .ZN(n790) );
  AND2_X1 U2261 ( .A1(n2202), .A2(n2203), .ZN(n2189) );
  AND2_X1 U2262 ( .A1(n2202), .A2(n2203), .ZN(n2188) );
  AND2_X1 U2263 ( .A1(n2202), .A2(n2203), .ZN(n301) );
  XOR2_X1 U2264 ( .A(n780), .B(n767), .Z(n2190) );
  XOR2_X1 U2265 ( .A(n778), .B(n2190), .Z(n763) );
  NAND2_X1 U2266 ( .A1(n778), .A2(n780), .ZN(n2191) );
  NAND2_X1 U2267 ( .A1(n778), .A2(n767), .ZN(n2192) );
  NAND2_X1 U2268 ( .A1(n780), .A2(n767), .ZN(n2193) );
  NAND3_X1 U2269 ( .A1(n2191), .A2(n2192), .A3(n2193), .ZN(n762) );
  INV_X1 U2270 ( .A(n2249), .ZN(n2245) );
  NAND2_X1 U2271 ( .A1(n672), .A2(n535), .ZN(n321) );
  INV_X1 U2272 ( .A(n2221), .ZN(n2220) );
  NAND2_X1 U2273 ( .A1(n897), .A2(n918), .ZN(n535) );
  INV_X1 U2274 ( .A(n439), .ZN(n445) );
  NAND2_X1 U2275 ( .A1(n1995), .A2(n940), .ZN(n543) );
  INV_X1 U2276 ( .A(n428), .ZN(n661) );
  OAI21_X1 U2277 ( .B1(n428), .B2(n436), .A(n429), .ZN(n427) );
  INV_X1 U2278 ( .A(n2281), .ZN(n2277) );
  OAI21_X1 U2279 ( .B1(n2042), .B2(n535), .A(n532), .ZN(n526) );
  NAND2_X1 U2280 ( .A1(n666), .A2(n2102), .ZN(n467) );
  INV_X1 U2281 ( .A(n2162), .ZN(n565) );
  INV_X1 U2282 ( .A(n490), .ZN(n492) );
  OAI21_X1 U2283 ( .B1(n495), .B2(n503), .A(n496), .ZN(n490) );
  CLKBUF_X1 U2284 ( .A(n2201), .Z(n2195) );
  NOR2_X1 U2285 ( .A1(n857), .A2(n876), .ZN(n520) );
  NOR2_X1 U2286 ( .A1(n491), .A2(n480), .ZN(n478) );
  OAI21_X1 U2287 ( .B1(n492), .B2(n480), .A(n481), .ZN(n479) );
  INV_X1 U2288 ( .A(n480), .ZN(n666) );
  NOR2_X1 U2289 ( .A1(n571), .A2(n569), .ZN(n567) );
  NAND2_X1 U2290 ( .A1(n1003), .A2(n1020), .ZN(n570) );
  NOR2_X1 U2291 ( .A1(n1003), .A2(n1020), .ZN(n569) );
  NAND2_X1 U2292 ( .A1(n709), .A2(n716), .ZN(n409) );
  NOR2_X1 U2293 ( .A1(n1935), .A2(n2051), .ZN(n545) );
  OAI21_X1 U2294 ( .B1(n555), .B2(n2051), .A(n550), .ZN(n546) );
  NAND2_X1 U2295 ( .A1(n941), .A2(n962), .ZN(n550) );
  NAND2_X1 U2296 ( .A1(n588), .A2(n2104), .ZN(n582) );
  AOI21_X1 U2297 ( .B1(n589), .B2(n2104), .A(n2107), .ZN(n583) );
  AOI21_X1 U2298 ( .B1(n565), .B2(n2043), .A(n2041), .ZN(n551) );
  INV_X1 U2299 ( .A(n2041), .ZN(n555) );
  NOR2_X1 U2300 ( .A1(n558), .A2(n563), .ZN(n552) );
  OAI21_X1 U2301 ( .B1(n1965), .B2(n564), .A(n559), .ZN(n553) );
  NAND2_X1 U2302 ( .A1(n996), .A2(n994), .ZN(n2196) );
  NAND2_X1 U2303 ( .A1(n996), .A2(n1217), .ZN(n2197) );
  NAND2_X1 U2304 ( .A1(n994), .A2(n1217), .ZN(n2198) );
  NAND3_X1 U2305 ( .A1(n2196), .A2(n2197), .A3(n2198), .ZN(n972) );
  OR2_X1 U2306 ( .A1(n2217), .A2(n1668), .ZN(n2199) );
  OR2_X1 U2307 ( .A1(n1667), .A2(n2150), .ZN(n2200) );
  NAND2_X1 U2308 ( .A1(n2199), .A2(n2200), .ZN(n1372) );
  AOI21_X1 U2309 ( .B1(n1997), .B2(n1936), .A(n2166), .ZN(n2201) );
  XNOR2_X1 U2310 ( .A(n2279), .B(b[12]), .ZN(n1668) );
  NOR2_X1 U2311 ( .A1(n590), .A2(n592), .ZN(n588) );
  INV_X1 U2312 ( .A(n383), .ZN(n381) );
  AOI21_X1 U2313 ( .B1(n383), .B2(n2164), .A(n376), .ZN(n372) );
  NAND2_X1 U2314 ( .A1(n552), .A2(n540), .ZN(n538) );
  OAI22_X1 U2315 ( .A1(n2077), .A2(n1508), .B1(n1507), .B2(n2225), .ZN(n682)
         );
  OAI22_X1 U2316 ( .A1(n2077), .A2(n1518), .B1(n1517), .B2(n2225), .ZN(n1228)
         );
  OAI22_X1 U2317 ( .A1(n2077), .A2(n1510), .B1(n1509), .B2(n2225), .ZN(n1220)
         );
  OAI22_X1 U2318 ( .A1(n2077), .A2(n1514), .B1(n1513), .B2(n2225), .ZN(n1224)
         );
  OAI22_X1 U2319 ( .A1(n2077), .A2(n1512), .B1(n1511), .B2(n2226), .ZN(n1222)
         );
  OAI22_X1 U2320 ( .A1(n2077), .A2(n2249), .B1(n1531), .B2(n2226), .ZN(n1183)
         );
  OAI22_X1 U2321 ( .A1(n2077), .A2(n1516), .B1(n1515), .B2(n2226), .ZN(n1226)
         );
  OAI21_X1 U2322 ( .B1(n337), .B2(n334), .A(n335), .ZN(n333) );
  NAND2_X1 U2323 ( .A1(n685), .A2(n688), .ZN(n369) );
  AOI21_X1 U2324 ( .B1(n595), .B2(n609), .A(n596), .ZN(n594) );
  NAND2_X1 U2325 ( .A1(n1171), .A2(n1174), .ZN(n634) );
  NOR2_X1 U2326 ( .A1(n1171), .A2(n1174), .ZN(n633) );
  OAI21_X1 U2327 ( .B1(n390), .B2(n384), .A(n387), .ZN(n383) );
  OAI21_X1 U2328 ( .B1(n456), .B2(n481), .A(n457), .ZN(n455) );
  NOR2_X1 U2329 ( .A1(n456), .A2(n480), .ZN(n454) );
  OAI22_X1 U2330 ( .A1(n2216), .A2(n1671), .B1(n2234), .B2(n1670), .ZN(n1375)
         );
  OAI22_X1 U2331 ( .A1(n2216), .A2(n1672), .B1(n1671), .B2(n2234), .ZN(n1376)
         );
  OAI22_X1 U2332 ( .A1(n2216), .A2(n1676), .B1(n1675), .B2(n2234), .ZN(n1380)
         );
  OAI22_X1 U2333 ( .A1(n2216), .A2(n1679), .B1(n2234), .B2(n1678), .ZN(n1383)
         );
  OAI22_X1 U2334 ( .A1(n2216), .A2(n1669), .B1(n2234), .B2(n1668), .ZN(n1373)
         );
  OAI22_X1 U2335 ( .A1(n2216), .A2(n1670), .B1(n1669), .B2(n2234), .ZN(n1374)
         );
  AOI21_X1 U2336 ( .B1(n2103), .B2(n2106), .A(n1941), .ZN(n572) );
  NAND2_X1 U2337 ( .A1(n1929), .A2(n2105), .ZN(n571) );
  INV_X1 U2338 ( .A(n2083), .ZN(n524) );
  AOI21_X1 U2339 ( .B1(n2083), .B2(n2160), .A(n2088), .ZN(n517) );
  AOI21_X1 U2340 ( .B1(n2102), .B2(n483), .A(n472), .ZN(n468) );
  AOI21_X1 U2341 ( .B1(n2114), .B2(n472), .A(n459), .ZN(n457) );
  INV_X1 U2342 ( .A(n2201), .ZN(n508) );
  NAND2_X1 U2343 ( .A1(n2159), .A2(n2160), .ZN(n516) );
  INV_X1 U2344 ( .A(n534), .ZN(n672) );
  NAND2_X1 U2345 ( .A1(n525), .A2(n511), .ZN(n505) );
  OAI21_X1 U2346 ( .B1(n620), .B2(n610), .A(n611), .ZN(n609) );
  NOR2_X1 U2347 ( .A1(n513), .A2(n520), .ZN(n511) );
  INV_X1 U2348 ( .A(n1982), .ZN(n491) );
  NAND2_X1 U2349 ( .A1(n454), .A2(n489), .ZN(n452) );
  NOR2_X1 U2350 ( .A1(n336), .A2(n334), .ZN(n332) );
  NAND2_X1 U2351 ( .A1(n717), .A2(n726), .ZN(n418) );
  NAND2_X1 U2352 ( .A1(n983), .A2(n1002), .ZN(n564) );
  OAI21_X1 U2353 ( .B1(n1933), .B2(n550), .A(n543), .ZN(n541) );
  XNOR2_X1 U2354 ( .A(b[21]), .B(n2256), .ZN(n1559) );
  XNOR2_X1 U2355 ( .A(b[17]), .B(n2256), .ZN(n1563) );
  XNOR2_X1 U2356 ( .A(b[15]), .B(n2256), .ZN(n1565) );
  XNOR2_X1 U2357 ( .A(b[19]), .B(n2256), .ZN(n1561) );
  XNOR2_X1 U2358 ( .A(b[11]), .B(n2256), .ZN(n1569) );
  XNOR2_X1 U2359 ( .A(b[13]), .B(n2256), .ZN(n1567) );
  INV_X1 U2360 ( .A(n382), .ZN(n380) );
  NAND2_X1 U2361 ( .A1(n382), .A2(n2164), .ZN(n371) );
  NOR2_X1 U2362 ( .A1(n389), .A2(n384), .ZN(n382) );
  XNOR2_X1 U2363 ( .A(b[17]), .B(n2245), .ZN(n1513) );
  XNOR2_X1 U2364 ( .A(b[21]), .B(n2245), .ZN(n1509) );
  XNOR2_X1 U2365 ( .A(b[19]), .B(n2245), .ZN(n1511) );
  XNOR2_X1 U2366 ( .A(b[11]), .B(n2245), .ZN(n1519) );
  XNOR2_X1 U2367 ( .A(b[13]), .B(n2245), .ZN(n1517) );
  XNOR2_X1 U2368 ( .A(b[15]), .B(n2245), .ZN(n1515) );
  NAND2_X1 U2369 ( .A1(n963), .A2(n982), .ZN(n559) );
  NOR2_X1 U2370 ( .A1(n918), .A2(n897), .ZN(n534) );
  NOR2_X1 U2371 ( .A1(n2063), .A2(n547), .ZN(n540) );
  OAI21_X1 U2372 ( .B1(n572), .B2(n1951), .A(n570), .ZN(n568) );
  OAI21_X1 U2373 ( .B1(n594), .B2(n582), .A(n583), .ZN(n581) );
  NAND2_X1 U2374 ( .A1(n2113), .A2(n2097), .ZN(n599) );
  NAND2_X1 U2375 ( .A1(n1071), .A2(n1084), .ZN(n591) );
  OAI22_X1 U2376 ( .A1(n2011), .A2(n1750), .B1(n2239), .B2(n1749), .ZN(n1451)
         );
  OAI22_X1 U2377 ( .A1(n2012), .A2(n1749), .B1(n1748), .B2(n2239), .ZN(n1450)
         );
  OAI22_X1 U2378 ( .A1(n2012), .A2(n1753), .B1(n1752), .B2(n2239), .ZN(n1454)
         );
  OAI22_X1 U2379 ( .A1(n2012), .A2(n1747), .B1(n1746), .B2(n2239), .ZN(n1448)
         );
  OAI22_X1 U2380 ( .A1(n2011), .A2(n1754), .B1(n2239), .B2(n1753), .ZN(n1455)
         );
  OAI22_X1 U2381 ( .A1(n2011), .A2(n1745), .B1(n1744), .B2(n2239), .ZN(n1446)
         );
  OAI22_X1 U2382 ( .A1(n2216), .A2(n1678), .B1(n1677), .B2(n2150), .ZN(n1382)
         );
  OAI22_X1 U2383 ( .A1(n2216), .A2(n1674), .B1(n1673), .B2(n2234), .ZN(n1378)
         );
  OAI22_X1 U2384 ( .A1(n2216), .A2(n1680), .B1(n1679), .B2(n2150), .ZN(n1384)
         );
  OAI22_X1 U2385 ( .A1(n2217), .A2(n1673), .B1(n2234), .B2(n1672), .ZN(n1377)
         );
  OAI22_X1 U2386 ( .A1(n2216), .A2(n1675), .B1(n2234), .B2(n1674), .ZN(n1379)
         );
  OAI22_X1 U2387 ( .A1(n2216), .A2(n1677), .B1(n2234), .B2(n1676), .ZN(n1381)
         );
  INV_X1 U2388 ( .A(n401), .ZN(n399) );
  AOI21_X1 U2389 ( .B1(n401), .B2(n2111), .A(n394), .ZN(n390) );
  OAI21_X1 U2390 ( .B1(n2139), .B2(n1994), .A(n2311), .ZN(n1338) );
  INV_X1 U2391 ( .A(n2194), .ZN(n2232) );
  OAI22_X1 U2392 ( .A1(n2012), .A2(n1751), .B1(n1750), .B2(n2239), .ZN(n1452)
         );
  OAI22_X1 U2393 ( .A1(n2012), .A2(n1755), .B1(n1754), .B2(n2239), .ZN(n1456)
         );
  OAI22_X1 U2394 ( .A1(n2011), .A2(n1752), .B1(n2239), .B2(n1751), .ZN(n1453)
         );
  OAI22_X1 U2395 ( .A1(n2012), .A2(n1746), .B1(n2239), .B2(n1745), .ZN(n1447)
         );
  OAI22_X1 U2396 ( .A1(n2012), .A2(n1744), .B1(n2239), .B2(n1743), .ZN(n1445)
         );
  OAI22_X1 U2397 ( .A1(n2012), .A2(n1748), .B1(n2239), .B2(n1747), .ZN(n1449)
         );
  AOI21_X1 U2398 ( .B1(n490), .B2(n2010), .A(n455), .ZN(n453) );
  INV_X1 U2399 ( .A(n874), .ZN(n875) );
  INV_X1 U2400 ( .A(n474), .ZN(n472) );
  NAND2_X1 U2401 ( .A1(n2102), .A2(n474), .ZN(n314) );
  AOI21_X1 U2402 ( .B1(n526), .B2(n2168), .A(n512), .ZN(n506) );
  OAI21_X1 U2403 ( .B1(n2056), .B2(n521), .A(n514), .ZN(n512) );
  OAI21_X1 U2404 ( .B1(n421), .B2(n402), .A(n405), .ZN(n401) );
  INV_X1 U2405 ( .A(n345), .ZN(n343) );
  NAND2_X1 U2406 ( .A1(n345), .A2(n2121), .ZN(n336) );
  XNOR2_X1 U2407 ( .A(b[19]), .B(n2272), .ZN(n1636) );
  XNOR2_X1 U2408 ( .A(b[21]), .B(n2272), .ZN(n1634) );
  XNOR2_X1 U2409 ( .A(b[11]), .B(n2272), .ZN(n1644) );
  XNOR2_X1 U2410 ( .A(b[17]), .B(n2272), .ZN(n1638) );
  XNOR2_X1 U2411 ( .A(b[13]), .B(n2272), .ZN(n1642) );
  XNOR2_X1 U2412 ( .A(b[15]), .B(n2272), .ZN(n1640) );
  OAI22_X1 U2413 ( .A1(n2011), .A2(n2297), .B1(n1756), .B2(n2239), .ZN(n1192)
         );
  OAI22_X1 U2414 ( .A1(n2011), .A2(n1738), .B1(n2239), .B2(n1737), .ZN(n1439)
         );
  OAI22_X1 U2415 ( .A1(n2012), .A2(n1741), .B1(n1740), .B2(n2238), .ZN(n1442)
         );
  OAI22_X1 U2416 ( .A1(n2155), .A2(n1734), .B1(n2238), .B2(n1733), .ZN(n1435)
         );
  OAI22_X1 U2417 ( .A1(n2012), .A2(n1739), .B1(n1738), .B2(n2238), .ZN(n1440)
         );
  OAI22_X1 U2418 ( .A1(n2011), .A2(n1740), .B1(n2238), .B2(n1739), .ZN(n1441)
         );
  OAI22_X1 U2419 ( .A1(n2220), .A2(n1736), .B1(n2238), .B2(n1735), .ZN(n1437)
         );
  OAI22_X1 U2420 ( .A1(n2155), .A2(n1735), .B1(n1734), .B2(n2238), .ZN(n1436)
         );
  OAI22_X1 U2421 ( .A1(n2220), .A2(n1742), .B1(n2238), .B2(n1741), .ZN(n1443)
         );
  OAI22_X1 U2422 ( .A1(n2155), .A2(n1737), .B1(n1736), .B2(n2238), .ZN(n1438)
         );
  OAI22_X1 U2423 ( .A1(n2012), .A2(n1743), .B1(n1742), .B2(n2238), .ZN(n1444)
         );
  OAI22_X1 U2424 ( .A1(n2096), .A2(n1705), .B1(n1704), .B2(n2235), .ZN(n1408)
         );
  OAI22_X1 U2425 ( .A1(n2218), .A2(n1703), .B1(n1702), .B2(n2236), .ZN(n1406)
         );
  AOI21_X1 U2426 ( .B1(n553), .B2(n540), .A(n541), .ZN(n539) );
  NAND2_X1 U2427 ( .A1(n400), .A2(n2111), .ZN(n389) );
  NAND2_X1 U2428 ( .A1(n2174), .A2(n2093), .ZN(n487) );
  NAND2_X1 U2429 ( .A1(n2174), .A2(n668), .ZN(n498) );
  NAND2_X1 U2430 ( .A1(n478), .A2(n2174), .ZN(n476) );
  NAND2_X1 U2431 ( .A1(n465), .A2(n2174), .ZN(n463) );
  NAND2_X1 U2432 ( .A1(n839), .A2(n856), .ZN(n514) );
  OAI22_X1 U2433 ( .A1(n2149), .A2(n2293), .B1(n1731), .B2(n2061), .ZN(n1191)
         );
  OAI22_X1 U2434 ( .A1(n2149), .A2(n1718), .B1(n1717), .B2(n2061), .ZN(n1420)
         );
  OAI22_X1 U2435 ( .A1(n1957), .A2(n1711), .B1(n1969), .B2(n1710), .ZN(n1413)
         );
  OAI22_X1 U2436 ( .A1(n2148), .A2(n1716), .B1(n1715), .B2(n1969), .ZN(n1418)
         );
  OAI22_X1 U2437 ( .A1(n1957), .A2(n1713), .B1(n2237), .B2(n1712), .ZN(n1415)
         );
  OAI22_X1 U2438 ( .A1(n1957), .A2(n1717), .B1(n2061), .B2(n1716), .ZN(n1419)
         );
  OAI22_X1 U2439 ( .A1(n2148), .A2(n1715), .B1(n2061), .B2(n1714), .ZN(n1417)
         );
  OAI22_X1 U2440 ( .A1(n1957), .A2(n1708), .B1(n1707), .B2(n2237), .ZN(n874)
         );
  OAI22_X1 U2441 ( .A1(n2148), .A2(n1709), .B1(n2237), .B2(n1708), .ZN(n1411)
         );
  OAI22_X1 U2442 ( .A1(n1957), .A2(n1710), .B1(n1709), .B2(n2237), .ZN(n1412)
         );
  OAI22_X1 U2443 ( .A1(n1957), .A2(n1714), .B1(n1713), .B2(n2237), .ZN(n1416)
         );
  OAI22_X1 U2444 ( .A1(n1957), .A2(n1712), .B1(n1711), .B2(n1969), .ZN(n1414)
         );
  NAND2_X1 U2445 ( .A1(n2102), .A2(n2114), .ZN(n456) );
  OAI21_X1 U2446 ( .B1(n638), .B2(n636), .A(n637), .ZN(n635) );
  NOR2_X1 U2447 ( .A1(n633), .A2(n631), .ZN(n629) );
  AOI21_X1 U2448 ( .B1(n508), .B2(n668), .A(n501), .ZN(n499) );
  AOI21_X1 U2449 ( .B1(n508), .B2(n465), .A(n466), .ZN(n464) );
  AOI21_X1 U2450 ( .B1(n508), .B2(n478), .A(n479), .ZN(n477) );
  AOI21_X1 U2451 ( .B1(n508), .B2(n2093), .A(n1979), .ZN(n488) );
  OAI22_X1 U2452 ( .A1(n2206), .A2(n1483), .B1(n1482), .B2(n2147), .ZN(n676)
         );
  OAI22_X1 U2453 ( .A1(n2206), .A2(n1485), .B1(n1484), .B2(n2147), .ZN(n1196)
         );
  OAI22_X1 U2454 ( .A1(n2206), .A2(n1491), .B1(n1490), .B2(n2147), .ZN(n1202)
         );
  OAI22_X1 U2455 ( .A1(n2206), .A2(n1487), .B1(n1486), .B2(n2147), .ZN(n1198)
         );
  OAI22_X1 U2456 ( .A1(n2206), .A2(n1489), .B1(n1488), .B2(n2147), .ZN(n1200)
         );
  XNOR2_X1 U2457 ( .A(n2034), .B(n2057), .ZN(n939) );
  OR2_X1 U2458 ( .A1(n1215), .A2(n1237), .ZN(n938) );
  OAI22_X1 U2459 ( .A1(n2206), .A2(n1493), .B1(n1492), .B2(n2147), .ZN(n1204)
         );
  OAI22_X1 U2460 ( .A1(n2206), .A2(n1949), .B1(n1506), .B2(n2147), .ZN(n1182)
         );
  OAI22_X1 U2461 ( .A1(n2212), .A2(n1613), .B1(n2231), .B2(n1612), .ZN(n1319)
         );
  INV_X1 U2462 ( .A(n746), .ZN(n747) );
  OAI22_X1 U2463 ( .A1(n2212), .A2(n1612), .B1(n1611), .B2(n2146), .ZN(n1318)
         );
  OAI22_X1 U2464 ( .A1(n2212), .A2(n2270), .B1(n1631), .B2(n2146), .ZN(n1187)
         );
  OAI22_X1 U2465 ( .A1(n2213), .A2(n1611), .B1(n2231), .B2(n1610), .ZN(n1317)
         );
  OAI22_X1 U2466 ( .A1(n2212), .A2(n1617), .B1(n2231), .B2(n1616), .ZN(n1323)
         );
  OAI22_X1 U2467 ( .A1(n2212), .A2(n1615), .B1(n2231), .B2(n1614), .ZN(n1321)
         );
  OAI22_X1 U2468 ( .A1(n2212), .A2(n1610), .B1(n1609), .B2(n2146), .ZN(n1316)
         );
  OAI22_X1 U2469 ( .A1(n2213), .A2(n1614), .B1(n1613), .B2(n2146), .ZN(n1320)
         );
  OAI22_X1 U2470 ( .A1(n2212), .A2(n1609), .B1(n2231), .B2(n1608), .ZN(n1315)
         );
  OAI22_X1 U2471 ( .A1(n2213), .A2(n1616), .B1(n1615), .B2(n2146), .ZN(n1322)
         );
  OAI22_X1 U2472 ( .A1(n2212), .A2(n1618), .B1(n1617), .B2(n2146), .ZN(n1324)
         );
  OAI22_X1 U2473 ( .A1(n2212), .A2(n1608), .B1(n1607), .B2(n2146), .ZN(n746)
         );
  NAND2_X1 U2474 ( .A1(n537), .A2(n450), .ZN(n2202) );
  INV_X1 U2475 ( .A(n451), .ZN(n2203) );
  OAI22_X1 U2476 ( .A1(n2011), .A2(n1733), .B1(n1732), .B2(n2238), .ZN(n2204)
         );
  OAI21_X1 U2477 ( .B1(n566), .B2(n538), .A(n539), .ZN(n537) );
  OAI22_X1 U2478 ( .A1(n2212), .A2(n1620), .B1(n1619), .B2(n1934), .ZN(n1326)
         );
  OAI22_X1 U2479 ( .A1(n2212), .A2(n1626), .B1(n1625), .B2(n1934), .ZN(n1332)
         );
  OAI22_X1 U2480 ( .A1(n2212), .A2(n1623), .B1(n2231), .B2(n1622), .ZN(n1329)
         );
  OAI22_X1 U2481 ( .A1(n2212), .A2(n1630), .B1(n1629), .B2(n2146), .ZN(n1336)
         );
  OAI22_X1 U2482 ( .A1(n2212), .A2(n1619), .B1(n2231), .B2(n1618), .ZN(n1325)
         );
  OAI22_X1 U2483 ( .A1(n2212), .A2(n1625), .B1(n2231), .B2(n1624), .ZN(n1331)
         );
  OAI22_X1 U2484 ( .A1(n2212), .A2(n1629), .B1(n1934), .B2(n1628), .ZN(n1335)
         );
  OAI22_X1 U2485 ( .A1(n2212), .A2(n1621), .B1(n1934), .B2(n1620), .ZN(n1327)
         );
  OAI22_X1 U2486 ( .A1(n2213), .A2(n1627), .B1(n2231), .B2(n1626), .ZN(n1333)
         );
  OAI22_X1 U2487 ( .A1(n2213), .A2(n1622), .B1(n1621), .B2(n2231), .ZN(n1328)
         );
  OAI22_X1 U2488 ( .A1(n2213), .A2(n1624), .B1(n1623), .B2(n2231), .ZN(n1330)
         );
  OAI22_X1 U2489 ( .A1(n2213), .A2(n1628), .B1(n1627), .B2(n2146), .ZN(n1334)
         );
  OAI21_X1 U2490 ( .B1(n506), .B2(n452), .A(n453), .ZN(n451) );
  NOR2_X1 U2491 ( .A1(n505), .A2(n452), .ZN(n450) );
  INV_X1 U2492 ( .A(n537), .ZN(n536) );
  OAI22_X1 U2493 ( .A1(n1930), .A2(n1652), .B1(n2232), .B2(n1651), .ZN(n1357)
         );
  OAI22_X1 U2494 ( .A1(n1930), .A2(n1649), .B1(n1648), .B2(n2232), .ZN(n1354)
         );
  OAI22_X1 U2495 ( .A1(n2072), .A2(n1653), .B1(n1652), .B2(n2154), .ZN(n1358)
         );
  OAI22_X1 U2496 ( .A1(n2072), .A2(n1648), .B1(n2232), .B2(n1647), .ZN(n1353)
         );
  OAI22_X1 U2497 ( .A1(n2073), .A2(n1647), .B1(n1646), .B2(n2232), .ZN(n1352)
         );
  OAI22_X1 U2498 ( .A1(n2215), .A2(n1645), .B1(n1644), .B2(n2232), .ZN(n1350)
         );
  OAI22_X1 U2499 ( .A1(n1931), .A2(n1654), .B1(n2232), .B2(n1653), .ZN(n1359)
         );
  OAI22_X1 U2500 ( .A1(n2072), .A2(n1650), .B1(n2232), .B2(n1649), .ZN(n1355)
         );
  OAI22_X1 U2501 ( .A1(n1931), .A2(n1644), .B1(n2233), .B2(n1643), .ZN(n1349)
         );
  OAI22_X1 U2502 ( .A1(n2073), .A2(n1655), .B1(n1654), .B2(n2154), .ZN(n1360)
         );
  OAI22_X1 U2503 ( .A1(n2214), .A2(n1646), .B1(n2233), .B2(n1645), .ZN(n1351)
         );
  OAI22_X1 U2504 ( .A1(n2072), .A2(n1651), .B1(n1650), .B2(n2232), .ZN(n1356)
         );
  XNOR2_X1 U2505 ( .A(b[17]), .B(n2277), .ZN(n1663) );
  XNOR2_X1 U2506 ( .A(b[11]), .B(n2277), .ZN(n1669) );
  XNOR2_X1 U2507 ( .A(b[19]), .B(n2277), .ZN(n1661) );
  XNOR2_X1 U2508 ( .A(b[13]), .B(n2277), .ZN(n1667) );
  XNOR2_X1 U2509 ( .A(b[15]), .B(n2277), .ZN(n1665) );
  XNOR2_X1 U2510 ( .A(b[21]), .B(n2277), .ZN(n1659) );
  OAI22_X1 U2511 ( .A1(n1977), .A2(n1571), .B1(n2153), .B2(n1570), .ZN(n1279)
         );
  OAI22_X1 U2512 ( .A1(n1976), .A2(n1570), .B1(n1569), .B2(n2228), .ZN(n1278)
         );
  OAI22_X1 U2513 ( .A1(n1977), .A2(n1575), .B1(n2228), .B2(n1574), .ZN(n1283)
         );
  OAI22_X1 U2514 ( .A1(n1977), .A2(n1580), .B1(n1579), .B2(n2153), .ZN(n1288)
         );
  OAI22_X1 U2515 ( .A1(n1977), .A2(n1579), .B1(n2228), .B2(n1578), .ZN(n1287)
         );
  OAI22_X1 U2516 ( .A1(n1976), .A2(n1573), .B1(n2228), .B2(n1572), .ZN(n1281)
         );
  OAI22_X1 U2517 ( .A1(n1976), .A2(n1569), .B1(n2228), .B2(n1568), .ZN(n1277)
         );
  OAI22_X1 U2518 ( .A1(n1976), .A2(n1578), .B1(n1577), .B2(n2153), .ZN(n1286)
         );
  OAI22_X1 U2519 ( .A1(n2210), .A2(n1577), .B1(n2228), .B2(n1576), .ZN(n1285)
         );
  OAI22_X1 U2520 ( .A1(n1977), .A2(n1572), .B1(n1571), .B2(n2228), .ZN(n1280)
         );
  XNOR2_X1 U2521 ( .A(b[21]), .B(n2264), .ZN(n1584) );
  XNOR2_X1 U2522 ( .A(b[17]), .B(n1961), .ZN(n1588) );
  OAI22_X1 U2523 ( .A1(n2210), .A2(n1574), .B1(n1573), .B2(n2228), .ZN(n1282)
         );
  OAI22_X1 U2524 ( .A1(n2209), .A2(n1576), .B1(n1575), .B2(n2228), .ZN(n1284)
         );
  XNOR2_X1 U2525 ( .A(b[15]), .B(n1960), .ZN(n1590) );
  XNOR2_X1 U2526 ( .A(b[13]), .B(n2264), .ZN(n1592) );
  XNOR2_X1 U2527 ( .A(b[19]), .B(n1961), .ZN(n1586) );
  XNOR2_X1 U2528 ( .A(b[11]), .B(n1961), .ZN(n1594) );
  OAI22_X1 U2529 ( .A1(n2156), .A2(n1535), .B1(n1534), .B2(n2151), .ZN(n1244)
         );
  OAI22_X1 U2530 ( .A1(n1537), .A2(n1990), .B1(n1536), .B2(n2151), .ZN(n1246)
         );
  OAI22_X1 U2531 ( .A1(n2157), .A2(n1533), .B1(n1532), .B2(n2151), .ZN(n692)
         );
  OAI22_X1 U2532 ( .A1(n2157), .A2(n1543), .B1(n1542), .B2(n2151), .ZN(n1252)
         );
  OAI22_X1 U2533 ( .A1(n2208), .A2(n1539), .B1(n1538), .B2(n2151), .ZN(n1248)
         );
  OAI22_X1 U2534 ( .A1(n1990), .A2(n2254), .B1(n1556), .B2(n2151), .ZN(n1184)
         );
  OAI22_X1 U2535 ( .A1(n2157), .A2(n1541), .B1(n1540), .B2(n2151), .ZN(n1250)
         );
  INV_X1 U2536 ( .A(n421), .ZN(n423) );
  OAI21_X1 U2537 ( .B1(n421), .B2(n347), .A(n348), .ZN(n346) );
  OAI22_X1 U2538 ( .A1(n2211), .A2(n1593), .B1(n1592), .B2(n2230), .ZN(n1300)
         );
  OAI22_X1 U2539 ( .A1(n2211), .A2(n1590), .B1(n2230), .B2(n1589), .ZN(n1297)
         );
  OAI22_X1 U2540 ( .A1(n2211), .A2(n1584), .B1(n2230), .B2(n1583), .ZN(n1291)
         );
  OAI22_X1 U2541 ( .A1(n2211), .A2(n1589), .B1(n1588), .B2(n2229), .ZN(n1296)
         );
  OAI22_X1 U2542 ( .A1(n2211), .A2(n1583), .B1(n1582), .B2(n2230), .ZN(n724)
         );
  OAI22_X1 U2543 ( .A1(n2015), .A2(n1588), .B1(n2230), .B2(n1587), .ZN(n1295)
         );
  OAI22_X1 U2544 ( .A1(n2211), .A2(n1585), .B1(n1584), .B2(n2229), .ZN(n1292)
         );
  OAI22_X1 U2545 ( .A1(n2015), .A2(n1592), .B1(n2230), .B2(n1591), .ZN(n1299)
         );
  OAI22_X1 U2546 ( .A1(n2015), .A2(n1587), .B1(n1586), .B2(n2230), .ZN(n1294)
         );
  OAI22_X1 U2547 ( .A1(n2211), .A2(n1591), .B1(n1590), .B2(n2229), .ZN(n1298)
         );
  OAI22_X1 U2548 ( .A1(n2211), .A2(n1586), .B1(n2230), .B2(n1585), .ZN(n1293)
         );
  OAI22_X1 U2549 ( .A1(n2211), .A2(n2265), .B1(n1606), .B2(n2229), .ZN(n1186)
         );
  XNOR2_X1 U2550 ( .A(b[19]), .B(n2267), .ZN(n1611) );
  XNOR2_X1 U2551 ( .A(b[11]), .B(n2267), .ZN(n1619) );
  XNOR2_X1 U2552 ( .A(b[17]), .B(n1988), .ZN(n1613) );
  XNOR2_X1 U2553 ( .A(b[13]), .B(n1989), .ZN(n1617) );
  XNOR2_X1 U2554 ( .A(b[21]), .B(n1989), .ZN(n1609) );
  XNOR2_X1 U2555 ( .A(b[15]), .B(n1988), .ZN(n1615) );
  NAND2_X1 U2556 ( .A1(n332), .A2(n2128), .ZN(n326) );
  AOI21_X1 U2557 ( .B1(n333), .B2(n2128), .A(n2129), .ZN(n327) );
  NAND2_X1 U2558 ( .A1(n356), .A2(n2120), .ZN(n347) );
  XNOR2_X1 U2559 ( .A(n437), .B(n311), .ZN(product[35]) );
  XNOR2_X1 U2560 ( .A(b[11]), .B(n2289), .ZN(n1719) );
  XNOR2_X1 U2561 ( .A(b[13]), .B(n2289), .ZN(n1717) );
  XNOR2_X1 U2562 ( .A(b[15]), .B(n2289), .ZN(n1715) );
  XNOR2_X1 U2563 ( .A(b[21]), .B(n2289), .ZN(n1709) );
  XNOR2_X1 U2564 ( .A(b[19]), .B(n2289), .ZN(n1711) );
  XNOR2_X1 U2565 ( .A(b[17]), .B(n2289), .ZN(n1713) );
  OAI22_X1 U2566 ( .A1(n2216), .A2(n1661), .B1(n2234), .B2(n1660), .ZN(n1365)
         );
  OAI22_X1 U2567 ( .A1(n2216), .A2(n1660), .B1(n1659), .B2(n2150), .ZN(n1364)
         );
  OAI22_X1 U2568 ( .A1(n2216), .A2(n1663), .B1(n2234), .B2(n1662), .ZN(n1367)
         );
  OAI22_X1 U2569 ( .A1(n2216), .A2(n1987), .B1(n1681), .B2(n2150), .ZN(n1189)
         );
  OAI22_X1 U2570 ( .A1(n2216), .A2(n1664), .B1(n1663), .B2(n2150), .ZN(n1368)
         );
  OAI22_X1 U2571 ( .A1(n2217), .A2(n1658), .B1(n1657), .B2(n2150), .ZN(n802)
         );
  OAI22_X1 U2572 ( .A1(n2216), .A2(n1667), .B1(n2234), .B2(n1666), .ZN(n1371)
         );
  OAI22_X1 U2573 ( .A1(n2217), .A2(n1665), .B1(n2234), .B2(n1664), .ZN(n1369)
         );
  OAI22_X1 U2574 ( .A1(n2217), .A2(n1662), .B1(n1661), .B2(n2150), .ZN(n1366)
         );
  OAI22_X1 U2575 ( .A1(n2217), .A2(n1666), .B1(n1665), .B2(n2150), .ZN(n1370)
         );
  OAI22_X1 U2576 ( .A1(n2217), .A2(n1659), .B1(n2234), .B2(n1658), .ZN(n1363)
         );
  XNOR2_X1 U2577 ( .A(b[17]), .B(n2283), .ZN(n1688) );
  XNOR2_X1 U2578 ( .A(b[19]), .B(n2283), .ZN(n1686) );
  XNOR2_X1 U2579 ( .A(b[15]), .B(n2283), .ZN(n1690) );
  XNOR2_X1 U2580 ( .A(b[21]), .B(n2283), .ZN(n1684) );
  XNOR2_X1 U2581 ( .A(b[11]), .B(n2283), .ZN(n1694) );
  XNOR2_X1 U2582 ( .A(b[13]), .B(n2283), .ZN(n1692) );
  XNOR2_X1 U2583 ( .A(n430), .B(n310), .ZN(product[36]) );
  OAI22_X1 U2584 ( .A1(n2156), .A2(n1544), .B1(n2227), .B2(n1543), .ZN(n1253)
         );
  OAI22_X1 U2585 ( .A1(n1546), .A2(n1990), .B1(n2227), .B2(n1545), .ZN(n1255)
         );
  OAI22_X1 U2586 ( .A1(n2208), .A2(n1552), .B1(n2227), .B2(n1551), .ZN(n1261)
         );
  OAI22_X1 U2587 ( .A1(n2207), .A2(n1548), .B1(n2227), .B2(n1547), .ZN(n1257)
         );
  OAI22_X1 U2588 ( .A1(n2157), .A2(n1549), .B1(n1548), .B2(n2151), .ZN(n1258)
         );
  OAI22_X1 U2589 ( .A1(n2157), .A2(n1555), .B1(n1554), .B2(n2151), .ZN(n1264)
         );
  OAI22_X1 U2590 ( .A1(n2207), .A2(n1547), .B1(n1546), .B2(n2151), .ZN(n1256)
         );
  OAI22_X1 U2591 ( .A1(n2156), .A2(n1545), .B1(n1544), .B2(n2227), .ZN(n1254)
         );
  OAI22_X1 U2592 ( .A1(n1990), .A2(n1550), .B1(n2227), .B2(n1549), .ZN(n1259)
         );
  OAI22_X1 U2593 ( .A1(n1554), .A2(n1990), .B1(n2227), .B2(n1553), .ZN(n1263)
         );
  OAI22_X1 U2594 ( .A1(n2208), .A2(n1551), .B1(n1550), .B2(n2227), .ZN(n1260)
         );
  XNOR2_X1 U2595 ( .A(n419), .B(n309), .ZN(product[37]) );
  OAI22_X1 U2596 ( .A1(n2205), .A2(n1497), .B1(n1496), .B2(n2224), .ZN(n1208)
         );
  OAI22_X1 U2597 ( .A1(n1970), .A2(n1496), .B1(n2147), .B2(n1495), .ZN(n1207)
         );
  OAI22_X1 U2598 ( .A1(n1970), .A2(n1495), .B1(n1494), .B2(n2224), .ZN(n1206)
         );
  OAI22_X1 U2599 ( .A1(n2205), .A2(n1502), .B1(n2224), .B2(n1501), .ZN(n1213)
         );
  OAI22_X1 U2600 ( .A1(n1970), .A2(n1500), .B1(n2224), .B2(n1499), .ZN(n1211)
         );
  OAI22_X1 U2601 ( .A1(n2205), .A2(n1501), .B1(n1500), .B2(n2224), .ZN(n1212)
         );
  OAI22_X1 U2602 ( .A1(n1970), .A2(n1494), .B1(n2147), .B2(n1493), .ZN(n1205)
         );
  OAI22_X1 U2603 ( .A1(n1970), .A2(n1499), .B1(n1498), .B2(n2224), .ZN(n1210)
         );
  OAI22_X1 U2604 ( .A1(n1970), .A2(n1498), .B1(n2224), .B2(n1497), .ZN(n1209)
         );
  OAI22_X1 U2605 ( .A1(n2205), .A2(n1505), .B1(n1504), .B2(n2147), .ZN(n1216)
         );
  OAI22_X1 U2606 ( .A1(n2205), .A2(n1503), .B1(n1502), .B2(n2147), .ZN(n1214)
         );
  OAI22_X1 U2607 ( .A1(n2205), .A2(n1504), .B1(n1503), .B2(n2224), .ZN(n1215)
         );
  OAI22_X1 U2608 ( .A1(n2077), .A2(n1522), .B1(n1521), .B2(n2226), .ZN(n1232)
         );
  OAI22_X1 U2609 ( .A1(n2077), .A2(n1521), .B1(n2226), .B2(n1520), .ZN(n1231)
         );
  OAI22_X1 U2610 ( .A1(n2077), .A2(n1520), .B1(n1519), .B2(n2225), .ZN(n1230)
         );
  OAI22_X1 U2611 ( .A1(n2077), .A2(n1519), .B1(n2226), .B2(n1518), .ZN(n1229)
         );
  XNOR2_X1 U2612 ( .A(b[21]), .B(n2251), .ZN(n1534) );
  XNOR2_X1 U2613 ( .A(b[19]), .B(n2251), .ZN(n1536) );
  OAI22_X1 U2614 ( .A1(n2077), .A2(n1525), .B1(n2225), .B2(n1524), .ZN(n1235)
         );
  OAI22_X1 U2615 ( .A1(n2077), .A2(n1523), .B1(n2226), .B2(n1522), .ZN(n1233)
         );
  OAI22_X1 U2616 ( .A1(n1529), .A2(n2077), .B1(n2225), .B2(n1528), .ZN(n1239)
         );
  OAI22_X1 U2617 ( .A1(n2077), .A2(n1524), .B1(n1523), .B2(n2226), .ZN(n1234)
         );
  OAI22_X1 U2618 ( .A1(n2077), .A2(n1526), .B1(n1525), .B2(n2226), .ZN(n1236)
         );
  OAI22_X1 U2619 ( .A1(n2077), .A2(n1530), .B1(n1529), .B2(n2226), .ZN(n1240)
         );
  OAI22_X1 U2620 ( .A1(n2077), .A2(n1528), .B1(n1527), .B2(n2225), .ZN(n1238)
         );
  OAI22_X1 U2621 ( .A1(n1956), .A2(n2077), .B1(n2225), .B2(n1526), .ZN(n1237)
         );
  XNOR2_X1 U2622 ( .A(b[13]), .B(n2251), .ZN(n1542) );
  XNOR2_X1 U2623 ( .A(b[11]), .B(n2251), .ZN(n1544) );
  XNOR2_X1 U2624 ( .A(b[15]), .B(n2251), .ZN(n1540) );
  XNOR2_X1 U2625 ( .A(b[17]), .B(n2251), .ZN(n1538) );
  INV_X1 U2626 ( .A(n346), .ZN(n344) );
  AOI21_X1 U2627 ( .B1(n346), .B2(n2121), .A(n339), .ZN(n337) );
  NAND2_X1 U2628 ( .A1(n694), .A2(n689), .ZN(n378) );
  XNOR2_X1 U2629 ( .A(n410), .B(n308), .ZN(product[38]) );
  NAND2_X1 U2630 ( .A1(n761), .A2(n774), .ZN(n461) );
  XNOR2_X1 U2631 ( .A(n397), .B(n307), .ZN(product[39]) );
  OAI22_X1 U2632 ( .A1(n2215), .A2(n1637), .B1(n1636), .B2(n2154), .ZN(n1342)
         );
  OAI22_X1 U2633 ( .A1(n2073), .A2(n1636), .B1(n2233), .B2(n1635), .ZN(n1341)
         );
  OAI22_X1 U2634 ( .A1(n2073), .A2(n1634), .B1(n2233), .B2(n1633), .ZN(n1339)
         );
  OAI22_X1 U2635 ( .A1(n2073), .A2(n1635), .B1(n1634), .B2(n2154), .ZN(n1340)
         );
  OAI22_X1 U2636 ( .A1(n1931), .A2(n1639), .B1(n1638), .B2(n2154), .ZN(n1344)
         );
  OAI22_X1 U2637 ( .A1(n2073), .A2(n1640), .B1(n2232), .B2(n1639), .ZN(n1345)
         );
  OAI22_X1 U2638 ( .A1(n1930), .A2(n1638), .B1(n2233), .B2(n1637), .ZN(n1343)
         );
  OAI22_X1 U2639 ( .A1(n1930), .A2(n1642), .B1(n2232), .B2(n1641), .ZN(n1347)
         );
  OAI22_X1 U2640 ( .A1(n1931), .A2(n1633), .B1(n1632), .B2(n2154), .ZN(n772)
         );
  OAI22_X1 U2641 ( .A1(n2214), .A2(n1641), .B1(n1640), .B2(n2154), .ZN(n1346)
         );
  OAI22_X1 U2642 ( .A1(n2215), .A2(n1643), .B1(n1642), .B2(n2154), .ZN(n1348)
         );
  OAI22_X1 U2643 ( .A1(n2215), .A2(n2275), .B1(n1656), .B2(n2154), .ZN(n1188)
         );
  XNOR2_X1 U2644 ( .A(n388), .B(n306), .ZN(product[40]) );
  OAI22_X1 U2645 ( .A1(n2015), .A2(n1602), .B1(n2229), .B2(n1601), .ZN(n1309)
         );
  OAI22_X1 U2646 ( .A1(n2211), .A2(n1600), .B1(n2230), .B2(n1599), .ZN(n1307)
         );
  OAI22_X1 U2647 ( .A1(n2211), .A2(n1601), .B1(n1600), .B2(n2229), .ZN(n1308)
         );
  OAI22_X1 U2648 ( .A1(n2015), .A2(n1594), .B1(n2230), .B2(n1593), .ZN(n1301)
         );
  OAI22_X1 U2649 ( .A1(n2015), .A2(n1596), .B1(n2230), .B2(n1595), .ZN(n1303)
         );
  OAI22_X1 U2650 ( .A1(n2015), .A2(n1598), .B1(n2229), .B2(n1597), .ZN(n1305)
         );
  OAI22_X1 U2651 ( .A1(n2015), .A2(n1597), .B1(n1596), .B2(n2229), .ZN(n1304)
         );
  OAI22_X1 U2652 ( .A1(n2015), .A2(n1603), .B1(n1602), .B2(n2229), .ZN(n1310)
         );
  OAI22_X1 U2653 ( .A1(n2015), .A2(n1595), .B1(n1594), .B2(n2230), .ZN(n1302)
         );
  OAI22_X1 U2654 ( .A1(n2015), .A2(n1604), .B1(n2229), .B2(n1603), .ZN(n1311)
         );
  OAI22_X1 U2655 ( .A1(n2015), .A2(n1599), .B1(n1598), .B2(n2229), .ZN(n1306)
         );
  OAI22_X1 U2656 ( .A1(n2015), .A2(n1605), .B1(n1604), .B2(n2230), .ZN(n1312)
         );
  XNOR2_X1 U2657 ( .A(n379), .B(n305), .ZN(product[41]) );
  NAND2_X1 U2658 ( .A1(n775), .A2(n788), .ZN(n474) );
  NAND2_X1 U2659 ( .A1(n805), .A2(n820), .ZN(n496) );
  XNOR2_X1 U2660 ( .A(b[17]), .B(n2299), .ZN(n1763) );
  XNOR2_X1 U2661 ( .A(b[21]), .B(n2299), .ZN(n1759) );
  XNOR2_X1 U2662 ( .A(b[13]), .B(n2299), .ZN(n1767) );
  XNOR2_X1 U2663 ( .A(b[19]), .B(n2299), .ZN(n1761) );
  XNOR2_X1 U2664 ( .A(b[15]), .B(n2299), .ZN(n1765) );
  XNOR2_X1 U2665 ( .A(b[11]), .B(n2299), .ZN(n1769) );
  XNOR2_X1 U2666 ( .A(n370), .B(n304), .ZN(product[42]) );
  INV_X1 U2667 ( .A(n916), .ZN(n917) );
  XNOR2_X1 U2668 ( .A(n353), .B(n303), .ZN(product[43]) );
  OAI22_X1 U2669 ( .A1(n2220), .A2(n1733), .B1(n1732), .B2(n2238), .ZN(n916)
         );
  XOR2_X1 U2670 ( .A(n1946), .B(n321), .Z(product[25]) );
  OAI21_X1 U2671 ( .B1(n1947), .B2(n1975), .A(n535), .ZN(n533) );
  OAI21_X1 U2672 ( .B1(n1946), .B2(n487), .A(n488), .ZN(n486) );
  OAI21_X1 U2673 ( .B1(n1948), .B2(n463), .A(n464), .ZN(n462) );
  OAI21_X1 U2674 ( .B1(n1947), .B2(n2035), .A(n524), .ZN(n522) );
  OAI21_X1 U2675 ( .B1(n1946), .B2(n476), .A(n477), .ZN(n475) );
  OAI21_X1 U2676 ( .B1(n1947), .B2(n516), .A(n517), .ZN(n515) );
  OAI21_X1 U2677 ( .B1(n1948), .B2(n2158), .A(n2195), .ZN(n504) );
  OAI21_X1 U2678 ( .B1(n1948), .B2(n498), .A(n499), .ZN(n497) );
  OAI22_X1 U2679 ( .A1(n2149), .A2(n1727), .B1(n2061), .B2(n1726), .ZN(n1429)
         );
  OAI22_X1 U2680 ( .A1(n2149), .A2(n1720), .B1(n1719), .B2(n2061), .ZN(n1422)
         );
  OAI22_X1 U2681 ( .A1(n2149), .A2(n1721), .B1(n1969), .B2(n1720), .ZN(n1423)
         );
  OAI22_X1 U2682 ( .A1(n2149), .A2(n1726), .B1(n1725), .B2(n2061), .ZN(n1428)
         );
  OAI22_X1 U2683 ( .A1(n2149), .A2(n1730), .B1(n1729), .B2(n1969), .ZN(n1432)
         );
  OAI22_X1 U2684 ( .A1(n2149), .A2(n1725), .B1(n2061), .B2(n1724), .ZN(n1427)
         );
  OAI22_X1 U2685 ( .A1(n2149), .A2(n1723), .B1(n1969), .B2(n1722), .ZN(n1425)
         );
  OAI22_X1 U2686 ( .A1(n2149), .A2(n1728), .B1(n1727), .B2(n1969), .ZN(n1430)
         );
  OAI22_X1 U2687 ( .A1(n2149), .A2(n1722), .B1(n1721), .B2(n2061), .ZN(n1424)
         );
  OAI22_X1 U2688 ( .A1(n2149), .A2(n1729), .B1(n2061), .B2(n1728), .ZN(n1431)
         );
  OAI22_X1 U2689 ( .A1(n1957), .A2(n1719), .B1(n1969), .B2(n1718), .ZN(n1421)
         );
  OAI22_X1 U2690 ( .A1(n1957), .A2(n1724), .B1(n1723), .B2(n2061), .ZN(n1426)
         );
  XNOR2_X1 U2691 ( .A(b[15]), .B(n1968), .ZN(n1740) );
  XNOR2_X1 U2692 ( .A(b[21]), .B(n2295), .ZN(n1734) );
  XNOR2_X1 U2693 ( .A(b[19]), .B(n2295), .ZN(n1736) );
  XNOR2_X1 U2694 ( .A(b[11]), .B(n1968), .ZN(n1744) );
  XNOR2_X1 U2695 ( .A(b[17]), .B(n2295), .ZN(n1738) );
  XNOR2_X1 U2696 ( .A(b[13]), .B(n2295), .ZN(n1742) );
  INV_X1 U2697 ( .A(n325), .ZN(product[47]) );
  AOI21_X1 U2698 ( .B1(n423), .B2(n356), .A(n359), .ZN(n355) );
  NAND2_X1 U2699 ( .A1(n422), .A2(n356), .ZN(n354) );
  OAI22_X1 U2700 ( .A1(n1977), .A2(n1563), .B1(n2153), .B2(n1562), .ZN(n1271)
         );
  OAI22_X1 U2701 ( .A1(n1977), .A2(n1566), .B1(n1565), .B2(n2153), .ZN(n1274)
         );
  OAI22_X1 U2702 ( .A1(n2209), .A2(n1561), .B1(n2228), .B2(n1560), .ZN(n1269)
         );
  OAI22_X1 U2703 ( .A1(n2209), .A2(n1567), .B1(n2228), .B2(n1566), .ZN(n1275)
         );
  OAI22_X1 U2704 ( .A1(n2209), .A2(n1564), .B1(n1563), .B2(n2153), .ZN(n1272)
         );
  OAI22_X1 U2705 ( .A1(n1976), .A2(n1560), .B1(n1559), .B2(n2153), .ZN(n1268)
         );
  OAI22_X1 U2706 ( .A1(n1976), .A2(n2260), .B1(n1581), .B2(n2153), .ZN(n1185)
         );
  OAI22_X1 U2707 ( .A1(n2209), .A2(n1559), .B1(n2228), .B2(n1558), .ZN(n1267)
         );
  OAI22_X1 U2708 ( .A1(n2210), .A2(n1565), .B1(n2228), .B2(n1564), .ZN(n1273)
         );
  INV_X1 U2709 ( .A(n706), .ZN(n707) );
  OAI22_X1 U2710 ( .A1(n2209), .A2(n1562), .B1(n1561), .B2(n2153), .ZN(n1270)
         );
  OAI22_X1 U2711 ( .A1(n2209), .A2(n1568), .B1(n1567), .B2(n2153), .ZN(n1276)
         );
  OAI22_X1 U2712 ( .A1(n1976), .A2(n1558), .B1(n1557), .B2(n2153), .ZN(n706)
         );
  XNOR2_X1 U2713 ( .A(n342), .B(n302), .ZN(product[44]) );
  OAI21_X1 U2714 ( .B1(n2189), .B2(n326), .A(n327), .ZN(n325) );
  OAI21_X1 U2715 ( .B1(n2188), .B2(n411), .A(n412), .ZN(n410) );
  OAI21_X1 U2716 ( .B1(n2188), .B2(n431), .A(n432), .ZN(n430) );
  OAI21_X1 U2717 ( .B1(n2189), .B2(n354), .A(n355), .ZN(n353) );
  OAI21_X1 U2718 ( .B1(n2181), .B2(n420), .A(n421), .ZN(n419) );
  OAI21_X1 U2719 ( .B1(n2189), .B2(n398), .A(n399), .ZN(n397) );
  OAI21_X1 U2720 ( .B1(n2181), .B2(n438), .A(n439), .ZN(n437) );
  OAI21_X1 U2721 ( .B1(n2181), .B2(n343), .A(n344), .ZN(n342) );
  OAI21_X1 U2722 ( .B1(n2188), .B2(n389), .A(n390), .ZN(n388) );
  OAI21_X1 U2723 ( .B1(n301), .B2(n371), .A(n372), .ZN(n370) );
  OAI21_X1 U2724 ( .B1(n301), .B2(n380), .A(n381), .ZN(n379) );
  OAI22_X1 U2725 ( .A1(n2095), .A2(n1691), .B1(n1690), .B2(n2235), .ZN(n1394)
         );
  OAI22_X1 U2726 ( .A1(n2096), .A2(n1686), .B1(n2236), .B2(n1685), .ZN(n1389)
         );
  OAI22_X1 U2727 ( .A1(n2095), .A2(n1689), .B1(n1688), .B2(n2236), .ZN(n1392)
         );
  OAI22_X1 U2728 ( .A1(n2219), .A2(n1690), .B1(n2235), .B2(n1689), .ZN(n1393)
         );
  OAI22_X1 U2729 ( .A1(n2218), .A2(n1687), .B1(n1686), .B2(n2236), .ZN(n1390)
         );
  OAI22_X1 U2730 ( .A1(n2096), .A2(n1692), .B1(n2235), .B2(n1691), .ZN(n1395)
         );
  OAI22_X1 U2731 ( .A1(n2004), .A2(n1685), .B1(n1684), .B2(n2236), .ZN(n1388)
         );
  OAI22_X1 U2732 ( .A1(n2004), .A2(n1688), .B1(n2236), .B2(n1687), .ZN(n1391)
         );
  INV_X1 U2733 ( .A(n836), .ZN(n837) );
  OAI22_X1 U2734 ( .A1(n2095), .A2(n1684), .B1(n2236), .B2(n1683), .ZN(n1387)
         );
  OAI22_X1 U2735 ( .A1(n2218), .A2(n2287), .B1(n1706), .B2(n2236), .ZN(n1190)
         );
  OAI22_X1 U2736 ( .A1(n2219), .A2(n1693), .B1(n1692), .B2(n1986), .ZN(n1396)
         );
  OAI22_X1 U2737 ( .A1(n2219), .A2(n1683), .B1(n1682), .B2(n1986), .ZN(n836)
         );
  INV_X2 U2738 ( .A(n2137), .ZN(n2211) );
  INV_X1 U2739 ( .A(n2194), .ZN(n2233) );
  INV_X1 U2740 ( .A(n2094), .ZN(n2236) );
  INV_X1 U2741 ( .A(n2250), .ZN(n2248) );
  INV_X1 U2742 ( .A(a[21]), .ZN(n2249) );
  INV_X1 U2743 ( .A(a[21]), .ZN(n2250) );
  INV_X1 U2744 ( .A(n2255), .ZN(n2253) );
  INV_X1 U2745 ( .A(a[19]), .ZN(n2254) );
  INV_X1 U2746 ( .A(a[19]), .ZN(n2255) );
  INV_X1 U2747 ( .A(n2261), .ZN(n2259) );
  INV_X1 U2748 ( .A(a[17]), .ZN(n2260) );
  INV_X1 U2749 ( .A(a[17]), .ZN(n2261) );
  INV_X1 U2750 ( .A(n2265), .ZN(n2264) );
  INV_X1 U2751 ( .A(a[15]), .ZN(n2265) );
  INV_X1 U2752 ( .A(a[15]), .ZN(n2266) );
  INV_X1 U2753 ( .A(n2271), .ZN(n2269) );
  INV_X1 U2754 ( .A(a[13]), .ZN(n2270) );
  INV_X1 U2755 ( .A(a[13]), .ZN(n2271) );
  INV_X1 U2756 ( .A(n2276), .ZN(n2274) );
  INV_X1 U2757 ( .A(a[11]), .ZN(n2275) );
  INV_X1 U2758 ( .A(a[11]), .ZN(n2276) );
  INV_X1 U2759 ( .A(n2281), .ZN(n2280) );
  INV_X1 U2760 ( .A(a[9]), .ZN(n2281) );
  INV_X1 U2761 ( .A(a[9]), .ZN(n2282) );
  INV_X1 U2762 ( .A(n2288), .ZN(n2286) );
  INV_X1 U2763 ( .A(a[7]), .ZN(n2287) );
  INV_X1 U2764 ( .A(a[7]), .ZN(n2288) );
  INV_X1 U2765 ( .A(n2294), .ZN(n2292) );
  INV_X1 U2766 ( .A(a[5]), .ZN(n2293) );
  INV_X1 U2767 ( .A(n1978), .ZN(n2294) );
  INV_X1 U2768 ( .A(n2298), .ZN(n2296) );
  INV_X1 U2769 ( .A(n1983), .ZN(n2297) );
  INV_X1 U2770 ( .A(a[3]), .ZN(n2298) );
  INV_X1 U2771 ( .A(n2304), .ZN(n2302) );
  INV_X1 U2772 ( .A(a[1]), .ZN(n2303) );
  INV_X1 U2773 ( .A(a[1]), .ZN(n2304) );
  INV_X2 U2774 ( .A(b[0]), .ZN(n2305) );
endmodule


module iir_filter_DW_mult_tc_3 ( a, b, product );
  input [23:0] a;
  input [23:0] b;
  output [47:0] product;
  wire   n251, n277, n281, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n325, n326, n327, n332, n333, n334, n335, n336, n337, n339,
         n341, n342, n343, n344, n345, n346, n347, n348, n350, n352, n353,
         n354, n355, n356, n359, n360, n361, n362, n363, n364, n365, n367,
         n369, n370, n371, n372, n376, n378, n379, n380, n381, n382, n383,
         n384, n387, n388, n389, n390, n394, n396, n397, n398, n399, n400,
         n401, n402, n405, n407, n409, n410, n411, n412, n416, n418, n419,
         n420, n421, n422, n423, n426, n427, n428, n429, n430, n431, n432,
         n434, n435, n436, n437, n438, n439, n445, n450, n451, n452, n453,
         n454, n455, n456, n457, n459, n461, n462, n463, n464, n465, n466,
         n467, n468, n472, n474, n475, n476, n477, n478, n479, n480, n481,
         n483, n486, n487, n488, n489, n490, n492, n495, n496, n497, n498,
         n499, n502, n503, n504, n505, n506, n507, n508, n511, n512, n513,
         n514, n515, n516, n517, n519, n520, n521, n522, n524, n525, n526,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n550, n551, n552, n553, n554,
         n555, n558, n559, n560, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n581, n582, n583, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n609, n610,
         n611, n620, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n643, n644, n645, n646, n657, n661,
         n662, n663, n667, n668, n670, n673, n674, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1806, n1807, n1809, n1810, n1817, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317;

  FA_X1 U546 ( .A(n1195), .B(n682), .CI(n1218), .CO(n678), .S(n679) );
  FA_X1 U547 ( .A(n683), .B(n1196), .CI(n686), .CO(n680), .S(n681) );
  FA_X1 U549 ( .A(n690), .B(n1242), .CI(n687), .CO(n684), .S(n685) );
  FA_X1 U550 ( .A(n1219), .B(n692), .CI(n1197), .CO(n686), .S(n687) );
  FA_X1 U551 ( .A(n691), .B(n698), .CI(n696), .CO(n688), .S(n689) );
  FA_X1 U552 ( .A(n1198), .B(n1220), .CI(n693), .CO(n690), .S(n691) );
  FA_X1 U554 ( .A(n702), .B(n699), .CI(n697), .CO(n694), .S(n695) );
  FA_X1 U555 ( .A(n1266), .B(n1243), .CI(n704), .CO(n696), .S(n697) );
  FA_X1 U556 ( .A(n1221), .B(n1199), .CI(n706), .CO(n698), .S(n699) );
  FA_X1 U557 ( .A(n710), .B(n712), .CI(n703), .CO(n700), .S(n701) );
  FA_X1 U558 ( .A(n714), .B(n1244), .CI(n705), .CO(n702), .S(n703) );
  FA_X1 U559 ( .A(n1222), .B(n1200), .CI(n707), .CO(n704), .S(n705) );
  FA_X1 U561 ( .A(n718), .B(n713), .CI(n711), .CO(n708), .S(n709) );
  FA_X1 U562 ( .A(n715), .B(n722), .CI(n720), .CO(n710), .S(n711) );
  FA_X1 U563 ( .A(n1245), .B(n1223), .CI(n1290), .CO(n712), .S(n713) );
  FA_X1 U564 ( .A(n1267), .B(n1201), .CI(n724), .CO(n714), .S(n715) );
  FA_X1 U565 ( .A(n728), .B(n721), .CI(n719), .CO(n716), .S(n717) );
  FA_X1 U566 ( .A(n723), .B(n732), .CI(n730), .CO(n718), .S(n719) );
  FA_X1 U567 ( .A(n1202), .B(n1246), .CI(n734), .CO(n720), .S(n721) );
  FA_X1 U568 ( .A(n1268), .B(n1224), .CI(n725), .CO(n722), .S(n723) );
  FA_X1 U570 ( .A(n738), .B(n731), .CI(n729), .CO(n726), .S(n727) );
  FA_X1 U571 ( .A(n735), .B(n733), .CI(n740), .CO(n728), .S(n729) );
  FA_X1 U572 ( .A(n744), .B(n1314), .CI(n742), .CO(n730), .S(n731) );
  FA_X1 U573 ( .A(n1225), .B(n1291), .CI(n1269), .CO(n732), .S(n733) );
  FA_X1 U574 ( .A(n746), .B(n1203), .CI(n1247), .CO(n734), .S(n735) );
  FA_X1 U575 ( .A(n750), .B(n741), .CI(n739), .CO(n736), .S(n737) );
  FA_X1 U576 ( .A(n754), .B(n745), .CI(n752), .CO(n738), .S(n739) );
  FA_X1 U577 ( .A(n756), .B(n758), .CI(n743), .CO(n740), .S(n741) );
  FA_X1 U578 ( .A(n1226), .B(n1204), .CI(n1270), .CO(n742), .S(n743) );
  FA_X1 U579 ( .A(n1292), .B(n1248), .CI(n747), .CO(n744), .S(n745) );
  FA_X1 U581 ( .A(n762), .B(n753), .CI(n751), .CO(n748), .S(n749) );
  FA_X1 U582 ( .A(n755), .B(n766), .CI(n764), .CO(n750), .S(n751) );
  FA_X1 U583 ( .A(n757), .B(n768), .CI(n759), .CO(n752), .S(n753) );
  FA_X1 U584 ( .A(n1338), .B(n1271), .CI(n770), .CO(n754), .S(n755) );
  FA_X1 U585 ( .A(n1249), .B(n1293), .CI(n1315), .CO(n756), .S(n757) );
  FA_X1 U586 ( .A(n772), .B(n1205), .CI(n1227), .CO(n758), .S(n759) );
  FA_X1 U587 ( .A(n776), .B(n765), .CI(n763), .CO(n760), .S(n761) );
  FA_X1 U588 ( .A(n767), .B(n780), .CI(n778), .CO(n762), .S(n763) );
  FA_X1 U589 ( .A(n771), .B(n769), .CI(n782), .CO(n764), .S(n765) );
  FA_X1 U590 ( .A(n786), .B(n1228), .CI(n784), .CO(n766), .S(n767) );
  FA_X1 U591 ( .A(n1294), .B(n1206), .CI(n1272), .CO(n768), .S(n769) );
  FA_X1 U592 ( .A(n1316), .B(n1250), .CI(n773), .CO(n770), .S(n771) );
  FA_X1 U594 ( .A(n777), .B(n779), .CI(n790), .CO(n774), .S(n775) );
  FA_X1 U595 ( .A(n781), .B(n794), .CI(n792), .CO(n776), .S(n777) );
  FA_X1 U596 ( .A(n796), .B(n787), .CI(n783), .CO(n778), .S(n779) );
  FA_X1 U597 ( .A(n798), .B(n800), .CI(n785), .CO(n780), .S(n781) );
  FA_X1 U598 ( .A(n1339), .B(n1229), .CI(n1362), .CO(n782), .S(n783) );
  FA_X1 U599 ( .A(n1273), .B(n1317), .CI(n1295), .CO(n784), .S(n785) );
  FA_X1 U600 ( .A(n1251), .B(n1207), .CI(n802), .CO(n786), .S(n787) );
  FA_X1 U601 ( .A(n806), .B(n793), .CI(n791), .CO(n788), .S(n789) );
  FA_X1 U602 ( .A(n795), .B(n810), .CI(n808), .CO(n790), .S(n791) );
  FA_X1 U604 ( .A(n814), .B(n816), .CI(n799), .CO(n794), .S(n795) );
  FA_X1 U606 ( .A(n1208), .B(n1318), .CI(n1230), .CO(n798), .S(n799) );
  FA_X1 U607 ( .A(n1340), .B(n1252), .CI(n803), .CO(n800), .S(n801) );
  FA_X1 U609 ( .A(n822), .B(n809), .CI(n807), .CO(n804), .S(n805) );
  FA_X1 U610 ( .A(n811), .B(n826), .CI(n824), .CO(n806), .S(n807) );
  FA_X1 U611 ( .A(n828), .B(n819), .CI(n813), .CO(n808), .S(n809) );
  FA_X1 U612 ( .A(n815), .B(n832), .CI(n817), .CO(n810), .S(n811) );
  FA_X1 U614 ( .A(n1319), .B(n1253), .CI(n1341), .CO(n814), .S(n815) );
  FA_X1 U615 ( .A(n1231), .B(n1297), .CI(n1275), .CO(n816), .S(n817) );
  FA_X1 U616 ( .A(n1363), .B(n1209), .CI(n2222), .CO(n818), .S(n819) );
  FA_X1 U617 ( .A(n840), .B(n825), .CI(n823), .CO(n820), .S(n821) );
  FA_X1 U619 ( .A(n846), .B(n848), .CI(n829), .CO(n824), .S(n825) );
  FA_X1 U620 ( .A(n835), .B(n831), .CI(n833), .CO(n826), .S(n827) );
  FA_X1 U621 ( .A(n852), .B(n854), .CI(n850), .CO(n828), .S(n829) );
  FA_X1 U622 ( .A(n1254), .B(n1320), .CI(n1298), .CO(n830), .S(n831) );
  FA_X1 U623 ( .A(n1232), .B(n1364), .CI(n1342), .CO(n832), .S(n833) );
  FA_X1 U626 ( .A(n843), .B(n858), .CI(n841), .CO(n838), .S(n839) );
  FA_X1 U627 ( .A(n845), .B(n847), .CI(n860), .CO(n840), .S(n841) );
  FA_X1 U629 ( .A(n855), .B(n853), .CI(n866), .CO(n844), .S(n845) );
  FA_X1 U630 ( .A(n868), .B(n870), .CI(n851), .CO(n846), .S(n847) );
  FA_X1 U631 ( .A(n1410), .B(n1365), .CI(n872), .CO(n848), .S(n849) );
  FA_X1 U632 ( .A(n1299), .B(n1277), .CI(n1343), .CO(n850), .S(n851) );
  FA_X1 U633 ( .A(n874), .B(n1255), .CI(n1321), .CO(n852), .S(n853) );
  FA_X1 U634 ( .A(n1211), .B(n1387), .CI(n1233), .CO(n854), .S(n855) );
  FA_X1 U638 ( .A(n888), .B(n873), .CI(n886), .CO(n862), .S(n863) );
  FA_X1 U639 ( .A(n869), .B(n890), .CI(n871), .CO(n864), .S(n865) );
  FA_X1 U640 ( .A(n894), .B(n1300), .CI(n892), .CO(n866), .S(n867) );
  FA_X1 U641 ( .A(n1234), .B(n1322), .CI(n1256), .CO(n868), .S(n869) );
  FA_X1 U642 ( .A(n1212), .B(n1366), .CI(n1344), .CO(n870), .S(n871) );
  FA_X1 U643 ( .A(n1388), .B(n1278), .CI(n875), .CO(n872), .S(n873) );
  FA_X1 U645 ( .A(n898), .B(n881), .CI(n879), .CO(n876), .S(n877) );
  FA_X1 U646 ( .A(n883), .B(n885), .CI(n900), .CO(n878), .S(n879) );
  FA_X1 U648 ( .A(n906), .B(n893), .CI(n889), .CO(n882), .S(n883) );
  FA_X1 U650 ( .A(n910), .B(n912), .CI(n914), .CO(n886), .S(n887) );
  FA_X1 U651 ( .A(n1367), .B(n1389), .CI(n1434), .CO(n888), .S(n889) );
  FA_X1 U652 ( .A(n1257), .B(n1301), .CI(n1345), .CO(n890), .S(n891) );
  FA_X1 U653 ( .A(n2214), .B(n1323), .CI(n1279), .CO(n892), .S(n893) );
  FA_X1 U654 ( .A(n1235), .B(n1411), .CI(n1213), .CO(n894), .S(n895) );
  FA_X1 U656 ( .A(n903), .B(n924), .CI(n922), .CO(n898), .S(n899) );
  FA_X1 U657 ( .A(n907), .B(n926), .CI(n905), .CO(n900), .S(n901) );
  FA_X1 U658 ( .A(n909), .B(n930), .CI(n928), .CO(n902), .S(n903) );
  FA_X1 U659 ( .A(n913), .B(n911), .CI(n915), .CO(n904), .S(n905) );
  FA_X1 U660 ( .A(n932), .B(n936), .CI(n934), .CO(n906), .S(n907) );
  FA_X1 U661 ( .A(n1368), .B(n1390), .CI(n938), .CO(n908), .S(n909) );
  FA_X1 U662 ( .A(n1324), .B(n1346), .CI(n1280), .CO(n910), .S(n911) );
  FA_X1 U663 ( .A(n1258), .B(n1412), .CI(n1236), .CO(n912), .S(n913) );
  FA_X1 U664 ( .A(n1302), .B(n1214), .CI(n917), .CO(n914), .S(n915) );
  FA_X1 U666 ( .A(n942), .B(n923), .CI(n921), .CO(n918), .S(n919) );
  FA_X1 U667 ( .A(n925), .B(n927), .CI(n944), .CO(n920), .S(n921) );
  FA_X1 U668 ( .A(n929), .B(n948), .CI(n946), .CO(n922), .S(n923) );
  FA_X1 U669 ( .A(n950), .B(n935), .CI(n931), .CO(n924), .S(n925) );
  FA_X1 U671 ( .A(n954), .B(n956), .CI(n958), .CO(n928), .S(n929) );
  FA_X1 U672 ( .A(n939), .B(n960), .CI(n1458), .CO(n930), .S(n931) );
  FA_X1 U673 ( .A(n1325), .B(n1435), .CI(n1413), .CO(n932), .S(n933) );
  FA_X1 U674 ( .A(n1281), .B(n1369), .CI(n1391), .CO(n934), .S(n935) );
  FA_X1 U678 ( .A(n964), .B(n945), .CI(n943), .CO(n940), .S(n941) );
  FA_X1 U679 ( .A(n947), .B(n949), .CI(n966), .CO(n942), .S(n943) );
  FA_X1 U680 ( .A(n951), .B(n970), .CI(n968), .CO(n944), .S(n945) );
  FA_X1 U681 ( .A(n972), .B(n959), .CI(n953), .CO(n946), .S(n947) );
  FA_X1 U682 ( .A(n955), .B(n974), .CI(n957), .CO(n948), .S(n949) );
  FA_X1 U683 ( .A(n976), .B(n980), .CI(n978), .CO(n950), .S(n951) );
  FA_X1 U684 ( .A(n1326), .B(n1392), .CI(n961), .CO(n952), .S(n953) );
  FA_X1 U686 ( .A(n1459), .B(n1370), .CI(n1436), .CO(n956), .S(n957) );
  FA_X1 U687 ( .A(n1260), .B(n1348), .CI(n1182), .CO(n958), .S(n959) );
  HA_X1 U688 ( .A(n1238), .B(n1216), .CO(n960), .S(n961) );
  FA_X1 U689 ( .A(n984), .B(n967), .CI(n965), .CO(n962), .S(n963) );
  FA_X1 U690 ( .A(n969), .B(n971), .CI(n986), .CO(n964), .S(n965) );
  FA_X1 U691 ( .A(n973), .B(n990), .CI(n988), .CO(n966), .S(n967) );
  FA_X1 U693 ( .A(n977), .B(n998), .CI(n979), .CO(n970), .S(n971) );
  FA_X1 U696 ( .A(n1305), .B(n1327), .CI(n1437), .CO(n976), .S(n977) );
  FA_X1 U697 ( .A(n1460), .B(n1371), .CI(n1283), .CO(n978), .S(n979) );
  FA_X1 U698 ( .A(n1261), .B(n1349), .CI(n1239), .CO(n980), .S(n981) );
  FA_X1 U699 ( .A(n1004), .B(n987), .CI(n985), .CO(n982), .S(n983) );
  FA_X1 U700 ( .A(n989), .B(n991), .CI(n1006), .CO(n984), .S(n985) );
  FA_X1 U701 ( .A(n993), .B(n1010), .CI(n1008), .CO(n986), .S(n987) );
  FA_X1 U702 ( .A(n999), .B(n997), .CI(n1012), .CO(n988), .S(n989) );
  FA_X1 U703 ( .A(n1014), .B(n1016), .CI(n995), .CO(n990), .S(n991) );
  FA_X1 U704 ( .A(n1001), .B(n1394), .CI(n1018), .CO(n992), .S(n993) );
  FA_X1 U707 ( .A(n1183), .B(n1350), .CI(n1461), .CO(n998), .S(n999) );
  FA_X1 U709 ( .A(n1022), .B(n1007), .CI(n1005), .CO(n1002), .S(n1003) );
  FA_X1 U710 ( .A(n1009), .B(n1011), .CI(n1024), .CO(n1004), .S(n1005) );
  FA_X1 U711 ( .A(n1013), .B(n1028), .CI(n1026), .CO(n1006), .S(n1007) );
  FA_X1 U712 ( .A(n1019), .B(n1015), .CI(n1017), .CO(n1008), .S(n1009) );
  FA_X1 U713 ( .A(n1030), .B(n1034), .CI(n1241), .CO(n1010), .S(n1011) );
  FA_X1 U714 ( .A(n1036), .B(n1439), .CI(n1032), .CO(n1012), .S(n1013) );
  FA_X1 U715 ( .A(n1417), .B(n1462), .CI(n1395), .CO(n1014), .S(n1015) );
  FA_X1 U716 ( .A(n1307), .B(n1373), .CI(n1329), .CO(n1016), .S(n1017) );
  FA_X1 U717 ( .A(n1263), .B(n1351), .CI(n1285), .CO(n1018), .S(n1019) );
  FA_X1 U718 ( .A(n1040), .B(n1025), .CI(n1023), .CO(n1020), .S(n1021) );
  FA_X1 U719 ( .A(n1027), .B(n1044), .CI(n1042), .CO(n1022), .S(n1023) );
  FA_X1 U720 ( .A(n1046), .B(n1035), .CI(n1029), .CO(n1024), .S(n1025) );
  FA_X1 U721 ( .A(n1031), .B(n1048), .CI(n1033), .CO(n1026), .S(n1027) );
  FA_X1 U722 ( .A(n1052), .B(n1037), .CI(n1050), .CO(n1028), .S(n1029) );
  FA_X1 U723 ( .A(n1418), .B(n1440), .CI(n1352), .CO(n1030), .S(n1031) );
  FA_X1 U725 ( .A(n1308), .B(n1374), .CI(n1184), .CO(n1034), .S(n1035) );
  HA_X1 U726 ( .A(n1264), .B(n1286), .CO(n1036), .S(n1037) );
  FA_X1 U727 ( .A(n1056), .B(n1043), .CI(n1041), .CO(n1038), .S(n1039) );
  FA_X1 U728 ( .A(n1058), .B(n1047), .CI(n1045), .CO(n1040), .S(n1041) );
  FA_X1 U730 ( .A(n1049), .B(n1265), .CI(n1051), .CO(n1044), .S(n1045) );
  FA_X1 U731 ( .A(n1064), .B(n1068), .CI(n1066), .CO(n1046), .S(n1047) );
  FA_X1 U732 ( .A(n1397), .B(n1441), .CI(n1419), .CO(n1048), .S(n1049) );
  FA_X1 U733 ( .A(n1331), .B(n1353), .CI(n1375), .CO(n1050), .S(n1051) );
  FA_X1 U734 ( .A(n1287), .B(n1464), .CI(n1309), .CO(n1052), .S(n1053) );
  FA_X1 U735 ( .A(n1072), .B(n1059), .CI(n1057), .CO(n1054), .S(n1055) );
  FA_X1 U736 ( .A(n1074), .B(n1063), .CI(n1061), .CO(n1056), .S(n1057) );
  FA_X1 U737 ( .A(n1067), .B(n1065), .CI(n1076), .CO(n1058), .S(n1059) );
  FA_X1 U739 ( .A(n1398), .B(n1420), .CI(n1069), .CO(n1062), .S(n1063) );
  FA_X1 U740 ( .A(n1442), .B(n1354), .CI(n1332), .CO(n1064), .S(n1065) );
  FA_X1 U741 ( .A(n1465), .B(n1376), .CI(n1185), .CO(n1066), .S(n1067) );
  HA_X1 U742 ( .A(n1288), .B(n1310), .CO(n1068), .S(n1069) );
  FA_X1 U743 ( .A(n1086), .B(n1075), .CI(n1073), .CO(n1070), .S(n1071) );
  FA_X1 U744 ( .A(n1088), .B(n1090), .CI(n1077), .CO(n1072), .S(n1073) );
  FA_X1 U745 ( .A(n1083), .B(n1081), .CI(n1079), .CO(n1074), .S(n1075) );
  FA_X1 U746 ( .A(n1092), .B(n1094), .CI(n1289), .CO(n1076), .S(n1077) );
  FA_X1 U747 ( .A(n1399), .B(n1421), .CI(n1096), .CO(n1078), .S(n1079) );
  FA_X1 U748 ( .A(n1355), .B(n1443), .CI(n1377), .CO(n1080), .S(n1081) );
  FA_X1 U749 ( .A(n1311), .B(n1466), .CI(n1333), .CO(n1082), .S(n1083) );
  FA_X1 U750 ( .A(n1100), .B(n1089), .CI(n1087), .CO(n1084), .S(n1085) );
  FA_X1 U751 ( .A(n1102), .B(n1104), .CI(n1091), .CO(n1086), .S(n1087) );
  FA_X1 U752 ( .A(n1093), .B(n1106), .CI(n1095), .CO(n1088), .S(n1089) );
  FA_X1 U753 ( .A(n1097), .B(n1422), .CI(n1108), .CO(n1090), .S(n1091) );
  FA_X1 U754 ( .A(n1444), .B(n1356), .CI(n1378), .CO(n1092), .S(n1093) );
  FA_X1 U755 ( .A(n1186), .B(n1400), .CI(n1467), .CO(n1094), .S(n1095) );
  HA_X1 U756 ( .A(n1312), .B(n1334), .CO(n1096), .S(n1097) );
  FA_X1 U757 ( .A(n1103), .B(n1112), .CI(n1101), .CO(n1098), .S(n1099) );
  FA_X1 U758 ( .A(n1114), .B(n1109), .CI(n1105), .CO(n1100), .S(n1101) );
  FA_X1 U759 ( .A(n1313), .B(n1116), .CI(n1107), .CO(n1102), .S(n1103) );
  FA_X1 U760 ( .A(n1120), .B(n1423), .CI(n1118), .CO(n1104), .S(n1105) );
  FA_X1 U761 ( .A(n1379), .B(n1445), .CI(n1401), .CO(n1106), .S(n1107) );
  FA_X1 U762 ( .A(n1335), .B(n1468), .CI(n1357), .CO(n1108), .S(n1109) );
  FA_X1 U763 ( .A(n1124), .B(n1115), .CI(n1113), .CO(n1110), .S(n1111) );
  FA_X1 U764 ( .A(n1119), .B(n1117), .CI(n1126), .CO(n1112), .S(n1113) );
  FA_X1 U765 ( .A(n1130), .B(n1121), .CI(n1128), .CO(n1114), .S(n1115) );
  FA_X1 U766 ( .A(n1424), .B(n1469), .CI(n1446), .CO(n1116), .S(n1117) );
  FA_X1 U767 ( .A(n1380), .B(n1402), .CI(n1187), .CO(n1118), .S(n1119) );
  HA_X1 U768 ( .A(n1336), .B(n1358), .CO(n1120), .S(n1121) );
  FA_X1 U769 ( .A(n1127), .B(n1134), .CI(n1125), .CO(n1122), .S(n1123) );
  FA_X1 U770 ( .A(n1131), .B(n1129), .CI(n1136), .CO(n1124), .S(n1125) );
  FA_X1 U771 ( .A(n1138), .B(n1140), .CI(n1337), .CO(n1126), .S(n1127) );
  FA_X1 U772 ( .A(n1403), .B(n1447), .CI(n1425), .CO(n1128), .S(n1129) );
  FA_X1 U773 ( .A(n1359), .B(n1470), .CI(n1381), .CO(n1130), .S(n1131) );
  FA_X1 U774 ( .A(n1144), .B(n1137), .CI(n1135), .CO(n1132), .S(n1133) );
  FA_X1 U775 ( .A(n1146), .B(n1148), .CI(n1139), .CO(n1134), .S(n1135) );
  FA_X1 U776 ( .A(n1404), .B(n1448), .CI(n1141), .CO(n1136), .S(n1137) );
  FA_X1 U777 ( .A(n1471), .B(n1426), .CI(n1188), .CO(n1138), .S(n1139) );
  HA_X1 U778 ( .A(n1360), .B(n1382), .CO(n1140), .S(n1141) );
  FA_X1 U779 ( .A(n1152), .B(n1147), .CI(n1145), .CO(n1142), .S(n1143) );
  FA_X1 U780 ( .A(n1361), .B(n1154), .CI(n1149), .CO(n1144), .S(n1145) );
  FA_X1 U781 ( .A(n1427), .B(n1449), .CI(n1156), .CO(n1146), .S(n1147) );
  FA_X1 U782 ( .A(n1383), .B(n1472), .CI(n1405), .CO(n1148), .S(n1149) );
  FA_X1 U783 ( .A(n1160), .B(n1155), .CI(n1153), .CO(n1150), .S(n1151) );
  FA_X1 U784 ( .A(n1157), .B(n1473), .CI(n1162), .CO(n1152), .S(n1153) );
  FA_X1 U785 ( .A(n1450), .B(n1428), .CI(n1189), .CO(n1154), .S(n1155) );
  HA_X1 U786 ( .A(n1384), .B(n1406), .CO(n1156), .S(n1157) );
  FA_X1 U787 ( .A(n1163), .B(n1385), .CI(n1164), .CO(n1158), .S(n1159) );
  FA_X1 U788 ( .A(n1168), .B(n1429), .CI(n1166), .CO(n1160), .S(n1161) );
  FA_X1 U789 ( .A(n1451), .B(n1474), .CI(n1407), .CO(n1162), .S(n1163) );
  FA_X1 U790 ( .A(n1172), .B(n1169), .CI(n1167), .CO(n1164), .S(n1165) );
  FA_X1 U791 ( .A(n1452), .B(n1475), .CI(n1190), .CO(n1166), .S(n1167) );
  HA_X1 U792 ( .A(n1408), .B(n1430), .CO(n1168), .S(n1169) );
  FA_X1 U793 ( .A(n1409), .B(n1176), .CI(n1173), .CO(n1170), .S(n1171) );
  FA_X1 U794 ( .A(n1476), .B(n1453), .CI(n1431), .CO(n1172), .S(n1173) );
  FA_X1 U795 ( .A(n1191), .B(n1454), .CI(n1177), .CO(n1174), .S(n1175) );
  HA_X1 U796 ( .A(n1432), .B(n1477), .CO(n1176), .S(n1177) );
  FA_X1 U797 ( .A(n1455), .B(n1478), .CI(n1180), .CO(n1178), .S(n1179) );
  HA_X1 U798 ( .A(n1456), .B(n1479), .CO(n1180), .S(n1181) );
  BUF_X1 U1448 ( .A(n568), .Z(n2060) );
  CLKBUF_X1 U1449 ( .A(n277), .Z(n2054) );
  XNOR2_X1 U1450 ( .A(n2106), .B(n1929), .ZN(product[34]) );
  AND2_X1 U1451 ( .A1(n663), .A2(n439), .ZN(n1929) );
  INV_X4 U1452 ( .A(n2030), .ZN(n2300) );
  INV_X2 U1453 ( .A(n2055), .ZN(n2056) );
  XNOR2_X1 U1454 ( .A(a[21]), .B(a[22]), .ZN(n1930) );
  INV_X2 U1455 ( .A(n1930), .ZN(n2205) );
  OR2_X4 U1456 ( .A1(n2146), .A2(n2149), .ZN(n2108) );
  BUF_X1 U1457 ( .A(n2099), .Z(n1949) );
  CLKBUF_X1 U1458 ( .A(n251), .Z(n2257) );
  BUF_X4 U1459 ( .A(n251), .Z(n2258) );
  INV_X1 U1460 ( .A(a[15]), .ZN(n1931) );
  CLKBUF_X1 U1461 ( .A(n2061), .Z(n2010) );
  INV_X1 U1462 ( .A(n2145), .ZN(n2231) );
  INV_X1 U1463 ( .A(n1964), .ZN(n2150) );
  NAND3_X1 U1464 ( .A1(n2077), .A2(n2078), .A3(n2079), .ZN(n884) );
  OR2_X1 U1465 ( .A1(n709), .A2(n716), .ZN(n2123) );
  NOR2_X1 U1466 ( .A1(n727), .A2(n736), .ZN(n428) );
  NAND3_X1 U1467 ( .A1(n2001), .A2(n2002), .A3(n2003), .ZN(n896) );
  AND2_X1 U1468 ( .A1(n1193), .A2(n1481), .ZN(n1932) );
  OR2_X1 U1469 ( .A1(n1457), .A2(n1480), .ZN(n1933) );
  OR2_X1 U1470 ( .A1(n1179), .A2(n1433), .ZN(n1934) );
  AND2_X1 U1471 ( .A1(n1151), .A2(n1158), .ZN(n1935) );
  AND2_X1 U1472 ( .A1(n1987), .A2(n1262), .ZN(n1936) );
  INV_X1 U1473 ( .A(n2167), .ZN(n2004) );
  AND2_X1 U1474 ( .A1(n1457), .A2(n1480), .ZN(n1937) );
  AND2_X1 U1475 ( .A1(n1179), .A2(n1433), .ZN(n1938) );
  AND2_X1 U1476 ( .A1(n1123), .A2(n1132), .ZN(n1939) );
  AND2_X1 U1477 ( .A1(n1133), .A2(n1142), .ZN(n1940) );
  AND2_X1 U1478 ( .A1(n1055), .A2(n1070), .ZN(n1941) );
  AND2_X1 U1479 ( .A1(n1021), .A2(n1038), .ZN(n1942) );
  OR2_X1 U1480 ( .A1(n1151), .A2(n1158), .ZN(n1943) );
  OR2_X1 U1481 ( .A1(n963), .A2(n982), .ZN(n1944) );
  CLKBUF_X1 U1482 ( .A(n2099), .Z(n2159) );
  CLKBUF_X1 U1483 ( .A(a[3]), .Z(n1945) );
  XNOR2_X1 U1484 ( .A(n551), .B(n1946), .ZN(product[23]) );
  AND2_X1 U1485 ( .A1(n674), .A2(n550), .ZN(n1946) );
  XNOR2_X1 U1486 ( .A(n560), .B(n1947), .ZN(product[22]) );
  AND2_X1 U1487 ( .A1(n1944), .A2(n559), .ZN(n1947) );
  NOR2_X1 U1488 ( .A1(n1003), .A2(n1020), .ZN(n1948) );
  XNOR2_X1 U1489 ( .A(a[0]), .B(n2051), .ZN(n1817) );
  BUF_X2 U1490 ( .A(n2099), .Z(n1950) );
  BUF_X1 U1491 ( .A(n536), .Z(n1951) );
  BUF_X1 U1492 ( .A(n536), .Z(n1953) );
  BUF_X1 U1493 ( .A(n536), .Z(n1952) );
  BUF_X1 U1494 ( .A(n506), .Z(n2091) );
  INV_X1 U1495 ( .A(n2056), .ZN(n1954) );
  INV_X2 U1496 ( .A(n2149), .ZN(n2253) );
  INV_X1 U1497 ( .A(n2167), .ZN(n1956) );
  INV_X1 U1498 ( .A(n2167), .ZN(n1955) );
  INV_X1 U1499 ( .A(n2202), .ZN(n2038) );
  CLKBUF_X3 U1500 ( .A(n277), .Z(n2191) );
  XNOR2_X1 U1501 ( .A(n996), .B(n1957), .ZN(n973) );
  XNOR2_X1 U1502 ( .A(n994), .B(n1217), .ZN(n1957) );
  XNOR2_X1 U1503 ( .A(n1958), .B(n1284), .ZN(n997) );
  XNOR2_X1 U1504 ( .A(n1438), .B(n1372), .ZN(n1958) );
  XNOR2_X1 U1505 ( .A(n899), .B(n1959), .ZN(n897) );
  XNOR2_X1 U1506 ( .A(n920), .B(n901), .ZN(n1959) );
  AND2_X1 U1507 ( .A1(n2257), .A2(n1817), .ZN(n2142) );
  INV_X1 U1508 ( .A(n2194), .ZN(n1961) );
  INV_X1 U1509 ( .A(n2194), .ZN(n1960) );
  INV_X1 U1510 ( .A(n2194), .ZN(n2243) );
  INV_X2 U1511 ( .A(n2037), .ZN(n2280) );
  OR2_X1 U1512 ( .A1(n2176), .A2(n2144), .ZN(n1962) );
  OR2_X1 U1513 ( .A1(n2176), .A2(n2144), .ZN(n277) );
  CLKBUF_X1 U1514 ( .A(a[10]), .Z(n1963) );
  OR2_X2 U1515 ( .A1(n2204), .A2(n2151), .ZN(n1964) );
  INV_X2 U1516 ( .A(n2205), .ZN(n2236) );
  XOR2_X1 U1517 ( .A(a[6]), .B(n2057), .Z(n1997) );
  CLKBUF_X1 U1518 ( .A(n2135), .Z(n2164) );
  INV_X1 U1519 ( .A(n2172), .ZN(n2266) );
  INV_X1 U1520 ( .A(n2172), .ZN(n2267) );
  CLKBUF_X1 U1521 ( .A(a[5]), .Z(n1965) );
  OR2_X1 U1522 ( .A1(n2151), .A2(n2204), .ZN(n1966) );
  CLKBUF_X3 U1523 ( .A(n1966), .Z(n2162) );
  XOR2_X1 U1524 ( .A(a[20]), .B(n2270), .Z(n1967) );
  INV_X1 U1525 ( .A(a[19]), .ZN(n2172) );
  INV_X1 U1526 ( .A(n2194), .ZN(n2244) );
  INV_X1 U1527 ( .A(n2147), .ZN(n1969) );
  INV_X2 U1528 ( .A(n2147), .ZN(n1968) );
  INV_X1 U1529 ( .A(n2147), .ZN(n2228) );
  NOR2_X1 U1530 ( .A1(n2206), .A2(n896), .ZN(n1970) );
  NAND3_X1 U1531 ( .A1(n2026), .A2(n2027), .A3(n2028), .ZN(n1971) );
  CLKBUF_X1 U1532 ( .A(n879), .Z(n2047) );
  XNOR2_X1 U1533 ( .A(a[12]), .B(n1993), .ZN(n1973) );
  XNOR2_X1 U1534 ( .A(a[12]), .B(n1993), .ZN(n1972) );
  XNOR2_X1 U1535 ( .A(a[12]), .B(n1993), .ZN(n2141) );
  INV_X1 U1536 ( .A(n1988), .ZN(n1974) );
  OR2_X1 U1537 ( .A1(n789), .A2(n804), .ZN(n1975) );
  OR2_X1 U1538 ( .A1(n2155), .A2(n2174), .ZN(n2042) );
  XNOR2_X1 U1539 ( .A(a[4]), .B(n1965), .ZN(n2146) );
  INV_X1 U1540 ( .A(n2241), .ZN(n1976) );
  CLKBUF_X3 U1541 ( .A(n2135), .Z(n2165) );
  INV_X1 U1542 ( .A(n281), .ZN(n1977) );
  OR2_X2 U1543 ( .A1(n1997), .A2(n2143), .ZN(n281) );
  INV_X1 U1544 ( .A(n492), .ZN(n1978) );
  INV_X1 U1545 ( .A(n2148), .ZN(n1979) );
  CLKBUF_X1 U1546 ( .A(n877), .Z(n1980) );
  CLKBUF_X1 U1547 ( .A(n1955), .Z(n1981) );
  AND2_X1 U1548 ( .A1(n1817), .A2(n2257), .ZN(n1982) );
  BUF_X1 U1549 ( .A(n2143), .Z(n1983) );
  XOR2_X1 U1550 ( .A(a[6]), .B(a[5]), .Z(n2143) );
  INV_X1 U1551 ( .A(n2202), .ZN(n1984) );
  INV_X1 U1552 ( .A(n2000), .ZN(n1985) );
  INV_X1 U1553 ( .A(n2148), .ZN(n2226) );
  INV_X1 U1554 ( .A(n2255), .ZN(n1986) );
  OAI22_X1 U1555 ( .A1(n1530), .A2(n1956), .B1(n1529), .B2(n2056), .ZN(n1987)
         );
  CLKBUF_X1 U1556 ( .A(n2204), .Z(n1988) );
  XNOR2_X1 U1557 ( .A(a[14]), .B(n2277), .ZN(n1810) );
  XOR2_X1 U1558 ( .A(a[12]), .B(n2037), .Z(n2157) );
  INV_X1 U1559 ( .A(n2282), .ZN(n2279) );
  CLKBUF_X1 U1560 ( .A(n1970), .Z(n1989) );
  NOR2_X1 U1561 ( .A1(n2206), .A2(n896), .ZN(n531) );
  INV_X1 U1562 ( .A(n2148), .ZN(n1991) );
  INV_X1 U1563 ( .A(n2148), .ZN(n1990) );
  INV_X1 U1564 ( .A(n2148), .ZN(n2225) );
  INV_X1 U1565 ( .A(n2277), .ZN(n2275) );
  INV_X2 U1566 ( .A(n1982), .ZN(n1992) );
  INV_X1 U1567 ( .A(n2142), .ZN(n2234) );
  INV_X1 U1568 ( .A(a[11]), .ZN(n1993) );
  XNOR2_X2 U1569 ( .A(n2301), .B(a[4]), .ZN(n2149) );
  INV_X1 U1570 ( .A(a[17]), .ZN(n1995) );
  INV_X1 U1571 ( .A(a[17]), .ZN(n1994) );
  INV_X1 U1572 ( .A(n2275), .ZN(n1996) );
  BUF_X1 U1573 ( .A(n1303), .Z(n1998) );
  INV_X1 U1574 ( .A(n2246), .ZN(n1999) );
  INV_X1 U1575 ( .A(n1930), .ZN(n2000) );
  INV_X1 U1576 ( .A(n2204), .ZN(n2249) );
  XOR2_X1 U1577 ( .A(a[7]), .B(a[8]), .Z(n2204) );
  XOR2_X1 U1578 ( .A(a[10]), .B(a[9]), .Z(n2169) );
  NAND2_X1 U1579 ( .A1(n899), .A2(n920), .ZN(n2001) );
  NAND2_X1 U1580 ( .A1(n899), .A2(n901), .ZN(n2002) );
  NAND2_X1 U1581 ( .A1(n920), .A2(n901), .ZN(n2003) );
  INV_X1 U1582 ( .A(n2167), .ZN(n2005) );
  OR2_X1 U1583 ( .A1(n502), .A2(n2188), .ZN(n2006) );
  XNOR2_X1 U1584 ( .A(a[16]), .B(a[15]), .ZN(n2085) );
  INV_X2 U1585 ( .A(n2298), .ZN(n2297) );
  INV_X2 U1586 ( .A(n2142), .ZN(n2235) );
  XNOR2_X1 U1587 ( .A(n1396), .B(n2007), .ZN(n1033) );
  XNOR2_X1 U1588 ( .A(n1463), .B(n1330), .ZN(n2007) );
  XNOR2_X1 U1589 ( .A(n859), .B(n2008), .ZN(n857) );
  XNOR2_X1 U1590 ( .A(n878), .B(n861), .ZN(n2008) );
  AND2_X2 U1591 ( .A1(n1809), .A2(n2085), .ZN(n2148) );
  XOR2_X1 U1592 ( .A(a[18]), .B(n2172), .Z(n2155) );
  XNOR2_X1 U1593 ( .A(a[8]), .B(a[9]), .ZN(n2151) );
  INV_X1 U1594 ( .A(a[9]), .ZN(n2290) );
  INV_X1 U1595 ( .A(n2265), .ZN(n2264) );
  CLKBUF_X3 U1596 ( .A(a[21]), .Z(n2039) );
  INV_X1 U1597 ( .A(n2098), .ZN(n2009) );
  XOR2_X1 U1598 ( .A(n904), .B(n887), .Z(n2011) );
  XOR2_X1 U1599 ( .A(n902), .B(n2011), .Z(n881) );
  NAND2_X1 U1600 ( .A1(n902), .A2(n904), .ZN(n2012) );
  NAND2_X1 U1601 ( .A1(n902), .A2(n887), .ZN(n2013) );
  NAND2_X1 U1602 ( .A1(n904), .A2(n887), .ZN(n2014) );
  NAND3_X1 U1603 ( .A1(n2012), .A2(n2013), .A3(n2014), .ZN(n880) );
  OR2_X1 U1604 ( .A1(n983), .A2(n1002), .ZN(n2015) );
  INV_X2 U1605 ( .A(n2295), .ZN(n2293) );
  OR2_X1 U1606 ( .A1(n897), .A2(n918), .ZN(n2016) );
  XOR2_X1 U1607 ( .A(n1274), .B(n1296), .Z(n2017) );
  XOR2_X1 U1608 ( .A(n2017), .B(n818), .Z(n797) );
  XOR2_X1 U1609 ( .A(n812), .B(n801), .Z(n2018) );
  XOR2_X1 U1610 ( .A(n2018), .B(n797), .Z(n793) );
  NAND2_X1 U1611 ( .A1(n1274), .A2(n1296), .ZN(n2019) );
  NAND2_X1 U1612 ( .A1(n1274), .A2(n818), .ZN(n2020) );
  NAND2_X1 U1613 ( .A1(n1296), .A2(n818), .ZN(n2021) );
  NAND3_X1 U1614 ( .A1(n2019), .A2(n2020), .A3(n2021), .ZN(n796) );
  NAND2_X1 U1615 ( .A1(n812), .A2(n801), .ZN(n2022) );
  NAND2_X1 U1616 ( .A1(n812), .A2(n797), .ZN(n2023) );
  NAND2_X1 U1617 ( .A1(n801), .A2(n797), .ZN(n2024) );
  NAND3_X1 U1618 ( .A1(n2022), .A2(n2023), .A3(n2024), .ZN(n792) );
  XOR2_X1 U1619 ( .A(n1080), .B(n1082), .Z(n2025) );
  XOR2_X1 U1620 ( .A(n1078), .B(n2025), .Z(n1061) );
  NAND2_X1 U1621 ( .A1(n1078), .A2(n1080), .ZN(n2026) );
  NAND2_X1 U1622 ( .A1(n1078), .A2(n1082), .ZN(n2027) );
  NAND2_X1 U1623 ( .A1(n1080), .A2(n1082), .ZN(n2028) );
  NAND3_X1 U1624 ( .A1(n2026), .A2(n2027), .A3(n2028), .ZN(n1060) );
  INV_X1 U1625 ( .A(n2191), .ZN(n2029) );
  INV_X1 U1626 ( .A(a[3]), .ZN(n2030) );
  XOR2_X1 U1627 ( .A(n849), .B(n864), .Z(n2031) );
  XOR2_X1 U1628 ( .A(n862), .B(n2031), .Z(n843) );
  NAND2_X1 U1629 ( .A1(n862), .A2(n849), .ZN(n2032) );
  NAND2_X1 U1630 ( .A1(n862), .A2(n864), .ZN(n2033) );
  NAND2_X1 U1631 ( .A1(n849), .A2(n864), .ZN(n2034) );
  NAND3_X1 U1632 ( .A1(n2032), .A2(n2033), .A3(n2034), .ZN(n842) );
  BUF_X1 U1633 ( .A(n495), .Z(n2035) );
  INV_X1 U1634 ( .A(a[3]), .ZN(n2301) );
  OAI21_X1 U1635 ( .B1(n535), .B2(n1989), .A(n532), .ZN(n2036) );
  INV_X1 U1636 ( .A(a[13]), .ZN(n2037) );
  INV_X2 U1637 ( .A(n1972), .ZN(n2246) );
  XOR2_X1 U1638 ( .A(a[1]), .B(a[2]), .Z(n2144) );
  INV_X1 U1639 ( .A(a[5]), .ZN(n2298) );
  NOR2_X1 U1640 ( .A1(n963), .A2(n982), .ZN(n2040) );
  NOR2_X1 U1641 ( .A1(n963), .A2(n982), .ZN(n558) );
  OR2_X2 U1642 ( .A1(n2155), .A2(n2174), .ZN(n2041) );
  OR2_X1 U1643 ( .A1(n2155), .A2(n2174), .ZN(n2062) );
  XOR2_X1 U1644 ( .A(n863), .B(n882), .Z(n2043) );
  XOR2_X1 U1645 ( .A(n880), .B(n2043), .Z(n859) );
  NAND2_X1 U1646 ( .A1(n880), .A2(n863), .ZN(n2044) );
  NAND2_X1 U1647 ( .A1(n880), .A2(n882), .ZN(n2045) );
  NAND2_X1 U1648 ( .A1(n863), .A2(n882), .ZN(n2046) );
  NAND3_X1 U1649 ( .A1(n2044), .A2(n2045), .A3(n2046), .ZN(n858) );
  INV_X1 U1650 ( .A(n2085), .ZN(n2202) );
  XOR2_X1 U1651 ( .A(n1240), .B(n1262), .Z(n1001) );
  BUF_X1 U1652 ( .A(n553), .Z(n2069) );
  XNOR2_X2 U1653 ( .A(a[18]), .B(n2274), .ZN(n2174) );
  INV_X2 U1654 ( .A(n2174), .ZN(n2240) );
  NAND2_X1 U1655 ( .A1(n859), .A2(n878), .ZN(n2048) );
  NAND2_X1 U1656 ( .A1(n859), .A2(n861), .ZN(n2049) );
  NAND2_X1 U1657 ( .A1(n878), .A2(n861), .ZN(n2050) );
  NAND3_X1 U1658 ( .A1(n2048), .A2(n2049), .A3(n2050), .ZN(n856) );
  INV_X1 U1659 ( .A(a[1]), .ZN(n2052) );
  INV_X1 U1660 ( .A(a[1]), .ZN(n2051) );
  CLKBUF_X1 U1661 ( .A(n505), .Z(n2053) );
  INV_X1 U1662 ( .A(n2062), .ZN(n2154) );
  NOR2_X2 U1663 ( .A1(n558), .A2(n563), .ZN(n552) );
  INV_X1 U1664 ( .A(n1967), .ZN(n2055) );
  INV_X1 U1665 ( .A(a[7]), .ZN(n2057) );
  OR2_X2 U1666 ( .A1(n2157), .A2(n2141), .ZN(n2059) );
  OR2_X2 U1667 ( .A1(n2157), .A2(n2141), .ZN(n2058) );
  OR2_X1 U1668 ( .A1(n2157), .A2(n1972), .ZN(n2107) );
  INV_X2 U1669 ( .A(n1973), .ZN(n2245) );
  INV_X1 U1670 ( .A(n2265), .ZN(n2263) );
  XNOR2_X1 U1671 ( .A(a[20]), .B(n2172), .ZN(n2203) );
  XNOR2_X1 U1672 ( .A(a[20]), .B(n2175), .ZN(n1807) );
  INV_X1 U1673 ( .A(a[7]), .ZN(n2295) );
  XOR2_X1 U1674 ( .A(n2286), .B(n1963), .Z(n2153) );
  INV_X1 U1675 ( .A(a[11]), .ZN(n2286) );
  INV_X1 U1676 ( .A(n2099), .ZN(n2152) );
  NOR2_X1 U1677 ( .A1(n940), .A2(n919), .ZN(n2061) );
  NOR2_X1 U1678 ( .A1(n919), .A2(n940), .ZN(n542) );
  NAND2_X1 U1679 ( .A1(n1330), .A2(n1396), .ZN(n2063) );
  NAND2_X1 U1680 ( .A1(n1463), .A2(n1396), .ZN(n2064) );
  NAND2_X1 U1681 ( .A1(n1330), .A2(n1463), .ZN(n2065) );
  NAND3_X1 U1682 ( .A1(n2063), .A2(n2064), .A3(n2065), .ZN(n1032) );
  INV_X1 U1683 ( .A(n674), .ZN(n2066) );
  OR2_X1 U1684 ( .A1(n2229), .A2(n1693), .ZN(n2067) );
  OR2_X1 U1685 ( .A1(n1692), .A2(n2251), .ZN(n2068) );
  NAND2_X1 U1686 ( .A1(n2067), .A2(n2068), .ZN(n1396) );
  NOR2_X1 U1687 ( .A1(n941), .A2(n962), .ZN(n547) );
  INV_X2 U1688 ( .A(n2298), .ZN(n2296) );
  XNOR2_X1 U1689 ( .A(a[16]), .B(n1994), .ZN(n1809) );
  INV_X1 U1690 ( .A(n1995), .ZN(n2272) );
  INV_X1 U1691 ( .A(a[17]), .ZN(n2274) );
  INV_X1 U1692 ( .A(n2230), .ZN(n2071) );
  INV_X1 U1693 ( .A(n2230), .ZN(n2070) );
  INV_X1 U1694 ( .A(n1977), .ZN(n2229) );
  XNOR2_X1 U1695 ( .A(n2072), .B(n975), .ZN(n969) );
  XNOR2_X1 U1696 ( .A(n992), .B(n981), .ZN(n2072) );
  NAND2_X1 U1697 ( .A1(n1438), .A2(n1284), .ZN(n2073) );
  NAND2_X1 U1698 ( .A1(n1284), .A2(n1372), .ZN(n2074) );
  NAND2_X1 U1699 ( .A1(n1438), .A2(n1372), .ZN(n2075) );
  NAND3_X1 U1700 ( .A1(n2073), .A2(n2074), .A3(n2075), .ZN(n996) );
  XOR2_X1 U1701 ( .A(n891), .B(n908), .Z(n2076) );
  XOR2_X1 U1702 ( .A(n2076), .B(n895), .Z(n885) );
  NAND2_X1 U1703 ( .A1(n891), .A2(n908), .ZN(n2077) );
  NAND2_X1 U1704 ( .A1(n891), .A2(n895), .ZN(n2078) );
  NAND2_X1 U1705 ( .A1(n908), .A2(n895), .ZN(n2079) );
  XOR2_X1 U1706 ( .A(n867), .B(n865), .Z(n2080) );
  XOR2_X1 U1707 ( .A(n2080), .B(n884), .Z(n861) );
  NAND2_X1 U1708 ( .A1(n865), .A2(n867), .ZN(n2081) );
  NAND2_X1 U1709 ( .A1(n867), .A2(n884), .ZN(n2082) );
  NAND2_X1 U1710 ( .A1(n865), .A2(n884), .ZN(n2083) );
  NAND3_X1 U1711 ( .A1(n2081), .A2(n2082), .A3(n2083), .ZN(n860) );
  OR2_X1 U1712 ( .A1(n839), .A2(n856), .ZN(n2084) );
  INV_X2 U1713 ( .A(n2202), .ZN(n2242) );
  INV_X1 U1714 ( .A(n2167), .ZN(n2224) );
  OR2_X2 U1715 ( .A1(n788), .A2(n775), .ZN(n2192) );
  INV_X1 U1716 ( .A(n2290), .ZN(n2287) );
  INV_X1 U1717 ( .A(n2016), .ZN(n2086) );
  XOR2_X1 U1718 ( .A(n1304), .B(n1414), .Z(n2087) );
  XOR2_X1 U1719 ( .A(n2087), .B(n1282), .Z(n955) );
  NAND2_X1 U1720 ( .A1(n1282), .A2(n1304), .ZN(n2088) );
  NAND2_X1 U1721 ( .A1(n1282), .A2(n1414), .ZN(n2089) );
  NAND2_X1 U1722 ( .A1(n1304), .A2(n1414), .ZN(n2090) );
  NAND3_X1 U1723 ( .A1(n2088), .A2(n2089), .A3(n2090), .ZN(n954) );
  XOR2_X1 U1724 ( .A(n1062), .B(n1053), .Z(n2092) );
  XOR2_X1 U1725 ( .A(n1971), .B(n2092), .Z(n1043) );
  NAND2_X1 U1726 ( .A1(n1971), .A2(n1062), .ZN(n2093) );
  NAND2_X1 U1727 ( .A1(n1060), .A2(n1053), .ZN(n2094) );
  NAND2_X1 U1728 ( .A1(n1062), .A2(n1053), .ZN(n2095) );
  NAND3_X1 U1729 ( .A1(n2093), .A2(n2094), .A3(n2095), .ZN(n1042) );
  AOI21_X1 U1730 ( .B1(n581), .B2(n567), .A(n2060), .ZN(n2096) );
  XNOR2_X1 U1731 ( .A(n2097), .B(n1936), .ZN(n975) );
  XNOR2_X1 U1732 ( .A(n1393), .B(n1415), .ZN(n2097) );
  AOI21_X1 U1733 ( .B1(n581), .B2(n567), .A(n568), .ZN(n566) );
  INV_X1 U1734 ( .A(n2059), .ZN(n2156) );
  OR2_X1 U1735 ( .A1(n534), .A2(n1989), .ZN(n2098) );
  OR2_X2 U1736 ( .A1(n2153), .A2(n2169), .ZN(n2099) );
  NOR2_X1 U1737 ( .A1(n839), .A2(n856), .ZN(n513) );
  NAND2_X1 U1738 ( .A1(n1393), .A2(n1415), .ZN(n2100) );
  NAND2_X1 U1739 ( .A1(n1393), .A2(n1936), .ZN(n2101) );
  NAND2_X1 U1740 ( .A1(n1415), .A2(n1936), .ZN(n2102) );
  NAND3_X1 U1741 ( .A1(n2100), .A2(n2101), .A3(n2102), .ZN(n974) );
  NAND2_X1 U1742 ( .A1(n992), .A2(n981), .ZN(n2103) );
  NAND2_X1 U1743 ( .A1(n981), .A2(n975), .ZN(n2104) );
  NAND2_X1 U1744 ( .A1(n992), .A2(n975), .ZN(n2105) );
  NAND3_X1 U1745 ( .A1(n2103), .A2(n2104), .A3(n2105), .ZN(n968) );
  AND2_X2 U1746 ( .A1(n2220), .A2(n2221), .ZN(n2106) );
  AND2_X2 U1747 ( .A1(n2220), .A2(n2221), .ZN(n301) );
  INV_X2 U1748 ( .A(n2057), .ZN(n2292) );
  XOR2_X1 U1749 ( .A(n827), .B(n844), .Z(n2109) );
  XOR2_X1 U1750 ( .A(n842), .B(n2109), .Z(n823) );
  NAND2_X1 U1751 ( .A1(n842), .A2(n827), .ZN(n2110) );
  NAND2_X1 U1752 ( .A1(n842), .A2(n844), .ZN(n2111) );
  NAND2_X1 U1753 ( .A1(n827), .A2(n844), .ZN(n2112) );
  NAND3_X1 U1754 ( .A1(n2110), .A2(n2111), .A3(n2112), .ZN(n822) );
  BUF_X2 U1755 ( .A(n2099), .Z(n2160) );
  XNOR2_X1 U1756 ( .A(n544), .B(n2113), .ZN(product[24]) );
  AND2_X1 U1757 ( .A1(n673), .A2(n543), .ZN(n2113) );
  NAND2_X1 U1758 ( .A1(n2122), .A2(n2123), .ZN(n402) );
  NOR2_X1 U1759 ( .A1(n695), .A2(n700), .ZN(n384) );
  AND2_X1 U1760 ( .A1(n1143), .A2(n1150), .ZN(n2114) );
  OR2_X1 U1761 ( .A1(n1143), .A2(n1150), .ZN(n2115) );
  XNOR2_X1 U1762 ( .A(n2130), .B(n1998), .ZN(n937) );
  XOR2_X1 U1763 ( .A(n2116), .B(n2138), .Z(n835) );
  XOR2_X1 U1764 ( .A(n1276), .B(n1210), .Z(n2116) );
  XOR2_X1 U1765 ( .A(n1416), .B(n2117), .Z(n995) );
  XOR2_X1 U1766 ( .A(n1306), .B(n1328), .Z(n2117) );
  OR2_X1 U1767 ( .A1(n679), .A2(n680), .ZN(n2134) );
  OR2_X1 U1768 ( .A1(n685), .A2(n688), .ZN(n2131) );
  INV_X2 U1769 ( .A(n2261), .ZN(n2259) );
  NAND2_X1 U1770 ( .A1(n465), .A2(n507), .ZN(n463) );
  INV_X1 U1771 ( .A(n505), .ZN(n507) );
  NOR2_X1 U1772 ( .A1(n2006), .A2(n467), .ZN(n465) );
  XNOR2_X1 U1773 ( .A(n522), .B(n319), .ZN(product[27]) );
  NAND2_X1 U1774 ( .A1(n478), .A2(n507), .ZN(n476) );
  NAND2_X1 U1775 ( .A1(n507), .A2(n668), .ZN(n498) );
  NAND2_X1 U1776 ( .A1(n662), .A2(n436), .ZN(n311) );
  OAI21_X1 U1777 ( .B1(n421), .B2(n402), .A(n405), .ZN(n401) );
  INV_X1 U1778 ( .A(n435), .ZN(n662) );
  NOR2_X1 U1779 ( .A1(n420), .A2(n402), .ZN(n400) );
  NAND2_X1 U1780 ( .A1(n667), .A2(n496), .ZN(n316) );
  AOI21_X1 U1781 ( .B1(n565), .B2(n2015), .A(n562), .ZN(n560) );
  AOI21_X1 U1782 ( .B1(n565), .B2(n545), .A(n546), .ZN(n544) );
  AOI21_X1 U1783 ( .B1(n2036), .B2(n670), .A(n519), .ZN(n517) );
  AOI21_X1 U1784 ( .B1(n662), .B2(n445), .A(n434), .ZN(n432) );
  INV_X1 U1785 ( .A(n436), .ZN(n434) );
  INV_X1 U1786 ( .A(n439), .ZN(n445) );
  XNOR2_X1 U1787 ( .A(n486), .B(n315), .ZN(product[31]) );
  NAND2_X1 U1788 ( .A1(n1975), .A2(n481), .ZN(n315) );
  XNOR2_X1 U1789 ( .A(n504), .B(n317), .ZN(product[29]) );
  XNOR2_X1 U1790 ( .A(n515), .B(n318), .ZN(product[28]) );
  NAND2_X1 U1791 ( .A1(n2084), .A2(n514), .ZN(n318) );
  NOR2_X1 U1792 ( .A1(n402), .A2(n360), .ZN(n356) );
  OAI21_X1 U1793 ( .B1(n492), .B2(n467), .A(n468), .ZN(n466) );
  INV_X1 U1794 ( .A(n481), .ZN(n483) );
  INV_X1 U1795 ( .A(n564), .ZN(n562) );
  INV_X1 U1796 ( .A(n438), .ZN(n663) );
  INV_X1 U1797 ( .A(n2036), .ZN(n524) );
  INV_X1 U1798 ( .A(n552), .ZN(n554) );
  INV_X1 U1799 ( .A(n382), .ZN(n380) );
  NOR2_X1 U1800 ( .A1(n789), .A2(n804), .ZN(n480) );
  AOI21_X1 U1801 ( .B1(n2123), .B2(n416), .A(n407), .ZN(n405) );
  INV_X1 U1802 ( .A(n409), .ZN(n407) );
  OR2_X1 U1803 ( .A1(n761), .A2(n774), .ZN(n2118) );
  AND2_X1 U1804 ( .A1(n1039), .A2(n1054), .ZN(n2119) );
  NAND2_X1 U1805 ( .A1(n2122), .A2(n418), .ZN(n309) );
  NOR2_X1 U1806 ( .A1(n384), .A2(n364), .ZN(n362) );
  NOR2_X1 U1807 ( .A1(n435), .A2(n428), .ZN(n426) );
  INV_X1 U1808 ( .A(n418), .ZN(n416) );
  INV_X1 U1809 ( .A(n383), .ZN(n381) );
  NAND2_X1 U1810 ( .A1(n2123), .A2(n409), .ZN(n308) );
  NAND2_X1 U1811 ( .A1(n422), .A2(n2122), .ZN(n411) );
  NAND2_X1 U1812 ( .A1(n657), .A2(n387), .ZN(n306) );
  INV_X1 U1813 ( .A(n384), .ZN(n657) );
  NAND2_X1 U1814 ( .A1(n2125), .A2(n396), .ZN(n307) );
  NAND2_X1 U1815 ( .A1(n661), .A2(n429), .ZN(n310) );
  NAND2_X1 U1816 ( .A1(n963), .A2(n982), .ZN(n559) );
  AOI21_X1 U1817 ( .B1(n423), .B2(n2122), .A(n416), .ZN(n412) );
  OAI21_X1 U1818 ( .B1(n535), .B2(n1970), .A(n532), .ZN(n526) );
  XNOR2_X1 U1819 ( .A(n533), .B(n320), .ZN(product[26]) );
  NOR2_X1 U1820 ( .A1(n389), .A2(n384), .ZN(n382) );
  INV_X1 U1821 ( .A(n396), .ZN(n394) );
  NAND2_X1 U1822 ( .A1(n362), .A2(n2125), .ZN(n360) );
  INV_X1 U1823 ( .A(n378), .ZN(n376) );
  NAND2_X1 U1824 ( .A1(n983), .A2(n1002), .ZN(n564) );
  OR2_X1 U1825 ( .A1(n1039), .A2(n1054), .ZN(n2120) );
  NAND2_X1 U1826 ( .A1(n1003), .A2(n1020), .ZN(n570) );
  OR2_X1 U1827 ( .A1(n1055), .A2(n1070), .ZN(n2121) );
  OR2_X2 U1828 ( .A1(n717), .A2(n726), .ZN(n2122) );
  INV_X1 U1829 ( .A(n352), .ZN(n350) );
  OAI21_X1 U1830 ( .B1(n638), .B2(n636), .A(n637), .ZN(n635) );
  OAI21_X1 U1831 ( .B1(n631), .B2(n634), .A(n632), .ZN(n630) );
  AND2_X1 U1832 ( .A1(n1111), .A2(n1122), .ZN(n2124) );
  OR2_X2 U1833 ( .A1(n701), .A2(n708), .ZN(n2125) );
  NAND2_X1 U1834 ( .A1(n2127), .A2(n2131), .ZN(n364) );
  NOR2_X1 U1835 ( .A1(n1099), .A2(n1110), .ZN(n597) );
  OR2_X1 U1836 ( .A1(n1133), .A2(n1142), .ZN(n2126) );
  NAND2_X1 U1837 ( .A1(n2131), .A2(n369), .ZN(n304) );
  NAND2_X1 U1838 ( .A1(n2134), .A2(n341), .ZN(n302) );
  NAND2_X1 U1839 ( .A1(n2133), .A2(n352), .ZN(n303) );
  NAND2_X1 U1840 ( .A1(n695), .A2(n700), .ZN(n387) );
  OAI21_X1 U1841 ( .B1(n405), .B2(n360), .A(n361), .ZN(n359) );
  AOI21_X1 U1842 ( .B1(n362), .B2(n394), .A(n363), .ZN(n361) );
  OAI21_X1 U1843 ( .B1(n364), .B2(n387), .A(n365), .ZN(n363) );
  AOI21_X1 U1844 ( .B1(n376), .B2(n2131), .A(n367), .ZN(n365) );
  NAND2_X1 U1845 ( .A1(n701), .A2(n708), .ZN(n396) );
  OR2_X1 U1846 ( .A1(n694), .A2(n689), .ZN(n2127) );
  INV_X1 U1847 ( .A(n369), .ZN(n367) );
  OR2_X1 U1848 ( .A1(n1111), .A2(n1122), .ZN(n2128) );
  AOI21_X1 U1849 ( .B1(n2126), .B2(n2114), .A(n1940), .ZN(n611) );
  NOR2_X1 U1850 ( .A1(n590), .A2(n592), .ZN(n588) );
  NOR2_X1 U1851 ( .A1(n1085), .A2(n1098), .ZN(n592) );
  OR2_X1 U1852 ( .A1(n1123), .A2(n1132), .ZN(n2129) );
  NAND2_X1 U1853 ( .A1(n1099), .A2(n1110), .ZN(n598) );
  NAND2_X1 U1854 ( .A1(n2115), .A2(n2126), .ZN(n610) );
  XNOR2_X1 U1855 ( .A(n1259), .B(n1347), .ZN(n2130) );
  AOI21_X1 U1856 ( .B1(n643), .B2(n1934), .A(n1938), .ZN(n638) );
  OAI21_X1 U1857 ( .B1(n646), .B2(n644), .A(n645), .ZN(n643) );
  NOR2_X1 U1858 ( .A1(n1165), .A2(n1170), .ZN(n631) );
  NAND2_X1 U1859 ( .A1(n678), .A2(n677), .ZN(n335) );
  INV_X1 U1860 ( .A(n341), .ZN(n339) );
  NOR2_X1 U1861 ( .A1(n1175), .A2(n1178), .ZN(n636) );
  XNOR2_X1 U1862 ( .A(n2132), .B(n834), .ZN(n813) );
  XNOR2_X1 U1863 ( .A(n1386), .B(n830), .ZN(n2132) );
  OR2_X2 U1864 ( .A1(n681), .A2(n684), .ZN(n2133) );
  NAND2_X1 U1865 ( .A1(n681), .A2(n684), .ZN(n352) );
  NAND2_X1 U1866 ( .A1(n679), .A2(n680), .ZN(n341) );
  NOR2_X1 U1867 ( .A1(n1171), .A2(n1174), .ZN(n633) );
  NOR2_X1 U1868 ( .A1(n1159), .A2(n1161), .ZN(n626) );
  NAND2_X1 U1869 ( .A1(n1175), .A2(n1178), .ZN(n637) );
  NAND2_X1 U1870 ( .A1(n1806), .A2(n1930), .ZN(n2135) );
  NAND2_X1 U1871 ( .A1(n1171), .A2(n1174), .ZN(n634) );
  NAND2_X1 U1872 ( .A1(n1159), .A2(n1161), .ZN(n627) );
  INV_X1 U1873 ( .A(n676), .ZN(n677) );
  NOR2_X1 U1874 ( .A1(n678), .A2(n677), .ZN(n334) );
  OR2_X1 U1875 ( .A1(n1194), .A2(n676), .ZN(n2136) );
  AND2_X1 U1876 ( .A1(n1194), .A2(n676), .ZN(n2137) );
  INV_X1 U1877 ( .A(n2270), .ZN(n2268) );
  INV_X1 U1878 ( .A(n1682), .ZN(n2309) );
  INV_X1 U1879 ( .A(n1507), .ZN(n2316) );
  INV_X1 U1880 ( .A(n682), .ZN(n683) );
  INV_X1 U1881 ( .A(n2144), .ZN(n2255) );
  AOI21_X1 U1882 ( .B1(n1933), .B2(n1932), .A(n1937), .ZN(n646) );
  NAND2_X1 U1883 ( .A1(n1181), .A2(n1192), .ZN(n645) );
  NOR2_X1 U1884 ( .A1(n1181), .A2(n1192), .ZN(n644) );
  NOR2_X1 U1885 ( .A1(n2139), .A2(n2140), .ZN(n2138) );
  NOR2_X1 U1886 ( .A1(n2193), .A2(n1683), .ZN(n2139) );
  NOR2_X1 U1887 ( .A1(n1682), .A2(n2252), .ZN(n2140) );
  INV_X1 U1888 ( .A(n724), .ZN(n725) );
  INV_X1 U1889 ( .A(n692), .ZN(n693) );
  INV_X1 U1890 ( .A(n1632), .ZN(n2311) );
  INV_X1 U1891 ( .A(n1532), .ZN(n2315) );
  INV_X1 U1892 ( .A(n1707), .ZN(n2308) );
  INV_X1 U1893 ( .A(n1607), .ZN(n2312) );
  INV_X1 U1894 ( .A(n1557), .ZN(n2314) );
  INV_X1 U1895 ( .A(n2173), .ZN(n2194) );
  INV_X1 U1896 ( .A(n802), .ZN(n803) );
  INV_X1 U1897 ( .A(n874), .ZN(n875) );
  INV_X1 U1898 ( .A(n1582), .ZN(n2313) );
  INV_X1 U1899 ( .A(n1732), .ZN(n2307) );
  INV_X1 U1900 ( .A(n1657), .ZN(n2310) );
  INV_X1 U1901 ( .A(n1482), .ZN(n2317) );
  XNOR2_X1 U1902 ( .A(n2303), .B(b[20]), .ZN(n1760) );
  XNOR2_X1 U1903 ( .A(n2300), .B(b[20]), .ZN(n1735) );
  XNOR2_X1 U1904 ( .A(n2269), .B(b[20]), .ZN(n1535) );
  XNOR2_X1 U1905 ( .A(n2273), .B(b[20]), .ZN(n1560) );
  XNOR2_X1 U1906 ( .A(n2276), .B(b[20]), .ZN(n1585) );
  XNOR2_X1 U1907 ( .A(n2264), .B(b[20]), .ZN(n1510) );
  XNOR2_X1 U1908 ( .A(n2284), .B(b[20]), .ZN(n1635) );
  XNOR2_X1 U1909 ( .A(n2297), .B(b[20]), .ZN(n1710) );
  XNOR2_X1 U1910 ( .A(n2281), .B(b[20]), .ZN(n1610) );
  XNOR2_X1 U1911 ( .A(n2294), .B(b[20]), .ZN(n1685) );
  XNOR2_X1 U1912 ( .A(n2289), .B(b[20]), .ZN(n1660) );
  XNOR2_X1 U1913 ( .A(n2299), .B(b[22]), .ZN(n1733) );
  XNOR2_X1 U1914 ( .A(n2303), .B(b[16]), .ZN(n1764) );
  XNOR2_X1 U1915 ( .A(n2299), .B(b[16]), .ZN(n1739) );
  XNOR2_X1 U1916 ( .A(n2264), .B(b[16]), .ZN(n1514) );
  XNOR2_X1 U1917 ( .A(n2273), .B(b[16]), .ZN(n1564) );
  XNOR2_X1 U1918 ( .A(n2269), .B(b[16]), .ZN(n1539) );
  XNOR2_X1 U1919 ( .A(n2275), .B(b[16]), .ZN(n1589) );
  XNOR2_X1 U1920 ( .A(n2281), .B(b[16]), .ZN(n1614) );
  XNOR2_X1 U1921 ( .A(n2171), .B(b[16]), .ZN(n1664) );
  XNOR2_X1 U1922 ( .A(n2285), .B(b[16]), .ZN(n1639) );
  XNOR2_X1 U1923 ( .A(n2294), .B(b[16]), .ZN(n1689) );
  XNOR2_X1 U1924 ( .A(n2302), .B(b[10]), .ZN(n1770) );
  XNOR2_X1 U1925 ( .A(n2280), .B(b[10]), .ZN(n1620) );
  XNOR2_X1 U1926 ( .A(n2285), .B(b[10]), .ZN(n1645) );
  XNOR2_X1 U1927 ( .A(n2170), .B(b[10]), .ZN(n1670) );
  XNOR2_X1 U1928 ( .A(n2276), .B(b[10]), .ZN(n1595) );
  XNOR2_X1 U1929 ( .A(n2268), .B(b[10]), .ZN(n1545) );
  XNOR2_X1 U1930 ( .A(n2293), .B(b[10]), .ZN(n1695) );
  XNOR2_X1 U1931 ( .A(n2300), .B(b[10]), .ZN(n1745) );
  XNOR2_X1 U1932 ( .A(n2297), .B(b[10]), .ZN(n1720) );
  XNOR2_X1 U1933 ( .A(n2304), .B(b[14]), .ZN(n1766) );
  XNOR2_X1 U1934 ( .A(n2303), .B(b[8]), .ZN(n1772) );
  XNOR2_X1 U1935 ( .A(n2304), .B(b[12]), .ZN(n1768) );
  XNOR2_X1 U1936 ( .A(b[23]), .B(n2300), .ZN(n1732) );
  XNOR2_X1 U1937 ( .A(n2276), .B(b[8]), .ZN(n1597) );
  XNOR2_X1 U1938 ( .A(n2284), .B(b[8]), .ZN(n1647) );
  XNOR2_X1 U1939 ( .A(n2296), .B(b[14]), .ZN(n1716) );
  XNOR2_X1 U1940 ( .A(n2293), .B(b[14]), .ZN(n1691) );
  XNOR2_X1 U1941 ( .A(n2280), .B(b[8]), .ZN(n1622) );
  XNOR2_X1 U1942 ( .A(n2268), .B(b[14]), .ZN(n1541) );
  XNOR2_X1 U1943 ( .A(n2268), .B(b[12]), .ZN(n1543) );
  XNOR2_X1 U1944 ( .A(n2284), .B(b[12]), .ZN(n1643) );
  XNOR2_X1 U1945 ( .A(n2271), .B(b[14]), .ZN(n1566) );
  XNOR2_X1 U1946 ( .A(n2285), .B(b[14]), .ZN(n1641) );
  XNOR2_X1 U1947 ( .A(n2280), .B(b[12]), .ZN(n1618) );
  XNOR2_X1 U1948 ( .A(n2293), .B(b[12]), .ZN(n1693) );
  XNOR2_X1 U1949 ( .A(n2276), .B(b[14]), .ZN(n1591) );
  XNOR2_X1 U1950 ( .A(n2296), .B(b[12]), .ZN(n1718) );
  XNOR2_X1 U1951 ( .A(n2300), .B(b[12]), .ZN(n1743) );
  XNOR2_X1 U1952 ( .A(n2293), .B(b[8]), .ZN(n1697) );
  XNOR2_X1 U1953 ( .A(n2273), .B(b[8]), .ZN(n1572) );
  XNOR2_X1 U1954 ( .A(n2280), .B(b[14]), .ZN(n1616) );
  XNOR2_X1 U1955 ( .A(n2268), .B(b[8]), .ZN(n1547) );
  XNOR2_X1 U1956 ( .A(n2275), .B(b[12]), .ZN(n1593) );
  XNOR2_X1 U1957 ( .A(n2300), .B(b[8]), .ZN(n1747) );
  XNOR2_X1 U1958 ( .A(n2303), .B(b[22]), .ZN(n1758) );
  XNOR2_X1 U1959 ( .A(n2302), .B(b[18]), .ZN(n1762) );
  XNOR2_X1 U1960 ( .A(n2302), .B(b[2]), .ZN(n1778) );
  XNOR2_X1 U1961 ( .A(n2304), .B(b[4]), .ZN(n1776) );
  XNOR2_X1 U1962 ( .A(n2268), .B(b[18]), .ZN(n1537) );
  XNOR2_X1 U1963 ( .A(n2300), .B(b[18]), .ZN(n1737) );
  XNOR2_X1 U1964 ( .A(n2275), .B(b[22]), .ZN(n1583) );
  XNOR2_X1 U1965 ( .A(n2264), .B(b[22]), .ZN(n1508) );
  XNOR2_X1 U1966 ( .A(n2273), .B(b[22]), .ZN(n1558) );
  XNOR2_X1 U1967 ( .A(n2275), .B(b[18]), .ZN(n1587) );
  XNOR2_X1 U1968 ( .A(n2269), .B(b[22]), .ZN(n1533) );
  XNOR2_X1 U1969 ( .A(n2268), .B(b[2]), .ZN(n1553) );
  XNOR2_X1 U1970 ( .A(n2281), .B(b[22]), .ZN(n1608) );
  XNOR2_X1 U1971 ( .A(n2268), .B(b[4]), .ZN(n1551) );
  XNOR2_X1 U1972 ( .A(n2275), .B(b[4]), .ZN(n1601) );
  XNOR2_X1 U1973 ( .A(n2275), .B(b[2]), .ZN(n1603) );
  XNOR2_X1 U1974 ( .A(n2293), .B(b[18]), .ZN(n1687) );
  XNOR2_X1 U1975 ( .A(n2285), .B(b[4]), .ZN(n1651) );
  XNOR2_X1 U1976 ( .A(n2280), .B(b[2]), .ZN(n1628) );
  XNOR2_X1 U1977 ( .A(n2284), .B(b[18]), .ZN(n1637) );
  XNOR2_X1 U1978 ( .A(n2293), .B(b[2]), .ZN(n1703) );
  XNOR2_X1 U1979 ( .A(n2170), .B(b[2]), .ZN(n1678) );
  XNOR2_X1 U1980 ( .A(n2280), .B(b[4]), .ZN(n1626) );
  XNOR2_X1 U1981 ( .A(n2293), .B(b[4]), .ZN(n1701) );
  XNOR2_X1 U1982 ( .A(n2280), .B(b[18]), .ZN(n1612) );
  XNOR2_X1 U1983 ( .A(n2300), .B(b[4]), .ZN(n1751) );
  XNOR2_X1 U1984 ( .A(n2296), .B(b[2]), .ZN(n1728) );
  XNOR2_X1 U1985 ( .A(n2304), .B(b[6]), .ZN(n1774) );
  XNOR2_X1 U1986 ( .A(n2276), .B(b[6]), .ZN(n1599) );
  XNOR2_X1 U1987 ( .A(n2268), .B(b[6]), .ZN(n1549) );
  XNOR2_X1 U1988 ( .A(n2280), .B(b[6]), .ZN(n1624) );
  XNOR2_X1 U1989 ( .A(n2293), .B(b[6]), .ZN(n1699) );
  XNOR2_X1 U1990 ( .A(n2300), .B(b[6]), .ZN(n1749) );
  XNOR2_X1 U1991 ( .A(b[23]), .B(n2288), .ZN(n1657) );
  XNOR2_X1 U1992 ( .A(b[23]), .B(n2271), .ZN(n1557) );
  XNOR2_X1 U1993 ( .A(b[1]), .B(n2259), .ZN(n1504) );
  XNOR2_X1 U1994 ( .A(b[1]), .B(n2285), .ZN(n1654) );
  XNOR2_X1 U1995 ( .A(b[3]), .B(n2259), .ZN(n1502) );
  XNOR2_X1 U1996 ( .A(b[3]), .B(n2284), .ZN(n1652) );
  XNOR2_X1 U1997 ( .A(b[3]), .B(n2171), .ZN(n1677) );
  XNOR2_X1 U1998 ( .A(b[3]), .B(n2299), .ZN(n1752) );
  XNOR2_X1 U1999 ( .A(b[1]), .B(n2299), .ZN(n1754) );
  XNOR2_X1 U2000 ( .A(b[1]), .B(n2293), .ZN(n1704) );
  XNOR2_X1 U2001 ( .A(b[9]), .B(n2284), .ZN(n1646) );
  XNOR2_X1 U2002 ( .A(b[9]), .B(n2259), .ZN(n1496) );
  XNOR2_X1 U2003 ( .A(b[7]), .B(n2259), .ZN(n1498) );
  XNOR2_X1 U2004 ( .A(b[7]), .B(n2288), .ZN(n1673) );
  XNOR2_X1 U2005 ( .A(b[7]), .B(n2285), .ZN(n1648) );
  XNOR2_X1 U2006 ( .A(b[9]), .B(n2271), .ZN(n1571) );
  XNOR2_X1 U2007 ( .A(b[5]), .B(n2259), .ZN(n1500) );
  XNOR2_X1 U2008 ( .A(b[5]), .B(n2299), .ZN(n1750) );
  XNOR2_X1 U2009 ( .A(b[21]), .B(n2259), .ZN(n1484) );
  XNOR2_X1 U2010 ( .A(b[11]), .B(n2259), .ZN(n1494) );
  XNOR2_X1 U2011 ( .A(b[15]), .B(n2259), .ZN(n1490) );
  XNOR2_X1 U2012 ( .A(b[13]), .B(n2259), .ZN(n1492) );
  XNOR2_X1 U2013 ( .A(b[19]), .B(n2259), .ZN(n1486) );
  XNOR2_X1 U2014 ( .A(b[17]), .B(n2259), .ZN(n1488) );
  NOR2_X1 U2015 ( .A1(n2146), .A2(n2149), .ZN(n2145) );
  AND2_X2 U2016 ( .A1(n2173), .A2(n1810), .ZN(n2147) );
  INV_X1 U2017 ( .A(a[13]), .ZN(n2282) );
  INV_X1 U2018 ( .A(a[23]), .ZN(n2261) );
  OAI21_X1 U2019 ( .B1(a[0]), .B2(n1982), .A(n2306), .ZN(n1458) );
  INV_X1 U2020 ( .A(n1757), .ZN(n2306) );
  XNOR2_X1 U2021 ( .A(b[23]), .B(n2259), .ZN(n1482) );
  XNOR2_X1 U2022 ( .A(n2039), .B(b[10]), .ZN(n1520) );
  XNOR2_X1 U2023 ( .A(n2039), .B(b[12]), .ZN(n1518) );
  XNOR2_X1 U2024 ( .A(n2264), .B(b[18]), .ZN(n1512) );
  XNOR2_X1 U2025 ( .A(n2039), .B(b[8]), .ZN(n1522) );
  XNOR2_X1 U2026 ( .A(n2039), .B(b[14]), .ZN(n1516) );
  XNOR2_X1 U2027 ( .A(n2263), .B(b[6]), .ZN(n1524) );
  XNOR2_X1 U2028 ( .A(n2263), .B(b[4]), .ZN(n1526) );
  XNOR2_X1 U2029 ( .A(n2263), .B(b[2]), .ZN(n1528) );
  INV_X1 U2030 ( .A(a[15]), .ZN(n2277) );
  OAI22_X1 U2031 ( .A1(n1969), .A2(n1584), .B1(n1960), .B2(n1583), .ZN(n1291)
         );
  OAI22_X1 U2032 ( .A1(n1968), .A2(n1590), .B1(n1961), .B2(n1589), .ZN(n1297)
         );
  OAI22_X1 U2033 ( .A1(n1968), .A2(n1588), .B1(n1961), .B2(n1587), .ZN(n1295)
         );
  OAI22_X1 U2034 ( .A1(n1968), .A2(n1586), .B1(n1960), .B2(n1585), .ZN(n1293)
         );
  OAI22_X1 U2035 ( .A1(n2227), .A2(n1592), .B1(n2244), .B2(n1591), .ZN(n1299)
         );
  CLKBUF_X1 U2036 ( .A(n2099), .Z(n2158) );
  CLKBUF_X1 U2037 ( .A(n1966), .Z(n2161) );
  CLKBUF_X1 U2038 ( .A(n2135), .Z(n2163) );
  OAI22_X1 U2039 ( .A1(n1992), .A2(n1772), .B1(n1771), .B2(n2258), .ZN(n1473)
         );
  OAI22_X1 U2040 ( .A1(n2235), .A2(n1780), .B1(n1779), .B2(n2258), .ZN(n1481)
         );
  OAI22_X1 U2041 ( .A1(n2235), .A2(n1777), .B1(n1776), .B2(n2258), .ZN(n1478)
         );
  OAI22_X1 U2042 ( .A1(n1992), .A2(n1776), .B1(n1775), .B2(n2258), .ZN(n1477)
         );
  OAI22_X1 U2043 ( .A1(n2235), .A2(n1779), .B1(n1778), .B2(n2258), .ZN(n1480)
         );
  OAI22_X1 U2044 ( .A1(n2235), .A2(n1775), .B1(n1774), .B2(n2258), .ZN(n1476)
         );
  OAI22_X1 U2045 ( .A1(n1992), .A2(n1773), .B1(n1772), .B2(n2258), .ZN(n1474)
         );
  OAI22_X1 U2046 ( .A1(n2235), .A2(n1778), .B1(n1777), .B2(n2258), .ZN(n1479)
         );
  OAI22_X1 U2047 ( .A1(n2235), .A2(n1774), .B1(n1773), .B2(n2258), .ZN(n1475)
         );
  OAI22_X1 U2048 ( .A1(n2235), .A2(n1769), .B1(n1768), .B2(n2258), .ZN(n1470)
         );
  OAI22_X1 U2049 ( .A1(n1992), .A2(n1771), .B1(n1770), .B2(n2258), .ZN(n1472)
         );
  XNOR2_X1 U2050 ( .A(b[9]), .B(n2292), .ZN(n1696) );
  XNOR2_X1 U2051 ( .A(b[3]), .B(n2292), .ZN(n1702) );
  XNOR2_X1 U2052 ( .A(b[7]), .B(n2292), .ZN(n1698) );
  XNOR2_X1 U2053 ( .A(b[5]), .B(n2292), .ZN(n1700) );
  INV_X1 U2054 ( .A(n508), .ZN(n2166) );
  AND2_X2 U2055 ( .A1(n1967), .A2(n1807), .ZN(n2167) );
  OR2_X1 U2056 ( .A1(n1021), .A2(n1038), .ZN(n2168) );
  XNOR2_X1 U2057 ( .A(n2272), .B(b[10]), .ZN(n1570) );
  XNOR2_X1 U2058 ( .A(b[3]), .B(n2272), .ZN(n1577) );
  XNOR2_X1 U2059 ( .A(n2283), .B(b[2]), .ZN(n1653) );
  XNOR2_X1 U2060 ( .A(n2283), .B(b[22]), .ZN(n1633) );
  XNOR2_X1 U2061 ( .A(b[23]), .B(n2283), .ZN(n1632) );
  XNOR2_X1 U2062 ( .A(n2283), .B(b[6]), .ZN(n1649) );
  XNOR2_X1 U2063 ( .A(b[5]), .B(n2285), .ZN(n1650) );
  INV_X1 U2064 ( .A(n2290), .ZN(n2171) );
  INV_X1 U2065 ( .A(n2290), .ZN(n2170) );
  INV_X1 U2066 ( .A(n2290), .ZN(n2288) );
  XNOR2_X1 U2067 ( .A(a[22]), .B(n2261), .ZN(n1806) );
  INV_X1 U2068 ( .A(n2149), .ZN(n2254) );
  XNOR2_X1 U2069 ( .A(n2299), .B(b[2]), .ZN(n1753) );
  XNOR2_X1 U2070 ( .A(b[7]), .B(n2300), .ZN(n1748) );
  XNOR2_X1 U2071 ( .A(b[9]), .B(n2300), .ZN(n1746) );
  XNOR2_X1 U2072 ( .A(n2300), .B(b[14]), .ZN(n1741) );
  INV_X2 U2073 ( .A(n2261), .ZN(n2260) );
  INV_X1 U2074 ( .A(a[19]), .ZN(n2270) );
  XOR2_X1 U2075 ( .A(a[14]), .B(n2282), .Z(n2173) );
  INV_X1 U2076 ( .A(n2169), .ZN(n2248) );
  INV_X1 U2077 ( .A(n2169), .ZN(n2247) );
  AOI21_X1 U2078 ( .B1(n2128), .B2(n1939), .A(n2124), .ZN(n600) );
  OAI22_X1 U2079 ( .A1(n1992), .A2(n1770), .B1(n1769), .B2(n2258), .ZN(n1471)
         );
  INV_X1 U2080 ( .A(a[0]), .ZN(n251) );
  NOR2_X1 U2081 ( .A1(n597), .A2(n599), .ZN(n595) );
  XNOR2_X1 U2082 ( .A(n2297), .B(b[4]), .ZN(n1726) );
  XNOR2_X1 U2083 ( .A(n2297), .B(b[8]), .ZN(n1722) );
  XNOR2_X1 U2084 ( .A(n2297), .B(b[6]), .ZN(n1724) );
  XNOR2_X1 U2085 ( .A(n2296), .B(b[22]), .ZN(n1708) );
  XNOR2_X1 U2086 ( .A(n2296), .B(b[18]), .ZN(n1712) );
  INV_X1 U2087 ( .A(a[21]), .ZN(n2175) );
  INV_X1 U2088 ( .A(a[21]), .ZN(n2265) );
  XNOR2_X1 U2089 ( .A(b[23]), .B(n2275), .ZN(n1582) );
  XNOR2_X1 U2090 ( .A(b[3]), .B(n2275), .ZN(n1602) );
  XNOR2_X1 U2091 ( .A(b[5]), .B(n2276), .ZN(n1600) );
  XNOR2_X1 U2092 ( .A(b[9]), .B(n2276), .ZN(n1596) );
  XNOR2_X1 U2093 ( .A(b[7]), .B(n2276), .ZN(n1598) );
  XNOR2_X1 U2094 ( .A(b[1]), .B(n2276), .ZN(n1604) );
  INV_X2 U2095 ( .A(n1931), .ZN(n2276) );
  INV_X1 U2096 ( .A(n2010), .ZN(n673) );
  OAI21_X1 U2097 ( .B1(n2147), .B2(n2194), .A(n2313), .ZN(n1290) );
  XNOR2_X1 U2098 ( .A(a[2]), .B(n1945), .ZN(n2176) );
  NAND2_X1 U2099 ( .A1(n1980), .A2(n896), .ZN(n2177) );
  NAND2_X1 U2100 ( .A1(n2009), .A2(n670), .ZN(n516) );
  NOR2_X1 U2101 ( .A1(n531), .A2(n534), .ZN(n525) );
  XNOR2_X1 U2102 ( .A(n2273), .B(b[18]), .ZN(n1562) );
  XNOR2_X1 U2103 ( .A(b[1]), .B(n2273), .ZN(n1579) );
  XNOR2_X1 U2104 ( .A(n2272), .B(b[2]), .ZN(n1578) );
  XNOR2_X1 U2105 ( .A(n2271), .B(b[12]), .ZN(n1568) );
  XNOR2_X1 U2106 ( .A(b[7]), .B(n2273), .ZN(n1573) );
  XNOR2_X1 U2107 ( .A(n2272), .B(b[6]), .ZN(n1574) );
  XNOR2_X1 U2108 ( .A(b[5]), .B(n2271), .ZN(n1575) );
  XNOR2_X1 U2109 ( .A(n2273), .B(b[4]), .ZN(n1576) );
  XNOR2_X1 U2110 ( .A(b[9]), .B(n2287), .ZN(n1671) );
  XNOR2_X1 U2111 ( .A(b[1]), .B(n2287), .ZN(n1679) );
  XNOR2_X1 U2112 ( .A(b[5]), .B(n2289), .ZN(n1675) );
  XNOR2_X1 U2113 ( .A(n2171), .B(b[8]), .ZN(n1672) );
  XNOR2_X1 U2114 ( .A(n2289), .B(b[4]), .ZN(n1676) );
  XNOR2_X1 U2115 ( .A(n2287), .B(b[6]), .ZN(n1674) );
  XNOR2_X1 U2116 ( .A(n2170), .B(b[22]), .ZN(n1658) );
  XNOR2_X1 U2117 ( .A(n2288), .B(b[18]), .ZN(n1662) );
  XNOR2_X1 U2118 ( .A(n2170), .B(b[14]), .ZN(n1666) );
  OAI21_X1 U2119 ( .B1(n2148), .B2(n2202), .A(n2314), .ZN(n1266) );
  AND2_X1 U2120 ( .A1(n821), .A2(n838), .ZN(n2178) );
  AND2_X1 U2121 ( .A1(n1806), .A2(n1930), .ZN(n2179) );
  NAND2_X1 U2122 ( .A1(n685), .A2(n688), .ZN(n369) );
  INV_X1 U2123 ( .A(n519), .ZN(n2180) );
  INV_X2 U2124 ( .A(n2174), .ZN(n2241) );
  NAND2_X1 U2125 ( .A1(n821), .A2(n838), .ZN(n503) );
  OAI21_X1 U2126 ( .B1(n2150), .B2(n1988), .A(n2310), .ZN(n1362) );
  NAND2_X1 U2127 ( .A1(n2213), .A2(n2177), .ZN(n320) );
  INV_X2 U2128 ( .A(n1983), .ZN(n2251) );
  NAND2_X1 U2129 ( .A1(n588), .A2(n2121), .ZN(n582) );
  XNOR2_X1 U2130 ( .A(n2047), .B(n2181), .ZN(n2206) );
  XNOR2_X1 U2131 ( .A(n898), .B(n881), .ZN(n2181) );
  OAI21_X1 U2132 ( .B1(n600), .B2(n597), .A(n598), .ZN(n596) );
  NOR2_X1 U2133 ( .A1(n2249), .A2(n2305), .ZN(n1385) );
  NOR2_X1 U2134 ( .A1(n2254), .A2(n2305), .ZN(n1433) );
  NOR2_X1 U2135 ( .A1(n2251), .A2(n2305), .ZN(n1409) );
  NOR2_X1 U2136 ( .A1(n2241), .A2(n2305), .ZN(n1265) );
  NOR2_X1 U2137 ( .A1(n2238), .A2(n2305), .ZN(n1241) );
  NAND2_X1 U2138 ( .A1(n2296), .A2(n2305), .ZN(n1731) );
  NOR2_X1 U2139 ( .A1(n2247), .A2(n2305), .ZN(n1361) );
  NAND2_X1 U2140 ( .A1(n2299), .A2(n2305), .ZN(n1756) );
  NOR2_X1 U2141 ( .A1(n1984), .A2(n2305), .ZN(n1289) );
  NOR2_X1 U2142 ( .A1(n1960), .A2(n2305), .ZN(n1313) );
  NOR2_X1 U2143 ( .A1(n2245), .A2(n2305), .ZN(n1337) );
  NOR2_X1 U2144 ( .A1(n2255), .A2(n2305), .ZN(n1457) );
  NAND2_X1 U2145 ( .A1(n2302), .A2(n2305), .ZN(n1781) );
  XNOR2_X1 U2146 ( .A(n2294), .B(b[0]), .ZN(n1705) );
  NAND2_X1 U2147 ( .A1(n2293), .A2(n2305), .ZN(n1706) );
  XNOR2_X1 U2148 ( .A(n2303), .B(b[0]), .ZN(n1780) );
  XNOR2_X1 U2149 ( .A(n2297), .B(b[0]), .ZN(n1730) );
  NAND2_X1 U2150 ( .A1(n2287), .A2(n2305), .ZN(n1681) );
  NAND2_X1 U2151 ( .A1(n2272), .A2(n2305), .ZN(n1581) );
  NAND2_X1 U2152 ( .A1(n2039), .A2(n2305), .ZN(n1531) );
  XNOR2_X1 U2153 ( .A(n2300), .B(b[0]), .ZN(n1755) );
  NAND2_X1 U2154 ( .A1(n2268), .A2(n2305), .ZN(n1556) );
  NAND2_X1 U2155 ( .A1(n2275), .A2(n2305), .ZN(n1606) );
  NAND2_X1 U2156 ( .A1(n2280), .A2(n2305), .ZN(n1631) );
  XNOR2_X1 U2157 ( .A(n2271), .B(b[0]), .ZN(n1580) );
  XNOR2_X1 U2158 ( .A(n2288), .B(b[0]), .ZN(n1680) );
  XNOR2_X1 U2159 ( .A(n2269), .B(b[0]), .ZN(n1555) );
  NAND2_X1 U2160 ( .A1(n2284), .A2(n2305), .ZN(n1656) );
  XNOR2_X1 U2161 ( .A(n2281), .B(b[0]), .ZN(n1630) );
  XNOR2_X1 U2162 ( .A(n2283), .B(b[0]), .ZN(n1655) );
  XNOR2_X1 U2163 ( .A(n2276), .B(b[0]), .ZN(n1605) );
  XNOR2_X1 U2164 ( .A(n2039), .B(b[0]), .ZN(n1530) );
  XNOR2_X1 U2165 ( .A(b[23]), .B(n2267), .ZN(n1532) );
  XNOR2_X1 U2166 ( .A(b[9]), .B(n2267), .ZN(n1546) );
  XNOR2_X1 U2167 ( .A(b[1]), .B(n2267), .ZN(n1554) );
  XNOR2_X1 U2168 ( .A(b[5]), .B(n2267), .ZN(n1550) );
  XNOR2_X1 U2169 ( .A(b[7]), .B(n2267), .ZN(n1548) );
  XNOR2_X1 U2170 ( .A(b[3]), .B(n2267), .ZN(n1552) );
  OAI22_X1 U2171 ( .A1(n2071), .A2(n1704), .B1(n2252), .B2(n1703), .ZN(n1407)
         );
  OAI22_X1 U2172 ( .A1(n2070), .A2(n1695), .B1(n1694), .B2(n2251), .ZN(n1398)
         );
  OAI22_X1 U2173 ( .A1(n2070), .A2(n1701), .B1(n1700), .B2(n2251), .ZN(n1404)
         );
  OAI22_X1 U2174 ( .A1(n2071), .A2(n1694), .B1(n2252), .B2(n1693), .ZN(n1397)
         );
  OAI22_X1 U2175 ( .A1(n2041), .A2(n1536), .B1(n2241), .B2(n1535), .ZN(n1245)
         );
  OAI22_X1 U2176 ( .A1(n2041), .A2(n1534), .B1(n2241), .B2(n1533), .ZN(n1243)
         );
  OAI22_X1 U2177 ( .A1(n2062), .A2(n1542), .B1(n2241), .B2(n1541), .ZN(n1251)
         );
  OAI22_X1 U2178 ( .A1(n2041), .A2(n1540), .B1(n2241), .B2(n1539), .ZN(n1249)
         );
  OAI22_X1 U2179 ( .A1(n2041), .A2(n1538), .B1(n2241), .B2(n1537), .ZN(n1247)
         );
  XNOR2_X1 U2180 ( .A(b[5]), .B(n2279), .ZN(n1625) );
  XNOR2_X1 U2181 ( .A(b[7]), .B(n2279), .ZN(n1623) );
  XNOR2_X1 U2182 ( .A(b[1]), .B(n2279), .ZN(n1629) );
  XNOR2_X1 U2183 ( .A(b[23]), .B(n2279), .ZN(n1607) );
  XNOR2_X1 U2184 ( .A(b[9]), .B(n2279), .ZN(n1621) );
  XNOR2_X1 U2185 ( .A(b[3]), .B(n2279), .ZN(n1627) );
  OAI21_X1 U2186 ( .B1(n2179), .B2(n2000), .A(n2317), .ZN(n1194) );
  XNOR2_X1 U2187 ( .A(n2260), .B(b[22]), .ZN(n1483) );
  XNOR2_X1 U2188 ( .A(n2260), .B(b[18]), .ZN(n1487) );
  XNOR2_X1 U2189 ( .A(n2260), .B(b[20]), .ZN(n1485) );
  XNOR2_X1 U2190 ( .A(n2260), .B(b[10]), .ZN(n1495) );
  XNOR2_X1 U2191 ( .A(n2260), .B(b[16]), .ZN(n1489) );
  XNOR2_X1 U2192 ( .A(n2260), .B(b[12]), .ZN(n1493) );
  XNOR2_X1 U2193 ( .A(n2260), .B(b[14]), .ZN(n1491) );
  XNOR2_X1 U2194 ( .A(n2260), .B(b[6]), .ZN(n1499) );
  NAND2_X1 U2195 ( .A1(n2260), .A2(n2305), .ZN(n1506) );
  XNOR2_X1 U2196 ( .A(n2260), .B(b[8]), .ZN(n1497) );
  XNOR2_X1 U2197 ( .A(n2260), .B(b[4]), .ZN(n1501) );
  XNOR2_X1 U2198 ( .A(n2260), .B(b[2]), .ZN(n1503) );
  XNOR2_X1 U2199 ( .A(n2260), .B(b[0]), .ZN(n1505) );
  XNOR2_X1 U2200 ( .A(b[3]), .B(n2296), .ZN(n1727) );
  XNOR2_X1 U2201 ( .A(b[1]), .B(n2296), .ZN(n1729) );
  XNOR2_X1 U2202 ( .A(b[5]), .B(n2297), .ZN(n1725) );
  XNOR2_X1 U2203 ( .A(b[9]), .B(n2296), .ZN(n1721) );
  XNOR2_X1 U2204 ( .A(b[23]), .B(n2297), .ZN(n1707) );
  XNOR2_X1 U2205 ( .A(b[7]), .B(n2297), .ZN(n1723) );
  NAND2_X1 U2206 ( .A1(n1210), .A2(n1276), .ZN(n2182) );
  NAND2_X1 U2207 ( .A1(n1210), .A2(n2138), .ZN(n2183) );
  NAND2_X1 U2208 ( .A1(n1276), .A2(n2138), .ZN(n2184) );
  NAND3_X1 U2209 ( .A1(n2182), .A2(n2183), .A3(n2184), .ZN(n834) );
  NAND2_X1 U2210 ( .A1(n1386), .A2(n830), .ZN(n2185) );
  NAND2_X1 U2211 ( .A1(n1386), .A2(n834), .ZN(n2186) );
  NAND2_X1 U2212 ( .A1(n830), .A2(n834), .ZN(n2187) );
  NAND3_X1 U2213 ( .A1(n2185), .A2(n2186), .A3(n2187), .ZN(n812) );
  OAI21_X1 U2214 ( .B1(n2230), .B2(n1983), .A(n2309), .ZN(n1386) );
  NOR2_X1 U2215 ( .A1(n805), .A2(n820), .ZN(n2188) );
  INV_X1 U2216 ( .A(n2006), .ZN(n2189) );
  INV_X1 U2217 ( .A(n2233), .ZN(n2190) );
  NOR2_X1 U2218 ( .A1(n805), .A2(n820), .ZN(n495) );
  NOR2_X1 U2219 ( .A1(n2188), .A2(n502), .ZN(n489) );
  INV_X2 U2220 ( .A(n1993), .ZN(n2283) );
  XNOR2_X1 U2221 ( .A(b[23]), .B(n2262), .ZN(n1507) );
  XNOR2_X1 U2222 ( .A(b[9]), .B(n2262), .ZN(n1521) );
  XNOR2_X1 U2223 ( .A(b[7]), .B(n2262), .ZN(n1523) );
  XNOR2_X1 U2224 ( .A(b[1]), .B(n2262), .ZN(n1529) );
  XNOR2_X1 U2225 ( .A(b[5]), .B(n2262), .ZN(n1525) );
  XNOR2_X1 U2226 ( .A(b[3]), .B(n2262), .ZN(n1527) );
  INV_X2 U2227 ( .A(n2175), .ZN(n2262) );
  BUF_X2 U2228 ( .A(n281), .Z(n2193) );
  INV_X1 U2229 ( .A(n281), .ZN(n2230) );
  XNOR2_X1 U2230 ( .A(n2294), .B(b[22]), .ZN(n1683) );
  XNOR2_X1 U2231 ( .A(b[23]), .B(n2292), .ZN(n1682) );
  INV_X1 U2232 ( .A(n2037), .ZN(n2278) );
  OAI21_X1 U2233 ( .B1(n2156), .B2(n1999), .A(n2312), .ZN(n1314) );
  XOR2_X1 U2234 ( .A(n933), .B(n952), .Z(n2195) );
  XOR2_X1 U2235 ( .A(n2195), .B(n937), .Z(n927) );
  NAND2_X1 U2236 ( .A1(n1259), .A2(n1347), .ZN(n2196) );
  NAND2_X1 U2237 ( .A1(n1259), .A2(n1303), .ZN(n2197) );
  NAND2_X1 U2238 ( .A1(n1347), .A2(n1303), .ZN(n2198) );
  NAND3_X1 U2239 ( .A1(n2196), .A2(n2197), .A3(n2198), .ZN(n936) );
  NAND2_X1 U2240 ( .A1(n933), .A2(n952), .ZN(n2199) );
  NAND2_X1 U2241 ( .A1(n933), .A2(n937), .ZN(n2200) );
  NAND2_X1 U2242 ( .A1(n952), .A2(n937), .ZN(n2201) );
  NAND3_X1 U2243 ( .A1(n2199), .A2(n2200), .A3(n2201), .ZN(n926) );
  NOR2_X1 U2244 ( .A1(n1003), .A2(n1020), .ZN(n569) );
  OAI21_X1 U2245 ( .B1(n620), .B2(n610), .A(n611), .ZN(n609) );
  OAI22_X1 U2246 ( .A1(n2071), .A2(n1702), .B1(n2251), .B2(n1701), .ZN(n1405)
         );
  NAND2_X1 U2247 ( .A1(n2168), .A2(n2120), .ZN(n571) );
  INV_X1 U2248 ( .A(n1962), .ZN(n2233) );
  INV_X2 U2249 ( .A(n1995), .ZN(n2271) );
  INV_X2 U2250 ( .A(n1994), .ZN(n2273) );
  OAI22_X1 U2251 ( .A1(n2193), .A2(n1696), .B1(n2252), .B2(n1695), .ZN(n1399)
         );
  OAI22_X1 U2252 ( .A1(n2193), .A2(n1698), .B1(n2251), .B2(n1697), .ZN(n1401)
         );
  OAI22_X1 U2253 ( .A1(n2193), .A2(n1700), .B1(n2252), .B2(n1699), .ZN(n1403)
         );
  OAI22_X1 U2254 ( .A1(n1699), .A2(n2193), .B1(n1698), .B2(n2251), .ZN(n1402)
         );
  AOI21_X1 U2255 ( .B1(n565), .B2(n552), .A(n2069), .ZN(n551) );
  INV_X1 U2256 ( .A(n2069), .ZN(n555) );
  OAI21_X1 U2257 ( .B1(n2040), .B2(n564), .A(n559), .ZN(n553) );
  NAND2_X1 U2258 ( .A1(n2118), .A2(n461), .ZN(n313) );
  INV_X1 U2259 ( .A(n461), .ZN(n459) );
  INV_X1 U2260 ( .A(n2233), .ZN(n2232) );
  INV_X1 U2261 ( .A(n2035), .ZN(n667) );
  OAI21_X1 U2262 ( .B1(n2152), .B2(n2169), .A(n2311), .ZN(n1338) );
  OAI21_X1 U2263 ( .B1(n2154), .B2(n1976), .A(n2315), .ZN(n1242) );
  INV_X1 U2264 ( .A(n2295), .ZN(n2291) );
  OAI21_X1 U2265 ( .B1(n2145), .B2(n2149), .A(n2308), .ZN(n1410) );
  NAND2_X1 U2266 ( .A1(n2192), .A2(n2118), .ZN(n456) );
  INV_X1 U2267 ( .A(n474), .ZN(n472) );
  INV_X1 U2268 ( .A(n547), .ZN(n674) );
  NOR2_X1 U2269 ( .A1(n554), .A2(n2066), .ZN(n545) );
  OAI21_X1 U2270 ( .B1(n555), .B2(n2066), .A(n550), .ZN(n546) );
  NAND2_X1 U2271 ( .A1(n941), .A2(n962), .ZN(n550) );
  OAI22_X1 U2272 ( .A1(n2235), .A2(n1764), .B1(n1763), .B2(n2258), .ZN(n1465)
         );
  OAI22_X1 U2273 ( .A1(n2234), .A2(n1759), .B1(n1758), .B2(n2257), .ZN(n1460)
         );
  OAI22_X1 U2274 ( .A1(n1992), .A2(n1768), .B1(n1767), .B2(n2258), .ZN(n1469)
         );
  OAI22_X1 U2275 ( .A1(n1992), .A2(n1767), .B1(n1766), .B2(n2258), .ZN(n1468)
         );
  OAI22_X1 U2276 ( .A1(n2235), .A2(n1760), .B1(n1759), .B2(n2258), .ZN(n1461)
         );
  OAI22_X1 U2277 ( .A1(n1992), .A2(n1763), .B1(n1762), .B2(n2258), .ZN(n1464)
         );
  OAI22_X1 U2278 ( .A1(n2234), .A2(n1761), .B1(n1760), .B2(n2257), .ZN(n1462)
         );
  OAI22_X1 U2279 ( .A1(n2234), .A2(n1758), .B1(n1757), .B2(n2257), .ZN(n1459)
         );
  OAI22_X1 U2280 ( .A1(n1992), .A2(n1765), .B1(n1764), .B2(n2258), .ZN(n1466)
         );
  XNOR2_X1 U2281 ( .A(b[1]), .B(n2302), .ZN(n1779) );
  OAI22_X1 U2282 ( .A1(n1992), .A2(n1766), .B1(n1765), .B2(n2258), .ZN(n1467)
         );
  XNOR2_X1 U2283 ( .A(b[5]), .B(n2304), .ZN(n1775) );
  XNOR2_X1 U2284 ( .A(b[7]), .B(n2302), .ZN(n1773) );
  OAI22_X1 U2285 ( .A1(n2234), .A2(n1762), .B1(n1761), .B2(n2257), .ZN(n1463)
         );
  XNOR2_X1 U2286 ( .A(b[3]), .B(n2303), .ZN(n1777) );
  XNOR2_X1 U2287 ( .A(b[9]), .B(n2302), .ZN(n1771) );
  XNOR2_X1 U2288 ( .A(b[23]), .B(n2303), .ZN(n1757) );
  INV_X1 U2289 ( .A(n2091), .ZN(n508) );
  INV_X1 U2290 ( .A(n520), .ZN(n670) );
  AOI21_X1 U2291 ( .B1(n526), .B2(n511), .A(n512), .ZN(n506) );
  NAND2_X1 U2292 ( .A1(n839), .A2(n856), .ZN(n514) );
  AOI21_X1 U2293 ( .B1(n595), .B2(n609), .A(n596), .ZN(n594) );
  AOI21_X1 U2294 ( .B1(n589), .B2(n2121), .A(n1941), .ZN(n583) );
  OAI21_X1 U2295 ( .B1(n2167), .B2(n1954), .A(n2316), .ZN(n1218) );
  INV_X1 U2296 ( .A(n2203), .ZN(n2238) );
  AOI21_X1 U2297 ( .B1(n2118), .B2(n472), .A(n459), .ZN(n457) );
  NOR2_X1 U2298 ( .A1(n838), .A2(n821), .ZN(n502) );
  NAND2_X1 U2299 ( .A1(n668), .A2(n503), .ZN(n317) );
  AOI21_X1 U2300 ( .B1(n2168), .B2(n2119), .A(n1942), .ZN(n572) );
  OAI22_X1 U2301 ( .A1(n2062), .A2(n1535), .B1(n1534), .B2(n2241), .ZN(n1244)
         );
  OAI22_X1 U2302 ( .A1(n2041), .A2(n1537), .B1(n1536), .B2(n2241), .ZN(n1246)
         );
  OAI22_X1 U2303 ( .A1(n2041), .A2(n1541), .B1(n1540), .B2(n2241), .ZN(n1250)
         );
  OAI22_X1 U2304 ( .A1(n2041), .A2(n1539), .B1(n1538), .B2(n2241), .ZN(n1248)
         );
  OAI22_X1 U2305 ( .A1(n2062), .A2(n1533), .B1(n1532), .B2(n2241), .ZN(n692)
         );
  OAI22_X1 U2306 ( .A1(n2062), .A2(n1543), .B1(n1542), .B2(n2241), .ZN(n1252)
         );
  OAI22_X1 U2307 ( .A1(n1556), .A2(n2241), .B1(n2041), .B2(n2172), .ZN(n1184)
         );
  NAND2_X1 U2308 ( .A1(n2127), .A2(n378), .ZN(n305) );
  NAND2_X1 U2309 ( .A1(n382), .A2(n2127), .ZN(n371) );
  AOI21_X1 U2310 ( .B1(n383), .B2(n2127), .A(n376), .ZN(n372) );
  INV_X1 U2311 ( .A(n490), .ZN(n492) );
  NOR2_X1 U2312 ( .A1(n983), .A2(n1002), .ZN(n563) );
  NAND2_X1 U2313 ( .A1(n1416), .A2(n1306), .ZN(n2207) );
  NAND2_X1 U2314 ( .A1(n1416), .A2(n1328), .ZN(n2208) );
  NAND2_X1 U2315 ( .A1(n1306), .A2(n1328), .ZN(n2209) );
  NAND3_X1 U2316 ( .A1(n2207), .A2(n2208), .A3(n2209), .ZN(n994) );
  CLKBUF_X1 U2317 ( .A(n535), .Z(n2210) );
  OR2_X1 U2318 ( .A1(n2108), .A2(n1714), .ZN(n2211) );
  OR2_X1 U2319 ( .A1(n1713), .A2(n2254), .ZN(n2212) );
  NAND2_X1 U2320 ( .A1(n2211), .A2(n2212), .ZN(n1416) );
  XNOR2_X1 U2321 ( .A(n2296), .B(b[16]), .ZN(n1714) );
  NAND2_X1 U2322 ( .A1(n877), .A2(n896), .ZN(n532) );
  AOI21_X1 U2323 ( .B1(n629), .B2(n635), .A(n630), .ZN(n628) );
  OAI21_X1 U2324 ( .B1(n628), .B2(n626), .A(n627), .ZN(n625) );
  AOI21_X1 U2325 ( .B1(n625), .B2(n1943), .A(n1935), .ZN(n620) );
  NAND2_X1 U2326 ( .A1(n670), .A2(n2180), .ZN(n319) );
  INV_X1 U2327 ( .A(n521), .ZN(n519) );
  NOR2_X1 U2328 ( .A1(n857), .A2(n876), .ZN(n520) );
  NAND2_X1 U2329 ( .A1(n857), .A2(n876), .ZN(n521) );
  XNOR2_X1 U2330 ( .A(n497), .B(n316), .ZN(product[30]) );
  NAND2_X1 U2331 ( .A1(n1085), .A2(n1098), .ZN(n593) );
  NAND2_X1 U2332 ( .A1(n897), .A2(n918), .ZN(n535) );
  XNOR2_X1 U2333 ( .A(b[19]), .B(n2266), .ZN(n1536) );
  XNOR2_X1 U2334 ( .A(b[21]), .B(n2266), .ZN(n1534) );
  XNOR2_X1 U2335 ( .A(b[17]), .B(n2266), .ZN(n1538) );
  XNOR2_X1 U2336 ( .A(b[13]), .B(n2266), .ZN(n1542) );
  XNOR2_X1 U2337 ( .A(b[15]), .B(n2266), .ZN(n1540) );
  XNOR2_X1 U2338 ( .A(b[11]), .B(n2266), .ZN(n1544) );
  NAND2_X1 U2339 ( .A1(n2128), .A2(n2129), .ZN(n599) );
  OR2_X1 U2340 ( .A1(n1980), .A2(n896), .ZN(n2213) );
  OAI22_X1 U2341 ( .A1(n2054), .A2(n1733), .B1(n1732), .B2(n2255), .ZN(n2214)
         );
  NOR2_X1 U2342 ( .A1(n336), .A2(n334), .ZN(n332) );
  NAND2_X1 U2343 ( .A1(n709), .A2(n716), .ZN(n409) );
  INV_X1 U2344 ( .A(n400), .ZN(n398) );
  NAND2_X1 U2345 ( .A1(n400), .A2(n2125), .ZN(n389) );
  NAND2_X1 U2346 ( .A1(n727), .A2(n736), .ZN(n429) );
  INV_X1 U2347 ( .A(n2286), .ZN(n2284) );
  INV_X1 U2348 ( .A(n537), .ZN(n536) );
  OAI21_X1 U2349 ( .B1(n590), .B2(n593), .A(n591), .ZN(n589) );
  NAND2_X1 U2350 ( .A1(n1071), .A2(n1084), .ZN(n591) );
  NOR2_X1 U2351 ( .A1(n1071), .A2(n1084), .ZN(n590) );
  NOR2_X1 U2352 ( .A1(n571), .A2(n569), .ZN(n567) );
  NAND2_X1 U2353 ( .A1(n996), .A2(n994), .ZN(n2215) );
  NAND2_X1 U2354 ( .A1(n996), .A2(n1217), .ZN(n2216) );
  NAND2_X1 U2355 ( .A1(n994), .A2(n1217), .ZN(n2217) );
  NAND3_X1 U2356 ( .A1(n2215), .A2(n2216), .A3(n2217), .ZN(n972) );
  OR2_X1 U2357 ( .A1(n1964), .A2(n1668), .ZN(n2218) );
  OR2_X1 U2358 ( .A1(n1667), .A2(n2249), .ZN(n2219) );
  NAND2_X1 U2359 ( .A1(n2218), .A2(n2219), .ZN(n1372) );
  NOR2_X1 U2360 ( .A1(n2236), .A2(n2305), .ZN(n1217) );
  XNOR2_X1 U2361 ( .A(n2289), .B(b[12]), .ZN(n1668) );
  OAI22_X1 U2362 ( .A1(n2070), .A2(n1705), .B1(n1704), .B2(n2252), .ZN(n1408)
         );
  NOR2_X1 U2363 ( .A1(n513), .A2(n520), .ZN(n511) );
  OAI21_X1 U2364 ( .B1(n513), .B2(n521), .A(n514), .ZN(n512) );
  INV_X1 U2365 ( .A(n2096), .ZN(n565) );
  NOR2_X1 U2366 ( .A1(n633), .A2(n631), .ZN(n629) );
  NAND2_X1 U2367 ( .A1(n507), .A2(n2189), .ZN(n487) );
  INV_X1 U2368 ( .A(n502), .ZN(n668) );
  OAI21_X1 U2369 ( .B1(n2029), .B2(n1986), .A(n2307), .ZN(n1434) );
  NOR2_X1 U2370 ( .A1(n2061), .A2(n547), .ZN(n540) );
  OAI22_X1 U2371 ( .A1(n2193), .A2(n1697), .B1(n1696), .B2(n2251), .ZN(n1400)
         );
  NAND2_X1 U2372 ( .A1(n2016), .A2(n2210), .ZN(n321) );
  OAI21_X1 U2373 ( .B1(n550), .B2(n542), .A(n543), .ZN(n541) );
  INV_X1 U2374 ( .A(n346), .ZN(n344) );
  OAI21_X1 U2375 ( .B1(n337), .B2(n334), .A(n335), .ZN(n333) );
  NAND2_X1 U2376 ( .A1(n717), .A2(n726), .ZN(n418) );
  OAI22_X1 U2377 ( .A1(n2193), .A2(n1703), .B1(n1702), .B2(n2251), .ZN(n1406)
         );
  INV_X1 U2378 ( .A(n2051), .ZN(n2302) );
  NAND2_X1 U2379 ( .A1(n789), .A2(n804), .ZN(n481) );
  NOR2_X1 U2380 ( .A1(n456), .A2(n480), .ZN(n454) );
  OAI21_X1 U2381 ( .B1(n492), .B2(n480), .A(n481), .ZN(n479) );
  NOR2_X1 U2382 ( .A1(n2006), .A2(n480), .ZN(n478) );
  OAI21_X1 U2383 ( .B1(n572), .B2(n1948), .A(n570), .ZN(n568) );
  OAI21_X1 U2384 ( .B1(n594), .B2(n582), .A(n583), .ZN(n581) );
  OAI21_X1 U2385 ( .B1(n456), .B2(n481), .A(n457), .ZN(n455) );
  INV_X1 U2386 ( .A(n2179), .ZN(n2223) );
  NAND2_X1 U2387 ( .A1(n919), .A2(n940), .ZN(n543) );
  OAI21_X1 U2388 ( .B1(n495), .B2(n503), .A(n496), .ZN(n490) );
  INV_X1 U2389 ( .A(n420), .ZN(n422) );
  NOR2_X1 U2390 ( .A1(n420), .A2(n347), .ZN(n345) );
  AOI21_X2 U2391 ( .B1(n426), .B2(n445), .A(n427), .ZN(n421) );
  NAND2_X1 U2392 ( .A1(n426), .A2(n663), .ZN(n420) );
  NAND2_X1 U2393 ( .A1(n737), .A2(n748), .ZN(n436) );
  NOR2_X1 U2394 ( .A1(n737), .A2(n748), .ZN(n435) );
  AOI21_X1 U2395 ( .B1(n508), .B2(n478), .A(n479), .ZN(n477) );
  AOI21_X1 U2396 ( .B1(n508), .B2(n465), .A(n466), .ZN(n464) );
  AOI21_X1 U2397 ( .B1(n508), .B2(n668), .A(n2178), .ZN(n499) );
  AOI21_X1 U2398 ( .B1(n508), .B2(n2189), .A(n1978), .ZN(n488) );
  NAND2_X1 U2399 ( .A1(n537), .A2(n450), .ZN(n2220) );
  INV_X1 U2400 ( .A(n451), .ZN(n2221) );
  OAI22_X1 U2401 ( .A1(n2229), .A2(n1683), .B1(n1682), .B2(n2251), .ZN(n2222)
         );
  INV_X1 U2402 ( .A(n401), .ZN(n399) );
  OAI21_X1 U2403 ( .B1(n390), .B2(n384), .A(n387), .ZN(n383) );
  AOI21_X1 U2404 ( .B1(n401), .B2(n2125), .A(n394), .ZN(n390) );
  NOR2_X1 U2405 ( .A1(n749), .A2(n760), .ZN(n438) );
  NAND2_X1 U2406 ( .A1(n749), .A2(n760), .ZN(n439) );
  INV_X1 U2407 ( .A(n2052), .ZN(n2303) );
  INV_X1 U2408 ( .A(n345), .ZN(n343) );
  NAND2_X1 U2409 ( .A1(n345), .A2(n2134), .ZN(n336) );
  NAND2_X1 U2410 ( .A1(n694), .A2(n689), .ZN(n378) );
  INV_X1 U2411 ( .A(n706), .ZN(n707) );
  XNOR2_X1 U2412 ( .A(n475), .B(n314), .ZN(product[32]) );
  XNOR2_X1 U2413 ( .A(n462), .B(n313), .ZN(product[33]) );
  NAND2_X1 U2414 ( .A1(n805), .A2(n820), .ZN(n496) );
  OAI22_X1 U2415 ( .A1(n1781), .A2(n2258), .B1(n1992), .B2(n2051), .ZN(n1193)
         );
  OAI22_X1 U2416 ( .A1(n1968), .A2(n1593), .B1(n1592), .B2(n1961), .ZN(n1300)
         );
  OAI22_X1 U2417 ( .A1(n1969), .A2(n1589), .B1(n1588), .B2(n2243), .ZN(n1296)
         );
  OAI22_X1 U2418 ( .A1(n2227), .A2(n1583), .B1(n1582), .B2(n1961), .ZN(n724)
         );
  OAI22_X1 U2419 ( .A1(n1968), .A2(n1591), .B1(n1590), .B2(n1961), .ZN(n1298)
         );
  OAI22_X1 U2420 ( .A1(n1969), .A2(n1587), .B1(n1586), .B2(n1961), .ZN(n1294)
         );
  OAI22_X1 U2421 ( .A1(n2227), .A2(n1585), .B1(n1584), .B2(n2243), .ZN(n1292)
         );
  OAI22_X1 U2422 ( .A1(n1606), .A2(n2243), .B1(n2228), .B2(n1996), .ZN(n1186)
         );
  NAND2_X1 U2423 ( .A1(n761), .A2(n774), .ZN(n461) );
  NAND2_X1 U2424 ( .A1(n663), .A2(n662), .ZN(n431) );
  INV_X1 U2425 ( .A(n772), .ZN(n773) );
  XNOR2_X1 U2426 ( .A(b[11]), .B(n2289), .ZN(n1669) );
  XNOR2_X1 U2427 ( .A(b[17]), .B(n2287), .ZN(n1663) );
  XNOR2_X1 U2428 ( .A(b[19]), .B(n2171), .ZN(n1661) );
  XNOR2_X1 U2429 ( .A(b[13]), .B(n2171), .ZN(n1667) );
  XNOR2_X1 U2430 ( .A(b[15]), .B(n2288), .ZN(n1665) );
  XNOR2_X1 U2431 ( .A(b[21]), .B(n2170), .ZN(n1659) );
  XNOR2_X1 U2432 ( .A(n437), .B(n311), .ZN(product[35]) );
  OAI22_X1 U2433 ( .A1(n1979), .A2(n1570), .B1(n1569), .B2(n1984), .ZN(n1278)
         );
  OAI22_X1 U2434 ( .A1(n1990), .A2(n1575), .B1(n2242), .B2(n1574), .ZN(n1283)
         );
  OAI22_X1 U2435 ( .A1(n1979), .A2(n1573), .B1(n1984), .B2(n1572), .ZN(n1281)
         );
  OAI22_X1 U2436 ( .A1(n2225), .A2(n1571), .B1(n2038), .B2(n1570), .ZN(n1279)
         );
  OAI22_X1 U2437 ( .A1(n2225), .A2(n1580), .B1(n1579), .B2(n2038), .ZN(n1288)
         );
  OAI22_X1 U2438 ( .A1(n1979), .A2(n1579), .B1(n2242), .B2(n1578), .ZN(n1287)
         );
  OAI22_X1 U2439 ( .A1(n2225), .A2(n1578), .B1(n1577), .B2(n2038), .ZN(n1286)
         );
  OAI22_X1 U2440 ( .A1(n2226), .A2(n1569), .B1(n2038), .B2(n1568), .ZN(n1277)
         );
  OAI22_X1 U2441 ( .A1(n2226), .A2(n1577), .B1(n2242), .B2(n1576), .ZN(n1285)
         );
  OAI22_X1 U2442 ( .A1(n1991), .A2(n1572), .B1(n1571), .B2(n2242), .ZN(n1280)
         );
  OAI22_X1 U2443 ( .A1(n2225), .A2(n1576), .B1(n1575), .B2(n2242), .ZN(n1284)
         );
  OAI22_X1 U2444 ( .A1(n1990), .A2(n1574), .B1(n1573), .B2(n2242), .ZN(n1282)
         );
  XNOR2_X1 U2445 ( .A(n430), .B(n310), .ZN(product[36]) );
  OAI22_X1 U2446 ( .A1(n2059), .A2(n1613), .B1(n2246), .B2(n1612), .ZN(n1319)
         );
  OAI22_X1 U2447 ( .A1(n2059), .A2(n1612), .B1(n1611), .B2(n2246), .ZN(n1318)
         );
  OAI22_X1 U2448 ( .A1(n2059), .A2(n1609), .B1(n2246), .B2(n1608), .ZN(n1315)
         );
  OAI22_X1 U2449 ( .A1(n2059), .A2(n1610), .B1(n1609), .B2(n2245), .ZN(n1316)
         );
  OAI22_X1 U2450 ( .A1(n2058), .A2(n1611), .B1(n2245), .B2(n1610), .ZN(n1317)
         );
  OAI22_X1 U2451 ( .A1(n1631), .A2(n2245), .B1(n2059), .B2(n2037), .ZN(n1187)
         );
  OAI22_X1 U2452 ( .A1(n2059), .A2(n1617), .B1(n2245), .B2(n1616), .ZN(n1323)
         );
  OAI22_X1 U2453 ( .A1(n2059), .A2(n1615), .B1(n2246), .B2(n1614), .ZN(n1321)
         );
  OAI22_X1 U2454 ( .A1(n2107), .A2(n1618), .B1(n1617), .B2(n2246), .ZN(n1324)
         );
  OAI22_X1 U2455 ( .A1(n2107), .A2(n1614), .B1(n1613), .B2(n2245), .ZN(n1320)
         );
  OAI22_X1 U2456 ( .A1(n2058), .A2(n1616), .B1(n1615), .B2(n2246), .ZN(n1322)
         );
  XNOR2_X1 U2457 ( .A(n419), .B(n309), .ZN(product[37]) );
  OAI22_X1 U2458 ( .A1(n2163), .A2(n1483), .B1(n1482), .B2(n2236), .ZN(n676)
         );
  OAI22_X1 U2459 ( .A1(n2165), .A2(n1484), .B1(n1985), .B2(n1483), .ZN(n1195)
         );
  OAI22_X1 U2460 ( .A1(n2165), .A2(n1485), .B1(n1484), .B2(n2236), .ZN(n1196)
         );
  OAI22_X1 U2461 ( .A1(n2165), .A2(n1491), .B1(n1490), .B2(n1985), .ZN(n1202)
         );
  OAI22_X1 U2462 ( .A1(n2165), .A2(n1486), .B1(n2236), .B2(n1485), .ZN(n1197)
         );
  OAI22_X1 U2463 ( .A1(n2163), .A2(n1488), .B1(n1985), .B2(n1487), .ZN(n1199)
         );
  OAI22_X1 U2464 ( .A1(n2165), .A2(n1490), .B1(n1985), .B2(n1489), .ZN(n1201)
         );
  OAI22_X1 U2465 ( .A1(n2163), .A2(n1487), .B1(n1486), .B2(n2236), .ZN(n1198)
         );
  OAI22_X1 U2466 ( .A1(n2163), .A2(n1492), .B1(n1985), .B2(n1491), .ZN(n1203)
         );
  OAI22_X1 U2467 ( .A1(n2163), .A2(n1493), .B1(n1492), .B2(n2237), .ZN(n1204)
         );
  OAI22_X1 U2468 ( .A1(n2165), .A2(n1489), .B1(n1488), .B2(n2236), .ZN(n1200)
         );
  OAI22_X1 U2469 ( .A1(n1506), .A2(n2237), .B1(n2164), .B2(n2261), .ZN(n1182)
         );
  INV_X1 U2470 ( .A(n428), .ZN(n661) );
  INV_X1 U2471 ( .A(n421), .ZN(n423) );
  OAI21_X1 U2472 ( .B1(n428), .B2(n436), .A(n429), .ZN(n427) );
  OAI22_X1 U2473 ( .A1(n2005), .A2(n1508), .B1(n1507), .B2(n2056), .ZN(n682)
         );
  OAI22_X1 U2474 ( .A1(n1955), .A2(n1513), .B1(n2239), .B2(n1512), .ZN(n1223)
         );
  OAI22_X1 U2475 ( .A1(n1981), .A2(n1518), .B1(n1517), .B2(n2056), .ZN(n1228)
         );
  OAI22_X1 U2476 ( .A1(n2005), .A2(n1509), .B1(n2239), .B2(n1508), .ZN(n1219)
         );
  OAI22_X1 U2477 ( .A1(n1956), .A2(n1514), .B1(n1513), .B2(n2056), .ZN(n1224)
         );
  OAI22_X1 U2478 ( .A1(n1956), .A2(n1511), .B1(n2238), .B2(n1510), .ZN(n1221)
         );
  OAI22_X1 U2479 ( .A1(n2005), .A2(n1515), .B1(n2239), .B2(n1514), .ZN(n1225)
         );
  OAI22_X1 U2480 ( .A1(n1955), .A2(n1510), .B1(n1509), .B2(n2056), .ZN(n1220)
         );
  OAI22_X1 U2481 ( .A1(n1531), .A2(n2056), .B1(n1955), .B2(n2265), .ZN(n1183)
         );
  OAI22_X1 U2482 ( .A1(n2004), .A2(n1517), .B1(n2239), .B2(n1516), .ZN(n1227)
         );
  OAI22_X1 U2483 ( .A1(n1981), .A2(n1512), .B1(n1511), .B2(n2056), .ZN(n1222)
         );
  OAI22_X1 U2484 ( .A1(n1955), .A2(n1516), .B1(n1515), .B2(n2056), .ZN(n1226)
         );
  OAI22_X1 U2485 ( .A1(n2160), .A2(n1652), .B1(n2247), .B2(n1651), .ZN(n1357)
         );
  OAI22_X1 U2486 ( .A1(n1950), .A2(n1649), .B1(n1648), .B2(n2248), .ZN(n1354)
         );
  OAI22_X1 U2487 ( .A1(n1949), .A2(n1645), .B1(n1644), .B2(n2248), .ZN(n1350)
         );
  OAI22_X1 U2488 ( .A1(n2158), .A2(n1647), .B1(n1646), .B2(n2247), .ZN(n1352)
         );
  OAI22_X1 U2489 ( .A1(n2160), .A2(n1653), .B1(n1652), .B2(n2247), .ZN(n1358)
         );
  OAI22_X1 U2490 ( .A1(n1950), .A2(n1648), .B1(n2247), .B2(n1647), .ZN(n1353)
         );
  OAI22_X1 U2491 ( .A1(n2099), .A2(n1644), .B1(n2248), .B2(n1643), .ZN(n1349)
         );
  OAI22_X1 U2492 ( .A1(n1949), .A2(n1654), .B1(n2248), .B2(n1653), .ZN(n1359)
         );
  OAI22_X1 U2493 ( .A1(n2160), .A2(n1650), .B1(n2247), .B2(n1649), .ZN(n1355)
         );
  OAI22_X1 U2494 ( .A1(n2158), .A2(n1655), .B1(n1654), .B2(n2247), .ZN(n1360)
         );
  OAI22_X1 U2495 ( .A1(n2099), .A2(n1646), .B1(n2247), .B2(n1645), .ZN(n1351)
         );
  OAI22_X1 U2496 ( .A1(n2099), .A2(n1651), .B1(n1650), .B2(n2247), .ZN(n1356)
         );
  OAI22_X1 U2497 ( .A1(n2108), .A2(n1718), .B1(n1717), .B2(n2254), .ZN(n1420)
         );
  OAI22_X1 U2498 ( .A1(n1731), .A2(n2254), .B1(n2231), .B2(n2298), .ZN(n1191)
         );
  OAI22_X1 U2499 ( .A1(n2108), .A2(n1716), .B1(n1715), .B2(n2253), .ZN(n1418)
         );
  OAI22_X1 U2500 ( .A1(n2108), .A2(n1715), .B1(n2253), .B2(n1714), .ZN(n1417)
         );
  OAI22_X1 U2501 ( .A1(n2108), .A2(n1713), .B1(n2254), .B2(n1712), .ZN(n1415)
         );
  OAI22_X1 U2502 ( .A1(n2108), .A2(n1717), .B1(n2254), .B2(n1716), .ZN(n1419)
         );
  OAI22_X1 U2503 ( .A1(n2108), .A2(n1708), .B1(n1707), .B2(n2254), .ZN(n874)
         );
  OAI22_X1 U2504 ( .A1(n2108), .A2(n1711), .B1(n2253), .B2(n1710), .ZN(n1413)
         );
  OAI22_X1 U2505 ( .A1(n2108), .A2(n1709), .B1(n2253), .B2(n1708), .ZN(n1411)
         );
  OAI22_X1 U2506 ( .A1(n2108), .A2(n1710), .B1(n1709), .B2(n2254), .ZN(n1412)
         );
  OAI22_X1 U2507 ( .A1(n2108), .A2(n1712), .B1(n1711), .B2(n2253), .ZN(n1414)
         );
  XNOR2_X1 U2508 ( .A(n410), .B(n308), .ZN(product[38]) );
  NAND2_X1 U2509 ( .A1(n775), .A2(n788), .ZN(n474) );
  XNOR2_X1 U2510 ( .A(b[17]), .B(n2304), .ZN(n1763) );
  XNOR2_X1 U2511 ( .A(b[21]), .B(n2302), .ZN(n1759) );
  XNOR2_X1 U2512 ( .A(b[13]), .B(n2303), .ZN(n1767) );
  XNOR2_X1 U2513 ( .A(b[19]), .B(n2304), .ZN(n1761) );
  XNOR2_X1 U2514 ( .A(b[15]), .B(n2302), .ZN(n1765) );
  XNOR2_X1 U2515 ( .A(b[11]), .B(n2304), .ZN(n1769) );
  NAND2_X1 U2516 ( .A1(n332), .A2(n2136), .ZN(n326) );
  AOI21_X1 U2517 ( .B1(n333), .B2(n2136), .A(n2137), .ZN(n327) );
  NAND2_X1 U2518 ( .A1(n1165), .A2(n1170), .ZN(n632) );
  OAI22_X1 U2519 ( .A1(n2191), .A2(n1753), .B1(n1752), .B2(n2256), .ZN(n1454)
         );
  OAI22_X1 U2520 ( .A1(n2191), .A2(n1747), .B1(n1746), .B2(n2255), .ZN(n1448)
         );
  OAI22_X1 U2521 ( .A1(n2191), .A2(n1750), .B1(n2255), .B2(n1749), .ZN(n1451)
         );
  OAI22_X1 U2522 ( .A1(n2191), .A2(n1749), .B1(n1748), .B2(n2256), .ZN(n1450)
         );
  OAI22_X1 U2523 ( .A1(n2191), .A2(n1745), .B1(n1744), .B2(n2256), .ZN(n1446)
         );
  OAI22_X1 U2524 ( .A1(n2191), .A2(n1748), .B1(n2255), .B2(n1747), .ZN(n1449)
         );
  OAI22_X1 U2525 ( .A1(n2190), .A2(n1744), .B1(n2255), .B2(n1743), .ZN(n1445)
         );
  OAI22_X1 U2526 ( .A1(n2190), .A2(n1746), .B1(n2255), .B2(n1745), .ZN(n1447)
         );
  OAI22_X1 U2527 ( .A1(n2191), .A2(n1754), .B1(n2256), .B2(n1753), .ZN(n1455)
         );
  OAI22_X1 U2528 ( .A1(n2191), .A2(n1752), .B1(n2256), .B2(n1751), .ZN(n1453)
         );
  OAI22_X1 U2529 ( .A1(n2191), .A2(n1751), .B1(n1750), .B2(n2256), .ZN(n1452)
         );
  OAI22_X1 U2530 ( .A1(n2191), .A2(n1755), .B1(n1754), .B2(n2255), .ZN(n1456)
         );
  XNOR2_X1 U2531 ( .A(n397), .B(n307), .ZN(product[39]) );
  OAI22_X1 U2532 ( .A1(n2004), .A2(n1522), .B1(n1521), .B2(n2238), .ZN(n1232)
         );
  OAI22_X1 U2533 ( .A1(n1955), .A2(n1521), .B1(n2238), .B2(n1520), .ZN(n1231)
         );
  OAI22_X1 U2534 ( .A1(n1956), .A2(n1519), .B1(n2239), .B2(n1518), .ZN(n1229)
         );
  OAI22_X1 U2535 ( .A1(n2005), .A2(n1520), .B1(n1519), .B2(n2238), .ZN(n1230)
         );
  XNOR2_X1 U2536 ( .A(n1237), .B(n1215), .ZN(n939) );
  OR2_X1 U2537 ( .A1(n1215), .A2(n1237), .ZN(n938) );
  OAI22_X1 U2538 ( .A1(n2004), .A2(n1525), .B1(n2238), .B2(n1524), .ZN(n1235)
         );
  OAI22_X1 U2539 ( .A1(n2004), .A2(n1523), .B1(n2239), .B2(n1522), .ZN(n1233)
         );
  OAI22_X1 U2540 ( .A1(n2224), .A2(n1529), .B1(n2239), .B2(n1528), .ZN(n1239)
         );
  OAI22_X1 U2541 ( .A1(n1956), .A2(n1526), .B1(n1525), .B2(n2238), .ZN(n1236)
         );
  OAI22_X1 U2542 ( .A1(n2224), .A2(n1524), .B1(n1523), .B2(n2238), .ZN(n1234)
         );
  OAI22_X1 U2543 ( .A1(n1528), .A2(n2224), .B1(n1527), .B2(n2056), .ZN(n1238)
         );
  OAI22_X1 U2544 ( .A1(n2005), .A2(n1527), .B1(n2239), .B2(n1526), .ZN(n1237)
         );
  OAI22_X1 U2545 ( .A1(n1964), .A2(n1669), .B1(n2250), .B2(n1668), .ZN(n1373)
         );
  OAI22_X1 U2546 ( .A1(n2162), .A2(n1670), .B1(n1669), .B2(n2249), .ZN(n1374)
         );
  OAI22_X1 U2547 ( .A1(n2162), .A2(n1671), .B1(n2249), .B2(n1670), .ZN(n1375)
         );
  OAI22_X1 U2548 ( .A1(n2162), .A2(n1672), .B1(n1671), .B2(n2250), .ZN(n1376)
         );
  OAI22_X1 U2549 ( .A1(n1964), .A2(n1679), .B1(n1974), .B2(n1678), .ZN(n1383)
         );
  OAI22_X1 U2550 ( .A1(n1964), .A2(n1677), .B1(n2249), .B2(n1676), .ZN(n1381)
         );
  OAI22_X1 U2551 ( .A1(n2162), .A2(n1675), .B1(n1974), .B2(n1674), .ZN(n1379)
         );
  OAI22_X1 U2552 ( .A1(n2162), .A2(n1673), .B1(n1974), .B2(n1672), .ZN(n1377)
         );
  OAI22_X1 U2553 ( .A1(n1964), .A2(n1676), .B1(n1675), .B2(n2249), .ZN(n1380)
         );
  OAI22_X1 U2554 ( .A1(n1964), .A2(n1680), .B1(n1679), .B2(n2249), .ZN(n1384)
         );
  OAI22_X1 U2555 ( .A1(n2162), .A2(n1674), .B1(n1673), .B2(n2249), .ZN(n1378)
         );
  OAI22_X1 U2556 ( .A1(n1964), .A2(n1678), .B1(n1677), .B2(n2249), .ZN(n1382)
         );
  XNOR2_X1 U2557 ( .A(b[17]), .B(n2291), .ZN(n1688) );
  XNOR2_X1 U2558 ( .A(b[15]), .B(n2291), .ZN(n1690) );
  XNOR2_X1 U2559 ( .A(b[19]), .B(n2291), .ZN(n1686) );
  XNOR2_X1 U2560 ( .A(b[11]), .B(n2291), .ZN(n1694) );
  XNOR2_X1 U2561 ( .A(b[21]), .B(n2291), .ZN(n1684) );
  XNOR2_X1 U2562 ( .A(b[13]), .B(n2291), .ZN(n1692) );
  AOI21_X1 U2563 ( .B1(n490), .B2(n454), .A(n455), .ZN(n453) );
  OAI21_X1 U2564 ( .B1(n538), .B2(n566), .A(n539), .ZN(n537) );
  XNOR2_X1 U2565 ( .A(n388), .B(n306), .ZN(product[40]) );
  XNOR2_X1 U2566 ( .A(n379), .B(n305), .ZN(product[41]) );
  OAI22_X1 U2567 ( .A1(n2158), .A2(n1637), .B1(n1636), .B2(n2248), .ZN(n1342)
         );
  OAI22_X1 U2568 ( .A1(n1950), .A2(n1636), .B1(n2248), .B2(n1635), .ZN(n1341)
         );
  OAI22_X1 U2569 ( .A1(n1949), .A2(n1634), .B1(n2247), .B2(n1633), .ZN(n1339)
         );
  OAI22_X1 U2570 ( .A1(n1949), .A2(n1635), .B1(n1634), .B2(n2248), .ZN(n1340)
         );
  OAI22_X1 U2571 ( .A1(n1950), .A2(n1639), .B1(n1638), .B2(n2248), .ZN(n1344)
         );
  OAI22_X1 U2572 ( .A1(n1950), .A2(n1640), .B1(n2248), .B2(n1639), .ZN(n1345)
         );
  OAI22_X1 U2573 ( .A1(n2160), .A2(n1642), .B1(n2248), .B2(n1641), .ZN(n1347)
         );
  OAI22_X1 U2574 ( .A1(n2160), .A2(n1633), .B1(n1632), .B2(n2247), .ZN(n772)
         );
  OAI22_X1 U2575 ( .A1(n2159), .A2(n1638), .B1(n2248), .B2(n1637), .ZN(n1343)
         );
  OAI22_X1 U2576 ( .A1(n2099), .A2(n1643), .B1(n1642), .B2(n2247), .ZN(n1348)
         );
  OAI22_X1 U2577 ( .A1(n2159), .A2(n1641), .B1(n1640), .B2(n2248), .ZN(n1346)
         );
  OAI22_X1 U2578 ( .A1(n1656), .A2(n2248), .B1(n1949), .B2(n1993), .ZN(n1188)
         );
  OAI21_X1 U2579 ( .B1(n506), .B2(n452), .A(n453), .ZN(n451) );
  XNOR2_X1 U2580 ( .A(n370), .B(n304), .ZN(product[42]) );
  OAI22_X1 U2581 ( .A1(n1756), .A2(n2255), .B1(n2191), .B2(n2030), .ZN(n1192)
         );
  OAI22_X1 U2582 ( .A1(n2191), .A2(n1738), .B1(n2256), .B2(n1737), .ZN(n1439)
         );
  OAI22_X1 U2583 ( .A1(n2191), .A2(n1741), .B1(n1740), .B2(n2255), .ZN(n1442)
         );
  OAI22_X1 U2584 ( .A1(n2054), .A2(n1739), .B1(n1738), .B2(n2255), .ZN(n1440)
         );
  OAI22_X1 U2585 ( .A1(n2191), .A2(n1740), .B1(n2256), .B2(n1739), .ZN(n1441)
         );
  OAI22_X1 U2586 ( .A1(n2190), .A2(n1736), .B1(n2256), .B2(n1735), .ZN(n1437)
         );
  OAI22_X1 U2587 ( .A1(n2191), .A2(n1742), .B1(n2256), .B2(n1741), .ZN(n1443)
         );
  OAI22_X1 U2588 ( .A1(n2054), .A2(n1735), .B1(n1734), .B2(n2256), .ZN(n1436)
         );
  INV_X1 U2589 ( .A(n916), .ZN(n917) );
  OAI22_X1 U2590 ( .A1(n2232), .A2(n1734), .B1(n2256), .B2(n1733), .ZN(n1435)
         );
  OAI22_X1 U2591 ( .A1(n2190), .A2(n1737), .B1(n1736), .B2(n2256), .ZN(n1438)
         );
  OAI22_X1 U2592 ( .A1(n2054), .A2(n1743), .B1(n1742), .B2(n2255), .ZN(n1444)
         );
  OAI22_X1 U2593 ( .A1(n2232), .A2(n1733), .B1(n1732), .B2(n2255), .ZN(n916)
         );
  NOR2_X1 U2594 ( .A1(n897), .A2(n918), .ZN(n534) );
  OAI22_X1 U2595 ( .A1(n2163), .A2(n1497), .B1(n1496), .B2(n1985), .ZN(n1208)
         );
  OAI22_X1 U2596 ( .A1(n2165), .A2(n1496), .B1(n2236), .B2(n1495), .ZN(n1207)
         );
  OAI22_X1 U2597 ( .A1(n2165), .A2(n1495), .B1(n1494), .B2(n2236), .ZN(n1206)
         );
  OAI22_X1 U2598 ( .A1(n2165), .A2(n1502), .B1(n2237), .B2(n1501), .ZN(n1213)
         );
  OAI22_X1 U2599 ( .A1(n2165), .A2(n1494), .B1(n1985), .B2(n1493), .ZN(n1205)
         );
  OAI22_X1 U2600 ( .A1(n2164), .A2(n1501), .B1(n1500), .B2(n2236), .ZN(n1212)
         );
  OAI22_X1 U2601 ( .A1(n2164), .A2(n1500), .B1(n2237), .B2(n1499), .ZN(n1211)
         );
  XNOR2_X1 U2602 ( .A(b[17]), .B(n2039), .ZN(n1513) );
  OAI22_X1 U2603 ( .A1(n2223), .A2(n1505), .B1(n1504), .B2(n2236), .ZN(n1216)
         );
  OAI22_X1 U2604 ( .A1(n2223), .A2(n1504), .B1(n2237), .B2(n1503), .ZN(n1215)
         );
  OAI22_X1 U2605 ( .A1(n2165), .A2(n1503), .B1(n1502), .B2(n2236), .ZN(n1214)
         );
  OAI22_X1 U2606 ( .A1(n2223), .A2(n1498), .B1(n2236), .B2(n1497), .ZN(n1209)
         );
  OAI22_X1 U2607 ( .A1(n2223), .A2(n1499), .B1(n1498), .B2(n2236), .ZN(n1210)
         );
  XNOR2_X1 U2608 ( .A(b[11]), .B(n2039), .ZN(n1519) );
  XNOR2_X1 U2609 ( .A(b[21]), .B(n2039), .ZN(n1509) );
  XNOR2_X1 U2610 ( .A(b[13]), .B(n2039), .ZN(n1517) );
  XNOR2_X1 U2611 ( .A(b[19]), .B(n2039), .ZN(n1511) );
  XNOR2_X1 U2612 ( .A(b[15]), .B(n2039), .ZN(n1515) );
  XNOR2_X1 U2613 ( .A(n353), .B(n303), .ZN(product[43]) );
  OAI22_X1 U2614 ( .A1(n1964), .A2(n1661), .B1(n2250), .B2(n1660), .ZN(n1365)
         );
  OAI22_X1 U2615 ( .A1(n1964), .A2(n1660), .B1(n1659), .B2(n2250), .ZN(n1364)
         );
  OAI22_X1 U2616 ( .A1(n1681), .A2(n1974), .B1(n2290), .B2(n1964), .ZN(n1189)
         );
  OAI22_X1 U2617 ( .A1(n1964), .A2(n1663), .B1(n2249), .B2(n1662), .ZN(n1367)
         );
  OAI22_X1 U2618 ( .A1(n2162), .A2(n1664), .B1(n1663), .B2(n1974), .ZN(n1368)
         );
  OAI22_X1 U2619 ( .A1(n2162), .A2(n1667), .B1(n1974), .B2(n1666), .ZN(n1371)
         );
  OAI22_X1 U2620 ( .A1(n2162), .A2(n1665), .B1(n2250), .B2(n1664), .ZN(n1369)
         );
  OAI22_X1 U2621 ( .A1(n2162), .A2(n1658), .B1(n1657), .B2(n2249), .ZN(n802)
         );
  OAI22_X1 U2622 ( .A1(n2161), .A2(n1662), .B1(n1661), .B2(n2249), .ZN(n1366)
         );
  OAI22_X1 U2623 ( .A1(n2161), .A2(n1666), .B1(n1665), .B2(n2250), .ZN(n1370)
         );
  OAI22_X1 U2624 ( .A1(n1964), .A2(n1659), .B1(n2249), .B2(n1658), .ZN(n1363)
         );
  OAI22_X1 U2625 ( .A1(n1968), .A2(n1600), .B1(n2243), .B2(n1599), .ZN(n1307)
         );
  OAI22_X1 U2626 ( .A1(n1969), .A2(n1602), .B1(n2243), .B2(n1601), .ZN(n1309)
         );
  OAI22_X1 U2627 ( .A1(n2227), .A2(n1601), .B1(n1600), .B2(n2243), .ZN(n1308)
         );
  OAI22_X1 U2628 ( .A1(n2227), .A2(n1603), .B1(n1602), .B2(n2243), .ZN(n1310)
         );
  OAI22_X1 U2629 ( .A1(n2228), .A2(n1598), .B1(n2244), .B2(n1597), .ZN(n1305)
         );
  OAI22_X1 U2630 ( .A1(n1968), .A2(n1604), .B1(n1961), .B2(n1603), .ZN(n1311)
         );
  OAI22_X1 U2631 ( .A1(n1969), .A2(n1594), .B1(n1960), .B2(n1593), .ZN(n1301)
         );
  OAI22_X1 U2632 ( .A1(n2227), .A2(n1596), .B1(n1960), .B2(n1595), .ZN(n1303)
         );
  OAI22_X1 U2633 ( .A1(n1969), .A2(n1597), .B1(n1596), .B2(n1960), .ZN(n1304)
         );
  OAI22_X1 U2634 ( .A1(n2228), .A2(n1605), .B1(n1604), .B2(n2244), .ZN(n1312)
         );
  OAI22_X1 U2635 ( .A1(n2227), .A2(n1595), .B1(n1594), .B2(n1960), .ZN(n1302)
         );
  OAI22_X1 U2636 ( .A1(n2228), .A2(n1599), .B1(n1598), .B2(n2244), .ZN(n1306)
         );
  XNOR2_X1 U2637 ( .A(b[19]), .B(n2278), .ZN(n1611) );
  XNOR2_X1 U2638 ( .A(b[21]), .B(n2278), .ZN(n1609) );
  XNOR2_X1 U2639 ( .A(b[11]), .B(n2278), .ZN(n1619) );
  XNOR2_X1 U2640 ( .A(b[13]), .B(n2278), .ZN(n1617) );
  XNOR2_X1 U2641 ( .A(b[17]), .B(n2278), .ZN(n1613) );
  XNOR2_X1 U2642 ( .A(b[15]), .B(n2278), .ZN(n1615) );
  NAND2_X1 U2643 ( .A1(n489), .A2(n454), .ZN(n452) );
  NAND2_X1 U2644 ( .A1(n511), .A2(n525), .ZN(n505) );
  INV_X1 U2645 ( .A(n746), .ZN(n747) );
  XNOR2_X1 U2646 ( .A(b[19]), .B(n2283), .ZN(n1636) );
  XNOR2_X1 U2647 ( .A(b[21]), .B(n2285), .ZN(n1634) );
  XNOR2_X1 U2648 ( .A(b[11]), .B(n2283), .ZN(n1644) );
  XNOR2_X1 U2649 ( .A(b[17]), .B(n2284), .ZN(n1638) );
  XNOR2_X1 U2650 ( .A(b[13]), .B(n2283), .ZN(n1642) );
  XNOR2_X1 U2651 ( .A(b[15]), .B(n2283), .ZN(n1640) );
  OAI22_X1 U2652 ( .A1(n1530), .A2(n2224), .B1(n1529), .B2(n2056), .ZN(n1240)
         );
  NAND2_X1 U2653 ( .A1(n540), .A2(n552), .ZN(n538) );
  AOI21_X1 U2654 ( .B1(n540), .B2(n553), .A(n541), .ZN(n539) );
  OAI22_X1 U2655 ( .A1(n2041), .A2(n1544), .B1(n2241), .B2(n1543), .ZN(n1253)
         );
  OAI22_X1 U2656 ( .A1(n2042), .A2(n1552), .B1(n2240), .B2(n1551), .ZN(n1261)
         );
  OAI22_X1 U2657 ( .A1(n2041), .A2(n1548), .B1(n2241), .B2(n1547), .ZN(n1257)
         );
  OAI22_X1 U2658 ( .A1(n2042), .A2(n1547), .B1(n1546), .B2(n2240), .ZN(n1256)
         );
  OAI22_X1 U2659 ( .A1(n2041), .A2(n1546), .B1(n2240), .B2(n1545), .ZN(n1255)
         );
  OAI22_X1 U2660 ( .A1(n2041), .A2(n1555), .B1(n1554), .B2(n2240), .ZN(n1264)
         );
  OAI22_X1 U2661 ( .A1(n2062), .A2(n1549), .B1(n1548), .B2(n2240), .ZN(n1258)
         );
  OAI22_X1 U2662 ( .A1(n2062), .A2(n1550), .B1(n2241), .B2(n1549), .ZN(n1259)
         );
  OAI22_X1 U2663 ( .A1(n2042), .A2(n1545), .B1(n1544), .B2(n2240), .ZN(n1254)
         );
  XNOR2_X1 U2664 ( .A(b[21]), .B(n2273), .ZN(n1559) );
  OAI22_X1 U2665 ( .A1(n2042), .A2(n1554), .B1(n2240), .B2(n1553), .ZN(n1263)
         );
  OAI22_X1 U2666 ( .A1(n2041), .A2(n1551), .B1(n1550), .B2(n2240), .ZN(n1260)
         );
  OAI22_X1 U2667 ( .A1(n2042), .A2(n1553), .B1(n1552), .B2(n2240), .ZN(n1262)
         );
  XNOR2_X1 U2668 ( .A(b[15]), .B(n2271), .ZN(n1565) );
  XNOR2_X1 U2669 ( .A(b[17]), .B(n2272), .ZN(n1563) );
  XNOR2_X1 U2670 ( .A(b[19]), .B(n2271), .ZN(n1561) );
  XNOR2_X1 U2671 ( .A(b[11]), .B(n2272), .ZN(n1569) );
  XNOR2_X1 U2672 ( .A(b[13]), .B(n2272), .ZN(n1567) );
  AOI21_X1 U2673 ( .B1(n346), .B2(n2134), .A(n339), .ZN(n337) );
  OAI21_X1 U2674 ( .B1(n421), .B2(n347), .A(n348), .ZN(n346) );
  NAND2_X1 U2675 ( .A1(n356), .A2(n2133), .ZN(n347) );
  AOI21_X1 U2676 ( .B1(n359), .B2(n2133), .A(n350), .ZN(n348) );
  OAI22_X1 U2677 ( .A1(n2059), .A2(n1608), .B1(n1607), .B2(n2245), .ZN(n746)
         );
  XNOR2_X1 U2678 ( .A(n342), .B(n302), .ZN(product[44]) );
  OAI22_X1 U2679 ( .A1(n2059), .A2(n1620), .B1(n1619), .B2(n2245), .ZN(n1326)
         );
  OAI22_X1 U2680 ( .A1(n2059), .A2(n1626), .B1(n1625), .B2(n2245), .ZN(n1332)
         );
  OAI22_X1 U2681 ( .A1(n2059), .A2(n1623), .B1(n2246), .B2(n1622), .ZN(n1329)
         );
  OAI22_X1 U2682 ( .A1(n2059), .A2(n1630), .B1(n1629), .B2(n2246), .ZN(n1336)
         );
  OAI22_X1 U2683 ( .A1(n2059), .A2(n1625), .B1(n2246), .B2(n1624), .ZN(n1331)
         );
  OAI22_X1 U2684 ( .A1(n2059), .A2(n1629), .B1(n2246), .B2(n1628), .ZN(n1335)
         );
  OAI22_X1 U2685 ( .A1(n2058), .A2(n1621), .B1(n2246), .B2(n1620), .ZN(n1327)
         );
  OAI22_X1 U2686 ( .A1(n2058), .A2(n1619), .B1(n2245), .B2(n1618), .ZN(n1325)
         );
  OAI22_X1 U2687 ( .A1(n2058), .A2(n1624), .B1(n1623), .B2(n2246), .ZN(n1330)
         );
  OAI22_X1 U2688 ( .A1(n2059), .A2(n1627), .B1(n2246), .B2(n1626), .ZN(n1333)
         );
  OAI22_X1 U2689 ( .A1(n2107), .A2(n1622), .B1(n1621), .B2(n2245), .ZN(n1328)
         );
  OAI22_X1 U2690 ( .A1(n2107), .A2(n1628), .B1(n1627), .B2(n2245), .ZN(n1334)
         );
  NOR2_X1 U2691 ( .A1(n505), .A2(n452), .ZN(n450) );
  XOR2_X1 U2692 ( .A(n1952), .B(n321), .Z(product[25]) );
  OAI21_X1 U2693 ( .B1(n1953), .B2(n2086), .A(n2210), .ZN(n533) );
  OAI21_X1 U2694 ( .B1(n1952), .B2(n487), .A(n488), .ZN(n486) );
  OAI21_X1 U2695 ( .B1(n1951), .B2(n463), .A(n464), .ZN(n462) );
  OAI21_X1 U2696 ( .B1(n1953), .B2(n2098), .A(n524), .ZN(n522) );
  OAI21_X1 U2697 ( .B1(n1953), .B2(n476), .A(n477), .ZN(n475) );
  OAI21_X1 U2698 ( .B1(n1951), .B2(n516), .A(n517), .ZN(n515) );
  OAI21_X1 U2699 ( .B1(n1952), .B2(n2053), .A(n2166), .ZN(n504) );
  OAI21_X1 U2700 ( .B1(n1951), .B2(n498), .A(n499), .ZN(n497) );
  OAI22_X1 U2701 ( .A1(n2231), .A2(n1727), .B1(n2253), .B2(n1726), .ZN(n1429)
         );
  OAI22_X1 U2702 ( .A1(n2231), .A2(n1720), .B1(n1719), .B2(n2253), .ZN(n1422)
         );
  OAI22_X1 U2703 ( .A1(n2231), .A2(n1721), .B1(n2253), .B2(n1720), .ZN(n1423)
         );
  OAI22_X1 U2704 ( .A1(n2231), .A2(n1726), .B1(n1725), .B2(n2253), .ZN(n1428)
         );
  OAI22_X1 U2705 ( .A1(n2231), .A2(n1730), .B1(n1729), .B2(n2254), .ZN(n1432)
         );
  OAI22_X1 U2706 ( .A1(n1725), .A2(n2108), .B1(n2253), .B2(n1724), .ZN(n1427)
         );
  OAI22_X1 U2707 ( .A1(n2108), .A2(n1723), .B1(n2254), .B2(n1722), .ZN(n1425)
         );
  OAI22_X1 U2708 ( .A1(n2231), .A2(n1728), .B1(n1727), .B2(n2253), .ZN(n1430)
         );
  OAI22_X1 U2709 ( .A1(n2108), .A2(n1729), .B1(n2254), .B2(n1728), .ZN(n1431)
         );
  OAI22_X1 U2710 ( .A1(n2108), .A2(n1722), .B1(n1721), .B2(n2253), .ZN(n1424)
         );
  OAI22_X1 U2711 ( .A1(n2108), .A2(n1719), .B1(n2253), .B2(n1718), .ZN(n1421)
         );
  OAI22_X1 U2712 ( .A1(n2108), .A2(n1724), .B1(n1723), .B2(n2253), .ZN(n1426)
         );
  XNOR2_X1 U2713 ( .A(b[15]), .B(n2300), .ZN(n1740) );
  XNOR2_X1 U2714 ( .A(b[21]), .B(n2300), .ZN(n1734) );
  XNOR2_X1 U2715 ( .A(b[19]), .B(n2299), .ZN(n1736) );
  XNOR2_X1 U2716 ( .A(b[11]), .B(n2299), .ZN(n1744) );
  XNOR2_X1 U2717 ( .A(b[17]), .B(n2299), .ZN(n1738) );
  XNOR2_X1 U2718 ( .A(b[13]), .B(n2300), .ZN(n1742) );
  INV_X1 U2719 ( .A(n325), .ZN(product[47]) );
  AOI21_X1 U2720 ( .B1(n423), .B2(n356), .A(n359), .ZN(n355) );
  NAND2_X1 U2721 ( .A1(n422), .A2(n356), .ZN(n354) );
  OAI22_X1 U2722 ( .A1(n1990), .A2(n1563), .B1(n2038), .B2(n1562), .ZN(n1271)
         );
  OAI22_X1 U2723 ( .A1(n1991), .A2(n1567), .B1(n1984), .B2(n1566), .ZN(n1275)
         );
  OAI22_X1 U2724 ( .A1(n1991), .A2(n1566), .B1(n1565), .B2(n2038), .ZN(n1274)
         );
  OAI22_X1 U2725 ( .A1(n1979), .A2(n1561), .B1(n2038), .B2(n1560), .ZN(n1269)
         );
  OAI22_X1 U2726 ( .A1(n1990), .A2(n1564), .B1(n1563), .B2(n1984), .ZN(n1272)
         );
  OAI22_X1 U2727 ( .A1(n2225), .A2(n1560), .B1(n1559), .B2(n2038), .ZN(n1268)
         );
  OAI22_X1 U2728 ( .A1(n1991), .A2(n1565), .B1(n2242), .B2(n1564), .ZN(n1273)
         );
  OAI22_X1 U2729 ( .A1(n1991), .A2(n1559), .B1(n2038), .B2(n1558), .ZN(n1267)
         );
  OAI22_X1 U2730 ( .A1(n1581), .A2(n2038), .B1(n1979), .B2(n1994), .ZN(n1185)
         );
  OAI22_X1 U2731 ( .A1(n1990), .A2(n1562), .B1(n1561), .B2(n2038), .ZN(n1270)
         );
  OAI22_X1 U2732 ( .A1(n2226), .A2(n1568), .B1(n1567), .B2(n1984), .ZN(n1276)
         );
  XNOR2_X1 U2733 ( .A(b[17]), .B(n2275), .ZN(n1588) );
  XNOR2_X1 U2734 ( .A(b[15]), .B(n2276), .ZN(n1590) );
  XNOR2_X1 U2735 ( .A(b[13]), .B(n2276), .ZN(n1592) );
  OAI22_X1 U2736 ( .A1(n2225), .A2(n1558), .B1(n1557), .B2(n2038), .ZN(n706)
         );
  XNOR2_X1 U2737 ( .A(b[19]), .B(n2275), .ZN(n1586) );
  XNOR2_X1 U2738 ( .A(b[21]), .B(n2275), .ZN(n1584) );
  XNOR2_X1 U2739 ( .A(b[11]), .B(n2276), .ZN(n1594) );
  OAI21_X1 U2740 ( .B1(n326), .B2(n2106), .A(n327), .ZN(n325) );
  NAND2_X1 U2741 ( .A1(n2192), .A2(n474), .ZN(n314) );
  OAI21_X1 U2742 ( .B1(n2106), .B2(n431), .A(n432), .ZN(n430) );
  OAI21_X1 U2743 ( .B1(n301), .B2(n420), .A(n421), .ZN(n419) );
  OAI21_X1 U2744 ( .B1(n301), .B2(n438), .A(n439), .ZN(n437) );
  OAI21_X1 U2745 ( .B1(n301), .B2(n411), .A(n412), .ZN(n410) );
  OAI21_X1 U2746 ( .B1(n2106), .B2(n354), .A(n355), .ZN(n353) );
  OAI21_X1 U2747 ( .B1(n301), .B2(n371), .A(n372), .ZN(n370) );
  OAI21_X1 U2748 ( .B1(n301), .B2(n380), .A(n381), .ZN(n379) );
  OAI21_X1 U2749 ( .B1(n2106), .B2(n343), .A(n344), .ZN(n342) );
  OAI21_X1 U2750 ( .B1(n2106), .B2(n398), .A(n399), .ZN(n397) );
  OAI21_X1 U2751 ( .B1(n301), .B2(n389), .A(n390), .ZN(n388) );
  AOI21_X1 U2752 ( .B1(n2192), .B2(n483), .A(n472), .ZN(n468) );
  NAND2_X1 U2753 ( .A1(n1975), .A2(n2192), .ZN(n467) );
  OAI22_X1 U2754 ( .A1(n2071), .A2(n1691), .B1(n1690), .B2(n2251), .ZN(n1394)
         );
  OAI22_X1 U2755 ( .A1(n2070), .A2(n1686), .B1(n2252), .B2(n1685), .ZN(n1389)
         );
  OAI22_X1 U2756 ( .A1(n2070), .A2(n1689), .B1(n1688), .B2(n2252), .ZN(n1392)
         );
  OAI22_X1 U2757 ( .A1(n2071), .A2(n1690), .B1(n2252), .B2(n1689), .ZN(n1393)
         );
  OAI22_X1 U2758 ( .A1(n2193), .A2(n1687), .B1(n1686), .B2(n2252), .ZN(n1390)
         );
  OAI22_X1 U2759 ( .A1(n2193), .A2(n1692), .B1(n2252), .B2(n1691), .ZN(n1395)
         );
  OAI22_X1 U2760 ( .A1(n2070), .A2(n1685), .B1(n1684), .B2(n2251), .ZN(n1388)
         );
  OAI22_X1 U2761 ( .A1(n2193), .A2(n1688), .B1(n2251), .B2(n1687), .ZN(n1391)
         );
  OAI22_X1 U2762 ( .A1(n2193), .A2(n1684), .B1(n2252), .B2(n1683), .ZN(n1387)
         );
  OAI22_X1 U2763 ( .A1(n1706), .A2(n2252), .B1(n2071), .B2(n2295), .ZN(n1190)
         );
  XNOR2_X1 U2764 ( .A(b[13]), .B(n2297), .ZN(n1717) );
  XNOR2_X1 U2765 ( .A(b[21]), .B(n2296), .ZN(n1709) );
  XNOR2_X1 U2766 ( .A(b[15]), .B(n2297), .ZN(n1715) );
  XNOR2_X1 U2767 ( .A(b[11]), .B(n2296), .ZN(n1719) );
  XNOR2_X1 U2768 ( .A(b[19]), .B(n2296), .ZN(n1711) );
  XNOR2_X1 U2769 ( .A(b[17]), .B(n2297), .ZN(n1713) );
  INV_X2 U2770 ( .A(n2147), .ZN(n2227) );
  INV_X1 U2771 ( .A(n2000), .ZN(n2237) );
  INV_X1 U2772 ( .A(n2203), .ZN(n2239) );
  INV_X1 U2773 ( .A(n1988), .ZN(n2250) );
  INV_X1 U2774 ( .A(n1983), .ZN(n2252) );
  INV_X1 U2775 ( .A(n2144), .ZN(n2256) );
  INV_X1 U2776 ( .A(n2172), .ZN(n2269) );
  INV_X1 U2777 ( .A(n2037), .ZN(n2281) );
  INV_X1 U2778 ( .A(n2286), .ZN(n2285) );
  INV_X1 U2779 ( .A(n2290), .ZN(n2289) );
  INV_X1 U2780 ( .A(n2295), .ZN(n2294) );
  INV_X1 U2781 ( .A(n2030), .ZN(n2299) );
  INV_X1 U2782 ( .A(n2052), .ZN(n2304) );
  INV_X2 U2783 ( .A(b[0]), .ZN(n2305) );
endmodule


module iir_filter_DW_mult_tc_2 ( a, b, product );
  input [23:0] a;
  input [23:0] b;
  output [47:0] product;
  wire   n251, n267, n277, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n325, n326, n327, n332, n333, n334, n335, n336, n337, n339,
         n341, n342, n343, n344, n345, n346, n347, n348, n350, n352, n353,
         n354, n355, n356, n359, n360, n361, n362, n363, n364, n365, n367,
         n369, n370, n371, n372, n376, n378, n379, n380, n381, n382, n383,
         n384, n387, n388, n389, n390, n394, n396, n397, n398, n399, n400,
         n401, n402, n405, n407, n409, n410, n411, n412, n416, n418, n419,
         n420, n421, n422, n423, n426, n427, n428, n429, n430, n431, n432,
         n434, n435, n436, n437, n438, n439, n445, n450, n451, n452, n453,
         n454, n455, n456, n457, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n483, n486, n487, n488, n489, n490, n492, n495, n496,
         n497, n498, n499, n501, n502, n503, n504, n505, n506, n507, n508,
         n511, n512, n513, n514, n515, n516, n517, n519, n520, n521, n522,
         n524, n525, n526, n531, n532, n533, n534, n535, n536, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n550, n551, n552,
         n553, n554, n555, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n581, n582, n583, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n609, n610, n611, n620, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n643, n644, n645,
         n646, n657, n661, n662, n663, n665, n666, n667, n668, n670, n672,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1807, n1809, n1813,
         n1817, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338;

  FA_X1 U546 ( .A(n1195), .B(n682), .CI(n1218), .CO(n678), .S(n679) );
  FA_X1 U547 ( .A(n683), .B(n1196), .CI(n686), .CO(n680), .S(n681) );
  FA_X1 U549 ( .A(n690), .B(n1242), .CI(n687), .CO(n684), .S(n685) );
  FA_X1 U550 ( .A(n1219), .B(n692), .CI(n1197), .CO(n686), .S(n687) );
  FA_X1 U551 ( .A(n691), .B(n698), .CI(n696), .CO(n688), .S(n689) );
  FA_X1 U552 ( .A(n1198), .B(n1220), .CI(n693), .CO(n690), .S(n691) );
  FA_X1 U554 ( .A(n702), .B(n699), .CI(n697), .CO(n694), .S(n695) );
  FA_X1 U555 ( .A(n1266), .B(n1243), .CI(n704), .CO(n696), .S(n697) );
  FA_X1 U556 ( .A(n1221), .B(n1199), .CI(n706), .CO(n698), .S(n699) );
  FA_X1 U557 ( .A(n710), .B(n712), .CI(n703), .CO(n700), .S(n701) );
  FA_X1 U558 ( .A(n714), .B(n1244), .CI(n705), .CO(n702), .S(n703) );
  FA_X1 U559 ( .A(n1222), .B(n1200), .CI(n707), .CO(n704), .S(n705) );
  FA_X1 U561 ( .A(n718), .B(n713), .CI(n711), .CO(n708), .S(n709) );
  FA_X1 U562 ( .A(n715), .B(n722), .CI(n720), .CO(n710), .S(n711) );
  FA_X1 U563 ( .A(n1245), .B(n1223), .CI(n1290), .CO(n712), .S(n713) );
  FA_X1 U564 ( .A(n1267), .B(n1201), .CI(n724), .CO(n714), .S(n715) );
  FA_X1 U565 ( .A(n728), .B(n721), .CI(n719), .CO(n716), .S(n717) );
  FA_X1 U566 ( .A(n723), .B(n732), .CI(n730), .CO(n718), .S(n719) );
  FA_X1 U567 ( .A(n1202), .B(n1246), .CI(n734), .CO(n720), .S(n721) );
  FA_X1 U568 ( .A(n1268), .B(n1224), .CI(n725), .CO(n722), .S(n723) );
  FA_X1 U570 ( .A(n738), .B(n731), .CI(n729), .CO(n726), .S(n727) );
  FA_X1 U571 ( .A(n735), .B(n733), .CI(n740), .CO(n728), .S(n729) );
  FA_X1 U572 ( .A(n744), .B(n1314), .CI(n742), .CO(n730), .S(n731) );
  FA_X1 U573 ( .A(n1225), .B(n1291), .CI(n1269), .CO(n732), .S(n733) );
  FA_X1 U574 ( .A(n746), .B(n1203), .CI(n1247), .CO(n734), .S(n735) );
  FA_X1 U575 ( .A(n750), .B(n741), .CI(n739), .CO(n736), .S(n737) );
  FA_X1 U576 ( .A(n754), .B(n745), .CI(n752), .CO(n738), .S(n739) );
  FA_X1 U577 ( .A(n756), .B(n758), .CI(n743), .CO(n740), .S(n741) );
  FA_X1 U578 ( .A(n1226), .B(n1204), .CI(n1270), .CO(n742), .S(n743) );
  FA_X1 U579 ( .A(n1292), .B(n1248), .CI(n747), .CO(n744), .S(n745) );
  FA_X1 U581 ( .A(n762), .B(n753), .CI(n751), .CO(n748), .S(n749) );
  FA_X1 U582 ( .A(n755), .B(n766), .CI(n764), .CO(n750), .S(n751) );
  FA_X1 U583 ( .A(n757), .B(n768), .CI(n759), .CO(n752), .S(n753) );
  FA_X1 U584 ( .A(n1338), .B(n1271), .CI(n770), .CO(n754), .S(n755) );
  FA_X1 U585 ( .A(n1249), .B(n1293), .CI(n1315), .CO(n756), .S(n757) );
  FA_X1 U586 ( .A(n772), .B(n1205), .CI(n1227), .CO(n758), .S(n759) );
  FA_X1 U587 ( .A(n776), .B(n765), .CI(n763), .CO(n760), .S(n761) );
  FA_X1 U588 ( .A(n767), .B(n780), .CI(n778), .CO(n762), .S(n763) );
  FA_X1 U589 ( .A(n771), .B(n769), .CI(n782), .CO(n764), .S(n765) );
  FA_X1 U590 ( .A(n786), .B(n1228), .CI(n784), .CO(n766), .S(n767) );
  FA_X1 U591 ( .A(n1294), .B(n1206), .CI(n1272), .CO(n768), .S(n769) );
  FA_X1 U592 ( .A(n1316), .B(n1250), .CI(n773), .CO(n770), .S(n771) );
  FA_X1 U594 ( .A(n790), .B(n779), .CI(n777), .CO(n774), .S(n775) );
  FA_X1 U595 ( .A(n781), .B(n794), .CI(n792), .CO(n776), .S(n777) );
  FA_X1 U596 ( .A(n783), .B(n787), .CI(n796), .CO(n778), .S(n779) );
  FA_X1 U597 ( .A(n798), .B(n800), .CI(n785), .CO(n780), .S(n781) );
  FA_X1 U598 ( .A(n1339), .B(n1229), .CI(n1362), .CO(n782), .S(n783) );
  FA_X1 U599 ( .A(n1273), .B(n1295), .CI(n1317), .CO(n784), .S(n785) );
  FA_X1 U600 ( .A(n1251), .B(n1207), .CI(n1996), .CO(n786), .S(n787) );
  FA_X1 U601 ( .A(n806), .B(n793), .CI(n791), .CO(n788), .S(n789) );
  FA_X1 U602 ( .A(n795), .B(n810), .CI(n808), .CO(n790), .S(n791) );
  FA_X1 U603 ( .A(n801), .B(n797), .CI(n812), .CO(n792), .S(n793) );
  FA_X1 U604 ( .A(n814), .B(n816), .CI(n799), .CO(n794), .S(n795) );
  FA_X1 U606 ( .A(n1208), .B(n1318), .CI(n1230), .CO(n798), .S(n799) );
  FA_X1 U607 ( .A(n1340), .B(n1252), .CI(n803), .CO(n800), .S(n801) );
  FA_X1 U609 ( .A(n822), .B(n809), .CI(n807), .CO(n804), .S(n805) );
  FA_X1 U610 ( .A(n811), .B(n826), .CI(n824), .CO(n806), .S(n807) );
  FA_X1 U611 ( .A(n828), .B(n819), .CI(n813), .CO(n808), .S(n809) );
  FA_X1 U612 ( .A(n815), .B(n832), .CI(n817), .CO(n810), .S(n811) );
  FA_X1 U613 ( .A(n830), .B(n1386), .CI(n834), .CO(n812), .S(n813) );
  FA_X1 U614 ( .A(n1319), .B(n1253), .CI(n1341), .CO(n814), .S(n815) );
  FA_X1 U615 ( .A(n1231), .B(n1297), .CI(n1275), .CO(n816), .S(n817) );
  FA_X1 U616 ( .A(n1209), .B(n1363), .CI(n2026), .CO(n818), .S(n819) );
  FA_X1 U617 ( .A(n840), .B(n825), .CI(n823), .CO(n820), .S(n821) );
  FA_X1 U619 ( .A(n846), .B(n848), .CI(n829), .CO(n824), .S(n825) );
  FA_X1 U620 ( .A(n835), .B(n831), .CI(n833), .CO(n826), .S(n827) );
  FA_X1 U621 ( .A(n850), .B(n854), .CI(n852), .CO(n828), .S(n829) );
  FA_X1 U622 ( .A(n1298), .B(n1320), .CI(n1254), .CO(n830), .S(n831) );
  FA_X1 U623 ( .A(n1232), .B(n1364), .CI(n1342), .CO(n832), .S(n833) );
  FA_X1 U624 ( .A(n1210), .B(n1276), .CI(n837), .CO(n834), .S(n835) );
  FA_X1 U626 ( .A(n858), .B(n843), .CI(n841), .CO(n838), .S(n839) );
  FA_X1 U627 ( .A(n845), .B(n847), .CI(n860), .CO(n840), .S(n841) );
  FA_X1 U628 ( .A(n864), .B(n849), .CI(n862), .CO(n842), .S(n843) );
  FA_X1 U629 ( .A(n855), .B(n853), .CI(n866), .CO(n844), .S(n845) );
  FA_X1 U630 ( .A(n868), .B(n870), .CI(n851), .CO(n846), .S(n847) );
  FA_X1 U631 ( .A(n1410), .B(n1365), .CI(n872), .CO(n848), .S(n849) );
  FA_X1 U632 ( .A(n1343), .B(n1277), .CI(n1299), .CO(n850), .S(n851) );
  FA_X1 U633 ( .A(n1255), .B(n1321), .CI(n874), .CO(n852), .S(n853) );
  FA_X1 U634 ( .A(n1387), .B(n1211), .CI(n1233), .CO(n854), .S(n855) );
  FA_X1 U635 ( .A(n878), .B(n861), .CI(n859), .CO(n856), .S(n857) );
  FA_X1 U637 ( .A(n884), .B(n867), .CI(n865), .CO(n860), .S(n861) );
  FA_X1 U639 ( .A(n869), .B(n890), .CI(n871), .CO(n864), .S(n865) );
  FA_X1 U640 ( .A(n894), .B(n1300), .CI(n892), .CO(n866), .S(n867) );
  FA_X1 U641 ( .A(n1234), .B(n1256), .CI(n1322), .CO(n868), .S(n869) );
  FA_X1 U642 ( .A(n1344), .B(n1366), .CI(n1212), .CO(n870), .S(n871) );
  FA_X1 U643 ( .A(n1388), .B(n1278), .CI(n875), .CO(n872), .S(n873) );
  FA_X1 U645 ( .A(n898), .B(n881), .CI(n879), .CO(n876), .S(n877) );
  FA_X1 U646 ( .A(n883), .B(n885), .CI(n900), .CO(n878), .S(n879) );
  FA_X1 U651 ( .A(n1367), .B(n1389), .CI(n1434), .CO(n888), .S(n889) );
  FA_X1 U652 ( .A(n1257), .B(n1301), .CI(n1345), .CO(n890), .S(n891) );
  FA_X1 U653 ( .A(n2237), .B(n1279), .CI(n1323), .CO(n892), .S(n893) );
  FA_X1 U654 ( .A(n1411), .B(n1213), .CI(n1235), .CO(n894), .S(n895) );
  FA_X1 U655 ( .A(n920), .B(n901), .CI(n899), .CO(n896), .S(n897) );
  FA_X1 U656 ( .A(n903), .B(n924), .CI(n922), .CO(n898), .S(n899) );
  FA_X1 U657 ( .A(n907), .B(n926), .CI(n905), .CO(n900), .S(n901) );
  FA_X1 U658 ( .A(n909), .B(n930), .CI(n928), .CO(n902), .S(n903) );
  FA_X1 U659 ( .A(n913), .B(n911), .CI(n915), .CO(n904), .S(n905) );
  FA_X1 U660 ( .A(n932), .B(n936), .CI(n934), .CO(n906), .S(n907) );
  FA_X1 U661 ( .A(n1368), .B(n1390), .CI(n938), .CO(n908), .S(n909) );
  FA_X1 U662 ( .A(n1280), .B(n1346), .CI(n1324), .CO(n910), .S(n911) );
  FA_X1 U663 ( .A(n1236), .B(n1412), .CI(n1258), .CO(n912), .S(n913) );
  FA_X1 U664 ( .A(n1214), .B(n1302), .CI(n917), .CO(n914), .S(n915) );
  FA_X1 U667 ( .A(n925), .B(n927), .CI(n944), .CO(n920), .S(n921) );
  FA_X1 U668 ( .A(n929), .B(n948), .CI(n946), .CO(n922), .S(n923) );
  FA_X1 U669 ( .A(n950), .B(n935), .CI(n931), .CO(n924), .S(n925) );
  FA_X1 U670 ( .A(n937), .B(n933), .CI(n952), .CO(n926), .S(n927) );
  FA_X1 U671 ( .A(n954), .B(n958), .CI(n956), .CO(n928), .S(n929) );
  FA_X1 U672 ( .A(n939), .B(n960), .CI(n1458), .CO(n930), .S(n931) );
  FA_X1 U673 ( .A(n1325), .B(n1435), .CI(n1413), .CO(n932), .S(n933) );
  FA_X1 U674 ( .A(n1281), .B(n1369), .CI(n1391), .CO(n934), .S(n935) );
  FA_X1 U675 ( .A(n1259), .B(n1303), .CI(n1347), .CO(n936), .S(n937) );
  FA_X1 U678 ( .A(n964), .B(n945), .CI(n943), .CO(n940), .S(n941) );
  FA_X1 U679 ( .A(n947), .B(n949), .CI(n966), .CO(n942), .S(n943) );
  FA_X1 U680 ( .A(n951), .B(n970), .CI(n968), .CO(n944), .S(n945) );
  FA_X1 U681 ( .A(n972), .B(n959), .CI(n953), .CO(n946), .S(n947) );
  FA_X1 U682 ( .A(n955), .B(n974), .CI(n957), .CO(n948), .S(n949) );
  FA_X1 U683 ( .A(n978), .B(n980), .CI(n976), .CO(n950), .S(n951) );
  FA_X1 U685 ( .A(n1282), .B(n1414), .CI(n1304), .CO(n954), .S(n955) );
  FA_X1 U686 ( .A(n1436), .B(n1459), .CI(n1370), .CO(n956), .S(n957) );
  FA_X1 U687 ( .A(n1348), .B(n1260), .CI(n1182), .CO(n958), .S(n959) );
  HA_X1 U688 ( .A(n1238), .B(n1939), .CO(n960), .S(n961) );
  FA_X1 U689 ( .A(n984), .B(n967), .CI(n965), .CO(n962), .S(n963) );
  FA_X1 U690 ( .A(n969), .B(n971), .CI(n986), .CO(n964), .S(n965) );
  FA_X1 U691 ( .A(n973), .B(n990), .CI(n988), .CO(n966), .S(n967) );
  FA_X1 U692 ( .A(n975), .B(n981), .CI(n992), .CO(n968), .S(n969) );
  FA_X1 U693 ( .A(n977), .B(n998), .CI(n979), .CO(n970), .S(n971) );
  FA_X1 U695 ( .A(n1393), .B(n1415), .CI(n1000), .CO(n974), .S(n975) );
  FA_X1 U696 ( .A(n1305), .B(n1437), .CI(n1327), .CO(n976), .S(n977) );
  FA_X1 U697 ( .A(n1460), .B(n1371), .CI(n1283), .CO(n978), .S(n979) );
  FA_X1 U698 ( .A(n1239), .B(n1349), .CI(n1261), .CO(n980), .S(n981) );
  FA_X1 U699 ( .A(n1004), .B(n987), .CI(n985), .CO(n982), .S(n983) );
  FA_X1 U700 ( .A(n989), .B(n991), .CI(n1006), .CO(n984), .S(n985) );
  FA_X1 U701 ( .A(n993), .B(n1010), .CI(n1008), .CO(n986), .S(n987) );
  FA_X1 U703 ( .A(n1014), .B(n1016), .CI(n995), .CO(n990), .S(n991) );
  FA_X1 U704 ( .A(n1001), .B(n1394), .CI(n1018), .CO(n992), .S(n993) );
  HA_X1 U708 ( .A(n1262), .B(n1240), .CO(n1000), .S(n1001) );
  FA_X1 U709 ( .A(n1022), .B(n1007), .CI(n1005), .CO(n1002), .S(n1003) );
  FA_X1 U710 ( .A(n1009), .B(n1011), .CI(n1024), .CO(n1004), .S(n1005) );
  FA_X1 U711 ( .A(n1013), .B(n1028), .CI(n1026), .CO(n1006), .S(n1007) );
  FA_X1 U712 ( .A(n1015), .B(n1019), .CI(n1017), .CO(n1008), .S(n1009) );
  FA_X1 U713 ( .A(n1030), .B(n1034), .CI(n1241), .CO(n1010), .S(n1011) );
  FA_X1 U714 ( .A(n1036), .B(n1439), .CI(n1032), .CO(n1012), .S(n1013) );
  FA_X1 U716 ( .A(n1307), .B(n1329), .CI(n1373), .CO(n1016), .S(n1017) );
  FA_X1 U717 ( .A(n1285), .B(n1351), .CI(n1263), .CO(n1018), .S(n1019) );
  FA_X1 U718 ( .A(n1040), .B(n1025), .CI(n1023), .CO(n1020), .S(n1021) );
  FA_X1 U719 ( .A(n1027), .B(n1044), .CI(n1042), .CO(n1022), .S(n1023) );
  FA_X1 U720 ( .A(n1046), .B(n1035), .CI(n1029), .CO(n1024), .S(n1025) );
  FA_X1 U722 ( .A(n1052), .B(n1037), .CI(n1050), .CO(n1028), .S(n1029) );
  FA_X1 U723 ( .A(n1352), .B(n1440), .CI(n1418), .CO(n1030), .S(n1031) );
  FA_X1 U724 ( .A(n1330), .B(n1463), .CI(n1396), .CO(n1032), .S(n1033) );
  FA_X1 U725 ( .A(n1308), .B(n1374), .CI(n1184), .CO(n1034), .S(n1035) );
  HA_X1 U726 ( .A(n1264), .B(n1286), .CO(n1036), .S(n1037) );
  FA_X1 U728 ( .A(n1058), .B(n1047), .CI(n1045), .CO(n1040), .S(n1041) );
  FA_X1 U730 ( .A(n1049), .B(n1265), .CI(n1051), .CO(n1044), .S(n1045) );
  FA_X1 U731 ( .A(n1064), .B(n1068), .CI(n1066), .CO(n1046), .S(n1047) );
  FA_X1 U732 ( .A(n1397), .B(n1441), .CI(n1419), .CO(n1048), .S(n1049) );
  FA_X1 U733 ( .A(n1331), .B(n1353), .CI(n1375), .CO(n1050), .S(n1051) );
  FA_X1 U734 ( .A(n1287), .B(n1464), .CI(n1309), .CO(n1052), .S(n1053) );
  FA_X1 U735 ( .A(n1072), .B(n1059), .CI(n1057), .CO(n1054), .S(n1055) );
  FA_X1 U736 ( .A(n1074), .B(n1063), .CI(n1061), .CO(n1056), .S(n1057) );
  FA_X1 U737 ( .A(n1067), .B(n1065), .CI(n1076), .CO(n1058), .S(n1059) );
  FA_X1 U739 ( .A(n1398), .B(n1420), .CI(n1069), .CO(n1062), .S(n1063) );
  FA_X1 U740 ( .A(n1442), .B(n1354), .CI(n1332), .CO(n1064), .S(n1065) );
  FA_X1 U741 ( .A(n1465), .B(n1376), .CI(n1185), .CO(n1066), .S(n1067) );
  HA_X1 U742 ( .A(n1288), .B(n1310), .CO(n1068), .S(n1069) );
  FA_X1 U743 ( .A(n1086), .B(n1075), .CI(n1073), .CO(n1070), .S(n1071) );
  FA_X1 U744 ( .A(n1088), .B(n1090), .CI(n1077), .CO(n1072), .S(n1073) );
  FA_X1 U745 ( .A(n1083), .B(n1081), .CI(n1079), .CO(n1074), .S(n1075) );
  FA_X1 U746 ( .A(n1092), .B(n1094), .CI(n1289), .CO(n1076), .S(n1077) );
  FA_X1 U748 ( .A(n1355), .B(n1443), .CI(n1377), .CO(n1080), .S(n1081) );
  FA_X1 U749 ( .A(n1311), .B(n1466), .CI(n1333), .CO(n1082), .S(n1083) );
  FA_X1 U750 ( .A(n1100), .B(n1089), .CI(n1087), .CO(n1084), .S(n1085) );
  FA_X1 U751 ( .A(n1102), .B(n1104), .CI(n1091), .CO(n1086), .S(n1087) );
  FA_X1 U752 ( .A(n1093), .B(n1106), .CI(n1095), .CO(n1088), .S(n1089) );
  FA_X1 U753 ( .A(n1097), .B(n1422), .CI(n1108), .CO(n1090), .S(n1091) );
  FA_X1 U754 ( .A(n1356), .B(n1444), .CI(n1378), .CO(n1092), .S(n1093) );
  FA_X1 U755 ( .A(n1186), .B(n1467), .CI(n1400), .CO(n1094), .S(n1095) );
  HA_X1 U756 ( .A(n1334), .B(n1312), .CO(n1096), .S(n1097) );
  FA_X1 U757 ( .A(n1103), .B(n1112), .CI(n1101), .CO(n1098), .S(n1099) );
  FA_X1 U758 ( .A(n1114), .B(n1109), .CI(n1105), .CO(n1100), .S(n1101) );
  FA_X1 U759 ( .A(n1313), .B(n1116), .CI(n1107), .CO(n1102), .S(n1103) );
  FA_X1 U760 ( .A(n1120), .B(n1423), .CI(n1118), .CO(n1104), .S(n1105) );
  FA_X1 U761 ( .A(n1379), .B(n1445), .CI(n1401), .CO(n1106), .S(n1107) );
  FA_X1 U762 ( .A(n1335), .B(n1468), .CI(n1357), .CO(n1108), .S(n1109) );
  FA_X1 U763 ( .A(n1124), .B(n1115), .CI(n1113), .CO(n1110), .S(n1111) );
  FA_X1 U764 ( .A(n1119), .B(n1117), .CI(n1126), .CO(n1112), .S(n1113) );
  FA_X1 U765 ( .A(n1130), .B(n1121), .CI(n1128), .CO(n1114), .S(n1115) );
  FA_X1 U766 ( .A(n1380), .B(n1446), .CI(n1424), .CO(n1116), .S(n1117) );
  FA_X1 U767 ( .A(n1469), .B(n1402), .CI(n1187), .CO(n1118), .S(n1119) );
  HA_X1 U768 ( .A(n1336), .B(n1358), .CO(n1120), .S(n1121) );
  FA_X1 U769 ( .A(n1127), .B(n1134), .CI(n1125), .CO(n1122), .S(n1123) );
  FA_X1 U770 ( .A(n1131), .B(n1129), .CI(n1136), .CO(n1124), .S(n1125) );
  FA_X1 U771 ( .A(n1138), .B(n1140), .CI(n1337), .CO(n1126), .S(n1127) );
  FA_X1 U772 ( .A(n1403), .B(n1447), .CI(n1425), .CO(n1128), .S(n1129) );
  FA_X1 U773 ( .A(n1359), .B(n1470), .CI(n1381), .CO(n1130), .S(n1131) );
  FA_X1 U774 ( .A(n1144), .B(n1137), .CI(n1135), .CO(n1132), .S(n1133) );
  FA_X1 U775 ( .A(n1146), .B(n1148), .CI(n1139), .CO(n1134), .S(n1135) );
  FA_X1 U776 ( .A(n1404), .B(n1448), .CI(n1141), .CO(n1136), .S(n1137) );
  FA_X1 U777 ( .A(n1471), .B(n1426), .CI(n1188), .CO(n1138), .S(n1139) );
  HA_X1 U778 ( .A(n1360), .B(n1382), .CO(n1140), .S(n1141) );
  FA_X1 U779 ( .A(n1152), .B(n1147), .CI(n1145), .CO(n1142), .S(n1143) );
  FA_X1 U780 ( .A(n1361), .B(n1154), .CI(n1149), .CO(n1144), .S(n1145) );
  FA_X1 U781 ( .A(n1427), .B(n1449), .CI(n1156), .CO(n1146), .S(n1147) );
  FA_X1 U782 ( .A(n1383), .B(n1472), .CI(n1405), .CO(n1148), .S(n1149) );
  FA_X1 U783 ( .A(n1160), .B(n1155), .CI(n1153), .CO(n1150), .S(n1151) );
  FA_X1 U784 ( .A(n1157), .B(n1473), .CI(n1162), .CO(n1152), .S(n1153) );
  FA_X1 U785 ( .A(n1450), .B(n1428), .CI(n1189), .CO(n1154), .S(n1155) );
  HA_X1 U786 ( .A(n1384), .B(n1406), .CO(n1156), .S(n1157) );
  FA_X1 U787 ( .A(n1163), .B(n1385), .CI(n1164), .CO(n1158), .S(n1159) );
  FA_X1 U788 ( .A(n1168), .B(n1429), .CI(n1166), .CO(n1160), .S(n1161) );
  FA_X1 U789 ( .A(n1407), .B(n1474), .CI(n1451), .CO(n1162), .S(n1163) );
  FA_X1 U790 ( .A(n1172), .B(n1169), .CI(n1167), .CO(n1164), .S(n1165) );
  FA_X1 U791 ( .A(n1452), .B(n1475), .CI(n1190), .CO(n1166), .S(n1167) );
  HA_X1 U792 ( .A(n1408), .B(n1430), .CO(n1168), .S(n1169) );
  FA_X1 U793 ( .A(n1409), .B(n1176), .CI(n1173), .CO(n1170), .S(n1171) );
  FA_X1 U794 ( .A(n1476), .B(n1453), .CI(n1431), .CO(n1172), .S(n1173) );
  FA_X1 U795 ( .A(n1191), .B(n1454), .CI(n1177), .CO(n1174), .S(n1175) );
  HA_X1 U796 ( .A(n1432), .B(n1477), .CO(n1176), .S(n1177) );
  FA_X1 U797 ( .A(n1455), .B(n1478), .CI(n1180), .CO(n1178), .S(n1179) );
  HA_X1 U798 ( .A(n1456), .B(n1479), .CO(n1180), .S(n1181) );
  XNOR2_X1 U1448 ( .A(n551), .B(n1929), .ZN(product[23]) );
  AND2_X1 U1449 ( .A1(n2093), .A2(n550), .ZN(n1929) );
  XNOR2_X1 U1450 ( .A(n544), .B(n1930), .ZN(product[24]) );
  AND2_X1 U1451 ( .A1(n2214), .A2(n543), .ZN(n1930) );
  INV_X1 U1452 ( .A(n2216), .ZN(n1931) );
  CLKBUF_X1 U1453 ( .A(n2197), .Z(n1932) );
  INV_X2 U1454 ( .A(n1932), .ZN(n2265) );
  CLKBUF_X1 U1455 ( .A(a[15]), .Z(n2175) );
  NOR2_X2 U1456 ( .A1(n1933), .A2(n2206), .ZN(n2151) );
  XNOR2_X1 U1457 ( .A(n1936), .B(n2164), .ZN(n1933) );
  OR2_X1 U1458 ( .A1(n2153), .A2(n2147), .ZN(n1955) );
  BUF_X1 U1459 ( .A(n512), .Z(n2105) );
  OR2_X2 U1460 ( .A1(n1983), .A2(n2143), .ZN(n1934) );
  INV_X1 U1461 ( .A(n2286), .ZN(n2283) );
  BUF_X1 U1462 ( .A(n2222), .Z(n1949) );
  CLKBUF_X1 U1463 ( .A(a[3]), .Z(n1935) );
  CLKBUF_X1 U1464 ( .A(a[22]), .Z(n1936) );
  OR2_X2 U1465 ( .A1(n2141), .A2(n2142), .ZN(n1284) );
  CLKBUF_X1 U1466 ( .A(n535), .Z(n1937) );
  XNOR2_X1 U1467 ( .A(a[8]), .B(n2306), .ZN(n1813) );
  XOR2_X1 U1468 ( .A(a[14]), .B(a[13]), .Z(n1938) );
  XOR2_X1 U1469 ( .A(a[14]), .B(a[13]), .Z(n2148) );
  NAND2_X1 U1470 ( .A1(n2220), .A2(n2221), .ZN(n1939) );
  INV_X2 U1471 ( .A(n1974), .ZN(n2247) );
  CLKBUF_X1 U1472 ( .A(n877), .Z(n1940) );
  BUF_X4 U1473 ( .A(n2249), .Z(n2162) );
  INV_X2 U1474 ( .A(n2325), .ZN(n2322) );
  OR2_X2 U1475 ( .A1(n2153), .A2(n2147), .ZN(n1941) );
  INV_X1 U1476 ( .A(n2272), .ZN(n1942) );
  BUF_X1 U1477 ( .A(n836), .Z(n2026) );
  INV_X1 U1478 ( .A(a[13]), .ZN(n1943) );
  INV_X1 U1479 ( .A(n1943), .ZN(n1945) );
  INV_X1 U1480 ( .A(n1943), .ZN(n1944) );
  INV_X1 U1481 ( .A(n1943), .ZN(n2296) );
  BUF_X4 U1482 ( .A(n2045), .Z(n1946) );
  BUF_X1 U1483 ( .A(n1979), .Z(n2020) );
  NAND3_X1 U1484 ( .A1(n2176), .A2(n2177), .A3(n2178), .ZN(n1947) );
  XNOR2_X1 U1485 ( .A(a[16]), .B(n2291), .ZN(n1809) );
  OR2_X2 U1486 ( .A1(n2159), .A2(n2143), .ZN(n1948) );
  INV_X1 U1487 ( .A(n2288), .ZN(n1950) );
  INV_X1 U1488 ( .A(n1950), .ZN(n1951) );
  INV_X1 U1489 ( .A(n1950), .ZN(n1953) );
  INV_X2 U1490 ( .A(n1950), .ZN(n1952) );
  XNOR2_X1 U1491 ( .A(a[10]), .B(n2302), .ZN(n2115) );
  OAI22_X1 U1492 ( .A1(n2247), .A2(n1683), .B1(n1682), .B2(n2268), .ZN(n1954)
         );
  XOR2_X1 U1493 ( .A(b[5]), .B(n2292), .Z(n1575) );
  INV_X1 U1494 ( .A(n2291), .ZN(n2288) );
  OAI22_X1 U1495 ( .A1(n2248), .A2(n1719), .B1(n2270), .B2(n1718), .ZN(n1421)
         );
  BUF_X2 U1496 ( .A(n1963), .Z(n2028) );
  INV_X1 U1497 ( .A(n2077), .ZN(n2216) );
  INV_X1 U1498 ( .A(n2145), .ZN(n2246) );
  XOR2_X1 U1499 ( .A(n2098), .B(n2202), .Z(n1043) );
  NAND3_X1 U1500 ( .A1(n2081), .A2(n2082), .A3(n2083), .ZN(n882) );
  NOR2_X1 U1501 ( .A1(n789), .A2(n804), .ZN(n480) );
  AND2_X1 U1502 ( .A1(n1193), .A2(n1481), .ZN(n1956) );
  AND2_X1 U1503 ( .A1(n1039), .A2(n1054), .ZN(n1957) );
  OR2_X1 U1504 ( .A1(n1457), .A2(n1480), .ZN(n1958) );
  OR2_X1 U1505 ( .A1(n1179), .A2(n1433), .ZN(n1959) );
  AND2_X1 U1506 ( .A1(n1143), .A2(n1150), .ZN(n1960) );
  AND2_X1 U1507 ( .A1(n1123), .A2(n1132), .ZN(n1961) );
  AND2_X1 U1508 ( .A1(n1151), .A2(n1158), .ZN(n1962) );
  OR2_X1 U1509 ( .A1(n2150), .A2(n1938), .ZN(n1963) );
  AND2_X1 U1510 ( .A1(n1457), .A2(n1480), .ZN(n1964) );
  AND2_X1 U1511 ( .A1(n1179), .A2(n1433), .ZN(n1965) );
  AND2_X1 U1512 ( .A1(n1133), .A2(n1142), .ZN(n1966) );
  AND2_X1 U1513 ( .A1(n1111), .A2(n1122), .ZN(n1967) );
  AND2_X1 U1514 ( .A1(n1055), .A2(n1070), .ZN(n1968) );
  AND2_X1 U1515 ( .A1(n1021), .A2(n1038), .ZN(n1969) );
  OR2_X1 U1516 ( .A1(n1151), .A2(n1158), .ZN(n1970) );
  OR2_X1 U1517 ( .A1(n1143), .A2(n1150), .ZN(n1971) );
  XNOR2_X1 U1518 ( .A(n560), .B(n1972), .ZN(product[22]) );
  AND2_X1 U1519 ( .A1(n2182), .A2(n559), .ZN(n1972) );
  XNOR2_X1 U1520 ( .A(n1949), .B(n1973), .ZN(product[34]) );
  AND2_X1 U1521 ( .A1(n663), .A2(n439), .ZN(n1973) );
  NOR2_X1 U1522 ( .A1(n2153), .A2(n2147), .ZN(n1974) );
  BUF_X1 U1523 ( .A(n536), .Z(n1976) );
  CLKBUF_X2 U1524 ( .A(n2013), .Z(n1988) );
  BUF_X2 U1525 ( .A(n2013), .Z(n1987) );
  CLKBUF_X1 U1526 ( .A(n552), .Z(n1975) );
  BUF_X1 U1527 ( .A(n505), .Z(n2196) );
  BUF_X1 U1528 ( .A(n536), .Z(n1978) );
  BUF_X1 U1529 ( .A(n536), .Z(n1977) );
  INV_X2 U1530 ( .A(n2010), .ZN(n2255) );
  XOR2_X1 U1531 ( .A(a[18]), .B(n2292), .Z(n1979) );
  XNOR2_X1 U1532 ( .A(a[0]), .B(n2324), .ZN(n1817) );
  INV_X1 U1533 ( .A(n2144), .ZN(n1981) );
  INV_X1 U1534 ( .A(n2144), .ZN(n1980) );
  INV_X1 U1535 ( .A(n2144), .ZN(n2252) );
  INV_X1 U1536 ( .A(n2284), .ZN(n1982) );
  INV_X2 U1537 ( .A(n2287), .ZN(n2284) );
  XOR2_X1 U1538 ( .A(a[18]), .B(n2286), .Z(n1983) );
  CLKBUF_X1 U1539 ( .A(n2273), .Z(n1985) );
  CLKBUF_X3 U1540 ( .A(n2273), .Z(n1984) );
  BUF_X1 U1541 ( .A(n251), .Z(n2273) );
  INV_X1 U1542 ( .A(n1987), .ZN(n1986) );
  BUF_X2 U1543 ( .A(n2239), .Z(n2168) );
  INV_X1 U1544 ( .A(n2276), .ZN(n1990) );
  INV_X1 U1545 ( .A(n2276), .ZN(n1989) );
  CLKBUF_X1 U1546 ( .A(n2258), .Z(n1991) );
  CLKBUF_X3 U1547 ( .A(n2258), .Z(n1992) );
  INV_X1 U1548 ( .A(n2260), .ZN(n2258) );
  INV_X2 U1549 ( .A(n2311), .ZN(n1994) );
  INV_X2 U1550 ( .A(n2311), .ZN(n1993) );
  INV_X1 U1551 ( .A(n2020), .ZN(n1995) );
  XNOR2_X1 U1552 ( .A(a[18]), .B(n2292), .ZN(n2143) );
  BUF_X1 U1553 ( .A(n1963), .Z(n2027) );
  BUF_X2 U1554 ( .A(n2297), .Z(n2029) );
  OAI22_X1 U1555 ( .A1(n2245), .A2(n1658), .B1(n1657), .B2(n2266), .ZN(n1996)
         );
  OR2_X2 U1556 ( .A1(n2160), .A2(n2157), .ZN(n1997) );
  INV_X1 U1557 ( .A(n2223), .ZN(n1998) );
  INV_X1 U1558 ( .A(n1955), .ZN(n1999) );
  INV_X1 U1559 ( .A(n2015), .ZN(n2157) );
  BUF_X1 U1560 ( .A(n1462), .Z(n2000) );
  INV_X1 U1561 ( .A(n2307), .ZN(n2002) );
  INV_X1 U1562 ( .A(n2307), .ZN(n2001) );
  OR2_X1 U1563 ( .A1(n2150), .A2(n2148), .ZN(n2013) );
  BUF_X1 U1564 ( .A(n1395), .Z(n2019) );
  XNOR2_X1 U1565 ( .A(n818), .B(n2003), .ZN(n797) );
  XNOR2_X1 U1566 ( .A(n1296), .B(n1274), .ZN(n2003) );
  INV_X1 U1567 ( .A(n2145), .ZN(n2245) );
  INV_X1 U1568 ( .A(n1934), .ZN(n2004) );
  INV_X1 U1569 ( .A(n2045), .ZN(n2201) );
  AND2_X1 U1570 ( .A1(n2045), .A2(n1807), .ZN(n2154) );
  INV_X1 U1571 ( .A(n2179), .ZN(n2005) );
  AND2_X2 U1572 ( .A1(n1809), .A2(n2257), .ZN(n2179) );
  FA_X1 U1573 ( .A(n776), .B(n765), .CI(n763), .S(n2006) );
  INV_X1 U1574 ( .A(n2089), .ZN(n2007) );
  OR2_X2 U1575 ( .A1(n2160), .A2(n2157), .ZN(n2022) );
  CLKBUF_X3 U1576 ( .A(n2175), .Z(n2008) );
  NOR2_X1 U1577 ( .A1(n520), .A2(n2007), .ZN(n2009) );
  CLKBUF_X1 U1578 ( .A(n2206), .Z(n2010) );
  CLKBUF_X1 U1579 ( .A(n525), .Z(n2011) );
  INV_X2 U1580 ( .A(n2307), .ZN(n2304) );
  INV_X1 U1581 ( .A(n2095), .ZN(n2012) );
  INV_X2 U1582 ( .A(n2295), .ZN(n2014) );
  XOR2_X1 U1583 ( .A(a[12]), .B(n2298), .Z(n2160) );
  XNOR2_X1 U1584 ( .A(a[12]), .B(a[11]), .ZN(n2015) );
  BUF_X4 U1585 ( .A(n2015), .Z(n2023) );
  CLKBUF_X3 U1586 ( .A(b[0]), .Z(n2016) );
  XNOR2_X1 U1587 ( .A(a[20]), .B(n2281), .ZN(n1807) );
  INV_X1 U1588 ( .A(n2316), .ZN(n2017) );
  INV_X1 U1589 ( .A(n672), .ZN(n2018) );
  BUF_X2 U1590 ( .A(n1979), .Z(n2021) );
  INV_X1 U1591 ( .A(n2303), .ZN(n2025) );
  INV_X1 U1592 ( .A(n2303), .ZN(n2024) );
  BUF_X1 U1593 ( .A(n2297), .Z(n2031) );
  CLKBUF_X3 U1594 ( .A(n2297), .Z(n2030) );
  NOR2_X1 U1595 ( .A1(n805), .A2(n820), .ZN(n2032) );
  NOR2_X1 U1596 ( .A1(n805), .A2(n820), .ZN(n495) );
  OR2_X1 U1597 ( .A1(n534), .A2(n531), .ZN(n2033) );
  NOR2_X1 U1598 ( .A1(n896), .A2(n877), .ZN(n2034) );
  INV_X2 U1599 ( .A(n2145), .ZN(n2036) );
  INV_X2 U1600 ( .A(n2145), .ZN(n2035) );
  INV_X1 U1601 ( .A(n2266), .ZN(n2037) );
  NOR2_X1 U1602 ( .A1(n839), .A2(n856), .ZN(n2038) );
  INV_X1 U1603 ( .A(n2022), .ZN(n2039) );
  OAI21_X1 U1604 ( .B1(n2034), .B2(n535), .A(n532), .ZN(n2040) );
  CLKBUF_X1 U1605 ( .A(n1997), .Z(n2041) );
  OR2_X1 U1606 ( .A1(n456), .A2(n481), .ZN(n2042) );
  NAND2_X1 U1607 ( .A1(n2042), .A2(n457), .ZN(n455) );
  OR2_X1 U1608 ( .A1(n2006), .A2(n774), .ZN(n2043) );
  XOR2_X1 U1609 ( .A(a[6]), .B(a[5]), .Z(n2044) );
  BUF_X2 U1610 ( .A(n2047), .Z(n2167) );
  NOR2_X2 U1611 ( .A1(n727), .A2(n736), .ZN(n428) );
  XNOR2_X1 U1612 ( .A(a[19]), .B(a[20]), .ZN(n2045) );
  BUF_X1 U1613 ( .A(n2239), .Z(n2166) );
  XNOR2_X1 U1614 ( .A(n880), .B(n2046), .ZN(n859) );
  XNOR2_X1 U1615 ( .A(n863), .B(n882), .ZN(n2046) );
  INV_X2 U1616 ( .A(n2280), .ZN(n2277) );
  INV_X2 U1617 ( .A(n2321), .ZN(n2318) );
  INV_X1 U1618 ( .A(n2151), .ZN(n2048) );
  INV_X1 U1619 ( .A(n2151), .ZN(n2047) );
  OR2_X1 U1620 ( .A1(n2238), .A2(n1499), .ZN(n2049) );
  OR2_X1 U1621 ( .A1(n1498), .A2(n2254), .ZN(n2050) );
  NAND2_X1 U1622 ( .A1(n2049), .A2(n2050), .ZN(n1210) );
  NAND2_X2 U1623 ( .A1(n1809), .A2(n2257), .ZN(n2138) );
  XOR2_X1 U1624 ( .A(a[7]), .B(a[8]), .Z(n2197) );
  NAND3_X1 U1625 ( .A1(n2086), .A2(n2087), .A3(n2088), .ZN(n2051) );
  XOR2_X1 U1626 ( .A(n1399), .B(n1421), .Z(n2052) );
  XOR2_X1 U1627 ( .A(n1096), .B(n2052), .Z(n1079) );
  NAND2_X1 U1628 ( .A1(n1096), .A2(n1399), .ZN(n2053) );
  NAND2_X1 U1629 ( .A1(n1096), .A2(n1421), .ZN(n2054) );
  NAND2_X1 U1630 ( .A1(n1399), .A2(n1421), .ZN(n2055) );
  NAND3_X1 U1631 ( .A1(n2053), .A2(n2054), .A3(n2055), .ZN(n1078) );
  XOR2_X1 U1632 ( .A(a[3]), .B(a[4]), .Z(n2158) );
  NAND2_X1 U1633 ( .A1(n2056), .A2(n2057), .ZN(n1306) );
  OR2_X1 U1634 ( .A1(n1988), .A2(n1599), .ZN(n2056) );
  OR2_X1 U1635 ( .A1(n1598), .A2(n2261), .ZN(n2057) );
  INV_X1 U1636 ( .A(n2324), .ZN(n2059) );
  INV_X1 U1637 ( .A(n2324), .ZN(n2058) );
  INV_X1 U1638 ( .A(n2144), .ZN(n2061) );
  INV_X1 U1639 ( .A(n2144), .ZN(n2060) );
  INV_X2 U1640 ( .A(n2311), .ZN(n2309) );
  CLKBUF_X3 U1641 ( .A(a[23]), .Z(n2165) );
  XOR2_X1 U1642 ( .A(n887), .B(n904), .Z(n2062) );
  XOR2_X1 U1643 ( .A(n902), .B(n2062), .Z(n881) );
  NAND2_X1 U1644 ( .A1(n902), .A2(n887), .ZN(n2063) );
  NAND2_X1 U1645 ( .A1(n902), .A2(n904), .ZN(n2064) );
  NAND2_X1 U1646 ( .A1(n887), .A2(n904), .ZN(n2065) );
  NAND3_X1 U1647 ( .A1(n2063), .A2(n2064), .A3(n2065), .ZN(n880) );
  CLKBUF_X1 U1648 ( .A(n473), .Z(n2066) );
  XNOR2_X1 U1649 ( .A(n2067), .B(n1183), .ZN(n999) );
  XNOR2_X1 U1650 ( .A(n1461), .B(n1350), .ZN(n2067) );
  INV_X1 U1651 ( .A(n2295), .ZN(n2294) );
  INV_X1 U1652 ( .A(n2144), .ZN(n2253) );
  INV_X1 U1653 ( .A(n2151), .ZN(n2238) );
  NAND2_X1 U1654 ( .A1(n880), .A2(n863), .ZN(n2068) );
  NAND2_X1 U1655 ( .A1(n880), .A2(n882), .ZN(n2069) );
  NAND2_X1 U1656 ( .A1(n863), .A2(n882), .ZN(n2070) );
  NAND3_X1 U1657 ( .A1(n2068), .A2(n2069), .A3(n2070), .ZN(n858) );
  XOR2_X1 U1658 ( .A(n1056), .B(n1043), .Z(n2071) );
  XOR2_X1 U1659 ( .A(n1041), .B(n2071), .Z(n1039) );
  NAND2_X1 U1660 ( .A1(n1041), .A2(n1056), .ZN(n2072) );
  NAND2_X1 U1661 ( .A1(n1041), .A2(n1043), .ZN(n2073) );
  NAND2_X1 U1662 ( .A1(n1056), .A2(n1043), .ZN(n2074) );
  NAND3_X1 U1663 ( .A1(n2072), .A2(n2073), .A3(n2074), .ZN(n1038) );
  AOI21_X1 U1664 ( .B1(n581), .B2(n567), .A(n568), .ZN(n2075) );
  NAND3_X1 U1665 ( .A1(n2189), .A2(n2190), .A3(n2191), .ZN(n2076) );
  XNOR2_X1 U1666 ( .A(a[9]), .B(a[10]), .ZN(n2077) );
  INV_X2 U1667 ( .A(n2216), .ZN(n2263) );
  BUF_X1 U1668 ( .A(n489), .Z(n2078) );
  CLKBUF_X1 U1669 ( .A(n490), .Z(n2079) );
  XOR2_X1 U1670 ( .A(n893), .B(n889), .Z(n2080) );
  XOR2_X1 U1671 ( .A(n906), .B(n2080), .Z(n883) );
  NAND2_X1 U1672 ( .A1(n906), .A2(n893), .ZN(n2081) );
  NAND2_X1 U1673 ( .A1(n906), .A2(n889), .ZN(n2082) );
  NAND2_X1 U1674 ( .A1(n893), .A2(n889), .ZN(n2083) );
  OR2_X1 U1675 ( .A1(n502), .A2(n495), .ZN(n2084) );
  BUF_X4 U1676 ( .A(n277), .Z(n2223) );
  OR2_X2 U1677 ( .A1(n2152), .A2(n2146), .ZN(n277) );
  XOR2_X1 U1678 ( .A(a[18]), .B(n2286), .Z(n2159) );
  AND2_X2 U1679 ( .A1(n1817), .A2(n251), .ZN(n2144) );
  XOR2_X1 U1680 ( .A(n1078), .B(n1080), .Z(n2085) );
  XOR2_X1 U1681 ( .A(n1082), .B(n2085), .Z(n1061) );
  NAND2_X1 U1682 ( .A1(n1082), .A2(n1078), .ZN(n2086) );
  NAND2_X1 U1683 ( .A1(n1080), .A2(n1082), .ZN(n2087) );
  NAND2_X1 U1684 ( .A1(n1078), .A2(n1080), .ZN(n2088) );
  NAND3_X1 U1685 ( .A1(n2086), .A2(n2087), .A3(n2088), .ZN(n1060) );
  OR2_X1 U1686 ( .A1(n839), .A2(n856), .ZN(n2089) );
  CLKBUF_X1 U1687 ( .A(n547), .Z(n2090) );
  NOR2_X1 U1688 ( .A1(n941), .A2(n962), .ZN(n547) );
  INV_X1 U1689 ( .A(n2197), .ZN(n2264) );
  NOR2_X1 U1690 ( .A1(n1003), .A2(n1020), .ZN(n2091) );
  CLKBUF_X1 U1691 ( .A(n521), .Z(n2092) );
  OR2_X1 U1692 ( .A1(n941), .A2(n962), .ZN(n2093) );
  BUF_X1 U1693 ( .A(a[23]), .Z(n2164) );
  INV_X1 U1694 ( .A(n2312), .ZN(n2310) );
  XOR2_X1 U1695 ( .A(a[22]), .B(a[21]), .Z(n2206) );
  INV_X1 U1696 ( .A(n2269), .ZN(n2094) );
  INV_X1 U1697 ( .A(n2094), .ZN(n2095) );
  INV_X1 U1698 ( .A(n2094), .ZN(n2097) );
  INV_X1 U1699 ( .A(n2094), .ZN(n2096) );
  AND2_X2 U1700 ( .A1(n2115), .A2(n2077), .ZN(n2149) );
  INV_X1 U1701 ( .A(n2206), .ZN(n2254) );
  NOR2_X1 U1702 ( .A1(n839), .A2(n856), .ZN(n513) );
  AOI21_X2 U1703 ( .B1(n426), .B2(n445), .A(n427), .ZN(n421) );
  BUF_X1 U1704 ( .A(n2249), .Z(n2161) );
  CLKBUF_X1 U1705 ( .A(n2051), .Z(n2098) );
  XOR2_X1 U1706 ( .A(n895), .B(n891), .Z(n2099) );
  XOR2_X1 U1707 ( .A(n908), .B(n2099), .Z(n885) );
  NAND2_X1 U1708 ( .A1(n908), .A2(n895), .ZN(n2100) );
  NAND2_X1 U1709 ( .A1(n908), .A2(n891), .ZN(n2101) );
  NAND2_X1 U1710 ( .A1(n895), .A2(n891), .ZN(n2102) );
  NAND3_X1 U1711 ( .A1(n2100), .A2(n2101), .A3(n2102), .ZN(n884) );
  XNOR2_X1 U1712 ( .A(n2103), .B(n999), .ZN(n989) );
  XNOR2_X1 U1713 ( .A(n1012), .B(n997), .ZN(n2103) );
  XOR2_X1 U1714 ( .A(n1238), .B(n1216), .Z(n2104) );
  INV_X2 U1715 ( .A(n2149), .ZN(n2244) );
  INV_X2 U1716 ( .A(n2149), .ZN(n2243) );
  NAND2_X1 U1717 ( .A1(n1461), .A2(n1350), .ZN(n2106) );
  NAND2_X1 U1718 ( .A1(n1461), .A2(n1183), .ZN(n2107) );
  NAND2_X1 U1719 ( .A1(n1350), .A2(n1183), .ZN(n2108) );
  NAND3_X1 U1720 ( .A1(n2106), .A2(n2107), .A3(n2108), .ZN(n998) );
  NAND2_X1 U1721 ( .A1(n1012), .A2(n997), .ZN(n2109) );
  NAND2_X1 U1722 ( .A1(n997), .A2(n999), .ZN(n2110) );
  NAND2_X1 U1723 ( .A1(n1012), .A2(n999), .ZN(n2111) );
  NAND3_X1 U1724 ( .A1(n2109), .A2(n2110), .A3(n2111), .ZN(n988) );
  OR2_X1 U1725 ( .A1(n2169), .A2(n2280), .ZN(n2112) );
  OR2_X1 U1726 ( .A1(n1531), .A2(n1946), .ZN(n2113) );
  NAND2_X1 U1727 ( .A1(n2112), .A2(n2113), .ZN(n1183) );
  BUF_X2 U1728 ( .A(n2241), .Z(n2170) );
  AND2_X2 U1729 ( .A1(n1813), .A2(n2264), .ZN(n2145) );
  BUF_X2 U1730 ( .A(n2241), .Z(n2169) );
  AND2_X2 U1731 ( .A1(n2235), .A2(n2236), .ZN(n2222) );
  AND2_X2 U1732 ( .A1(n2235), .A2(n2236), .ZN(n301) );
  INV_X1 U1733 ( .A(n2295), .ZN(n2293) );
  XNOR2_X1 U1734 ( .A(n1031), .B(n2114), .ZN(n1027) );
  XNOR2_X1 U1735 ( .A(n1033), .B(n1048), .ZN(n2114) );
  INV_X2 U1736 ( .A(n2317), .ZN(n2313) );
  INV_X2 U1737 ( .A(b[0]), .ZN(n2326) );
  INV_X1 U1738 ( .A(n2179), .ZN(n2117) );
  INV_X1 U1739 ( .A(n2179), .ZN(n2116) );
  NOR2_X1 U1740 ( .A1(n2084), .A2(n467), .ZN(n465) );
  NAND2_X1 U1741 ( .A1(n663), .A2(n662), .ZN(n431) );
  OAI21_X1 U1742 ( .B1(n492), .B2(n467), .A(n468), .ZN(n466) );
  INV_X1 U1743 ( .A(n481), .ZN(n483) );
  NOR2_X1 U1744 ( .A1(n502), .A2(n2032), .ZN(n489) );
  INV_X1 U1745 ( .A(n435), .ZN(n662) );
  INV_X1 U1746 ( .A(n503), .ZN(n501) );
  INV_X1 U1747 ( .A(n438), .ZN(n663) );
  NAND2_X1 U1748 ( .A1(n666), .A2(n481), .ZN(n315) );
  NAND2_X1 U1749 ( .A1(n667), .A2(n496), .ZN(n316) );
  NAND2_X1 U1750 ( .A1(n668), .A2(n503), .ZN(n317) );
  NAND2_X1 U1751 ( .A1(n2089), .A2(n514), .ZN(n318) );
  NAND2_X1 U1752 ( .A1(n662), .A2(n436), .ZN(n311) );
  NOR2_X1 U1753 ( .A1(n420), .A2(n402), .ZN(n400) );
  NAND2_X1 U1754 ( .A1(n426), .A2(n663), .ZN(n420) );
  AOI21_X1 U1755 ( .B1(n662), .B2(n445), .A(n434), .ZN(n432) );
  INV_X1 U1756 ( .A(n436), .ZN(n434) );
  NOR2_X1 U1757 ( .A1(n402), .A2(n360), .ZN(n356) );
  INV_X1 U1758 ( .A(n564), .ZN(n562) );
  INV_X1 U1759 ( .A(n563), .ZN(n561) );
  INV_X1 U1760 ( .A(n382), .ZN(n380) );
  AOI21_X1 U1761 ( .B1(n2121), .B2(n416), .A(n407), .ZN(n405) );
  INV_X1 U1762 ( .A(n409), .ZN(n407) );
  NOR2_X1 U1763 ( .A1(n435), .A2(n428), .ZN(n426) );
  NOR2_X1 U1764 ( .A1(n597), .A2(n599), .ZN(n595) );
  OAI21_X1 U1765 ( .B1(n620), .B2(n610), .A(n611), .ZN(n609) );
  NOR2_X1 U1766 ( .A1(n384), .A2(n364), .ZN(n362) );
  NAND2_X1 U1767 ( .A1(n661), .A2(n429), .ZN(n310) );
  NOR2_X1 U1768 ( .A1(n983), .A2(n1002), .ZN(n563) );
  NAND2_X1 U1769 ( .A1(n821), .A2(n838), .ZN(n503) );
  NAND2_X1 U1770 ( .A1(n2180), .A2(n532), .ZN(n320) );
  NAND2_X1 U1771 ( .A1(n2121), .A2(n409), .ZN(n308) );
  NAND2_X1 U1772 ( .A1(n422), .A2(n2120), .ZN(n411) );
  NAND2_X1 U1773 ( .A1(n2181), .A2(n378), .ZN(n305) );
  NAND2_X1 U1774 ( .A1(n657), .A2(n387), .ZN(n306) );
  INV_X1 U1775 ( .A(n384), .ZN(n657) );
  NAND2_X1 U1776 ( .A1(n2122), .A2(n396), .ZN(n307) );
  AOI21_X1 U1777 ( .B1(n565), .B2(n561), .A(n562), .ZN(n560) );
  AOI21_X1 U1778 ( .B1(n565), .B2(n545), .A(n546), .ZN(n544) );
  NAND2_X1 U1779 ( .A1(n963), .A2(n982), .ZN(n559) );
  AOI21_X1 U1780 ( .B1(n423), .B2(n2120), .A(n416), .ZN(n412) );
  NAND2_X1 U1781 ( .A1(n789), .A2(n804), .ZN(n481) );
  NOR2_X1 U1782 ( .A1(n389), .A2(n384), .ZN(n382) );
  INV_X1 U1783 ( .A(n378), .ZN(n376) );
  NAND2_X1 U1784 ( .A1(n737), .A2(n748), .ZN(n436) );
  INV_X1 U1785 ( .A(n396), .ZN(n394) );
  NAND2_X1 U1786 ( .A1(n362), .A2(n2122), .ZN(n360) );
  NAND2_X1 U1787 ( .A1(n2120), .A2(n2121), .ZN(n402) );
  OR2_X1 U1788 ( .A1(n1055), .A2(n1070), .ZN(n2118) );
  NAND2_X1 U1789 ( .A1(n1003), .A2(n1020), .ZN(n570) );
  XNOR2_X1 U1790 ( .A(n921), .B(n2119), .ZN(n919) );
  XNOR2_X1 U1791 ( .A(n942), .B(n923), .ZN(n2119) );
  NOR2_X1 U1792 ( .A1(n695), .A2(n700), .ZN(n384) );
  INV_X1 U1793 ( .A(n352), .ZN(n350) );
  AOI21_X1 U1794 ( .B1(n625), .B2(n1970), .A(n1962), .ZN(n620) );
  NOR2_X1 U1795 ( .A1(n1099), .A2(n1110), .ZN(n597) );
  OR2_X1 U1796 ( .A1(n717), .A2(n726), .ZN(n2120) );
  OR2_X1 U1797 ( .A1(n709), .A2(n716), .ZN(n2121) );
  OAI21_X1 U1798 ( .B1(n638), .B2(n636), .A(n637), .ZN(n635) );
  NOR2_X1 U1799 ( .A1(n633), .A2(n631), .ZN(n629) );
  OR2_X1 U1800 ( .A1(n694), .A2(n689), .ZN(n2181) );
  OR2_X1 U1801 ( .A1(n701), .A2(n708), .ZN(n2122) );
  OR2_X1 U1802 ( .A1(n1123), .A2(n1132), .ZN(n2123) );
  AOI21_X1 U1803 ( .B1(n2125), .B2(n1960), .A(n1966), .ZN(n611) );
  XNOR2_X1 U1804 ( .A(n842), .B(n2124), .ZN(n823) );
  XNOR2_X1 U1805 ( .A(n827), .B(n844), .ZN(n2124) );
  AOI21_X1 U1806 ( .B1(n2127), .B2(n1961), .A(n1967), .ZN(n600) );
  OR2_X1 U1807 ( .A1(n1133), .A2(n1142), .ZN(n2125) );
  NAND2_X1 U1808 ( .A1(n2129), .A2(n369), .ZN(n304) );
  NAND2_X1 U1809 ( .A1(n2135), .A2(n341), .ZN(n302) );
  NAND2_X1 U1810 ( .A1(n2134), .A2(n352), .ZN(n303) );
  OR2_X1 U1811 ( .A1(n1021), .A2(n1038), .ZN(n2126) );
  NAND2_X1 U1812 ( .A1(n695), .A2(n700), .ZN(n387) );
  OAI21_X1 U1813 ( .B1(n405), .B2(n360), .A(n361), .ZN(n359) );
  AOI21_X1 U1814 ( .B1(n362), .B2(n394), .A(n363), .ZN(n361) );
  OAI21_X1 U1815 ( .B1(n364), .B2(n387), .A(n365), .ZN(n363) );
  AOI21_X1 U1816 ( .B1(n376), .B2(n2129), .A(n367), .ZN(n365) );
  OR2_X1 U1817 ( .A1(n1111), .A2(n1122), .ZN(n2127) );
  NAND2_X1 U1818 ( .A1(n701), .A2(n708), .ZN(n396) );
  NAND2_X1 U1819 ( .A1(n2181), .A2(n2129), .ZN(n364) );
  INV_X1 U1820 ( .A(n369), .ZN(n367) );
  NAND2_X1 U1821 ( .A1(n1971), .A2(n2125), .ZN(n610) );
  OR2_X1 U1822 ( .A1(n1039), .A2(n1054), .ZN(n2128) );
  INV_X1 U1823 ( .A(n2179), .ZN(n2242) );
  NOR2_X1 U1824 ( .A1(n1165), .A2(n1170), .ZN(n631) );
  OR2_X1 U1825 ( .A1(n685), .A2(n688), .ZN(n2129) );
  BUF_X1 U1826 ( .A(n2077), .Z(n2163) );
  NAND2_X1 U1827 ( .A1(n678), .A2(n677), .ZN(n335) );
  INV_X1 U1828 ( .A(n341), .ZN(n339) );
  AOI21_X1 U1829 ( .B1(n1958), .B2(n1956), .A(n1964), .ZN(n646) );
  AOI21_X1 U1830 ( .B1(n643), .B2(n1959), .A(n1965), .ZN(n638) );
  OAI21_X1 U1831 ( .B1(n646), .B2(n644), .A(n645), .ZN(n643) );
  XNOR2_X1 U1832 ( .A(n994), .B(n2130), .ZN(n973) );
  XNOR2_X1 U1833 ( .A(n1947), .B(n1217), .ZN(n2130) );
  XNOR2_X1 U1834 ( .A(n2104), .B(n2131), .ZN(n953) );
  XNOR2_X1 U1835 ( .A(n1326), .B(n1392), .ZN(n2131) );
  XNOR2_X1 U1836 ( .A(n1284), .B(n2132), .ZN(n997) );
  XNOR2_X1 U1837 ( .A(n1372), .B(n1438), .ZN(n2132) );
  XNOR2_X1 U1838 ( .A(n1417), .B(n2133), .ZN(n1015) );
  XNOR2_X1 U1839 ( .A(n1395), .B(n1462), .ZN(n2133) );
  OR2_X1 U1840 ( .A1(n681), .A2(n684), .ZN(n2134) );
  OR2_X1 U1841 ( .A1(n679), .A2(n680), .ZN(n2135) );
  NAND2_X1 U1842 ( .A1(n681), .A2(n684), .ZN(n352) );
  NAND2_X1 U1843 ( .A1(n679), .A2(n680), .ZN(n341) );
  INV_X1 U1844 ( .A(n676), .ZN(n677) );
  NOR2_X1 U1845 ( .A1(n678), .A2(n677), .ZN(n334) );
  OR2_X1 U1846 ( .A1(n1194), .A2(n676), .ZN(n2136) );
  AND2_X1 U1847 ( .A1(n1194), .A2(n676), .ZN(n2137) );
  INV_X1 U1848 ( .A(n2303), .ZN(n2299) );
  INV_X1 U1849 ( .A(n2281), .ZN(n2278) );
  INV_X1 U1850 ( .A(n2321), .ZN(n2319) );
  INV_X1 U1851 ( .A(n2317), .ZN(n2314) );
  INV_X1 U1852 ( .A(n2148), .ZN(n2261) );
  INV_X1 U1853 ( .A(n2303), .ZN(n2300) );
  INV_X1 U1854 ( .A(n2291), .ZN(n2289) );
  INV_X1 U1855 ( .A(n2276), .ZN(n2275) );
  OAI22_X1 U1856 ( .A1(n2247), .A2(n1683), .B1(n1682), .B2(n2268), .ZN(n836)
         );
  INV_X1 U1857 ( .A(n2044), .ZN(n2268) );
  INV_X1 U1858 ( .A(n1507), .ZN(n2337) );
  INV_X1 U1859 ( .A(n682), .ZN(n683) );
  INV_X1 U1860 ( .A(n2146), .ZN(n2272) );
  INV_X1 U1861 ( .A(n2143), .ZN(n2256) );
  INV_X1 U1862 ( .A(n2311), .ZN(n2308) );
  INV_X1 U1863 ( .A(n2260), .ZN(n2259) );
  OR2_X1 U1864 ( .A1(n2139), .A2(n2140), .ZN(n1417) );
  NOR2_X1 U1865 ( .A1(n2161), .A2(n1715), .ZN(n2139) );
  NOR2_X1 U1866 ( .A1(n2097), .A2(n1714), .ZN(n2140) );
  NOR2_X1 U1867 ( .A1(n2138), .A2(n1576), .ZN(n2141) );
  NOR2_X1 U1868 ( .A1(n1575), .A2(n1991), .ZN(n2142) );
  INV_X1 U1869 ( .A(n724), .ZN(n725) );
  INV_X1 U1870 ( .A(n1632), .ZN(n2332) );
  OAI22_X1 U1871 ( .A1(n2028), .A2(n1586), .B1(n2261), .B2(n1585), .ZN(n1293)
         );
  INV_X1 U1872 ( .A(n1532), .ZN(n2336) );
  OAI22_X1 U1873 ( .A1(n2028), .A2(n1584), .B1(n2261), .B2(n1583), .ZN(n1291)
         );
  INV_X1 U1874 ( .A(n1682), .ZN(n2330) );
  INV_X1 U1875 ( .A(n692), .ZN(n693) );
  OAI21_X1 U1876 ( .B1(n2145), .B2(n2037), .A(n2331), .ZN(n1362) );
  OAI22_X1 U1877 ( .A1(n2028), .A2(n1588), .B1(n2261), .B2(n1587), .ZN(n1295)
         );
  OAI22_X1 U1878 ( .A1(n2028), .A2(n1592), .B1(n2261), .B2(n1591), .ZN(n1299)
         );
  OAI22_X1 U1879 ( .A1(n2028), .A2(n1590), .B1(n2261), .B2(n1589), .ZN(n1297)
         );
  INV_X1 U1880 ( .A(n1707), .ZN(n2329) );
  INV_X1 U1881 ( .A(n1557), .ZN(n2335) );
  INV_X1 U1882 ( .A(n1607), .ZN(n2333) );
  INV_X1 U1883 ( .A(n1657), .ZN(n2331) );
  CLKBUF_X1 U1884 ( .A(n251), .Z(n2274) );
  INV_X1 U1885 ( .A(n1582), .ZN(n2334) );
  INV_X1 U1886 ( .A(n1732), .ZN(n2328) );
  INV_X1 U1887 ( .A(n1482), .ZN(n2338) );
  XNOR2_X1 U1888 ( .A(n2320), .B(b[22]), .ZN(n1733) );
  XNOR2_X1 U1889 ( .A(n2310), .B(b[22]), .ZN(n1683) );
  XNOR2_X1 U1890 ( .A(n2008), .B(b[20]), .ZN(n1585) );
  XNOR2_X1 U1891 ( .A(n2008), .B(b[22]), .ZN(n1583) );
  XNOR2_X1 U1892 ( .A(n2008), .B(b[18]), .ZN(n1587) );
  XNOR2_X1 U1893 ( .A(n2008), .B(b[16]), .ZN(n1589) );
  XNOR2_X1 U1894 ( .A(n2322), .B(b[18]), .ZN(n1762) );
  XNOR2_X1 U1895 ( .A(n2322), .B(b[10]), .ZN(n1770) );
  XNOR2_X1 U1896 ( .A(n2323), .B(b[20]), .ZN(n1760) );
  XNOR2_X1 U1897 ( .A(n2323), .B(b[22]), .ZN(n1758) );
  XNOR2_X1 U1898 ( .A(n2322), .B(b[12]), .ZN(n1768) );
  XNOR2_X1 U1899 ( .A(n2322), .B(b[2]), .ZN(n1778) );
  XNOR2_X1 U1900 ( .A(n2309), .B(b[12]), .ZN(n1693) );
  XNOR2_X1 U1901 ( .A(n1993), .B(b[2]), .ZN(n1703) );
  XNOR2_X1 U1902 ( .A(n2024), .B(b[10]), .ZN(n1645) );
  XNOR2_X1 U1903 ( .A(n2031), .B(b[2]), .ZN(n1628) );
  XNOR2_X1 U1904 ( .A(n2284), .B(b[2]), .ZN(n1553) );
  XNOR2_X1 U1905 ( .A(n2313), .B(b[18]), .ZN(n1712) );
  XNOR2_X1 U1906 ( .A(n2319), .B(b[12]), .ZN(n1743) );
  XNOR2_X1 U1907 ( .A(n2165), .B(b[2]), .ZN(n1503) );
  XNOR2_X1 U1908 ( .A(n1993), .B(b[10]), .ZN(n1695) );
  XNOR2_X1 U1909 ( .A(n2319), .B(b[18]), .ZN(n1737) );
  XNOR2_X1 U1910 ( .A(n2304), .B(b[12]), .ZN(n1668) );
  XNOR2_X1 U1911 ( .A(n2290), .B(b[12]), .ZN(n1568) );
  XNOR2_X1 U1912 ( .A(n2030), .B(b[22]), .ZN(n1608) );
  XNOR2_X1 U1913 ( .A(n2300), .B(b[12]), .ZN(n1643) );
  XNOR2_X1 U1914 ( .A(n2315), .B(b[22]), .ZN(n1708) );
  XNOR2_X1 U1915 ( .A(n2008), .B(b[2]), .ZN(n1603) );
  XNOR2_X1 U1916 ( .A(n2008), .B(b[10]), .ZN(n1595) );
  XNOR2_X1 U1917 ( .A(n2305), .B(b[18]), .ZN(n1662) );
  XNOR2_X1 U1918 ( .A(n2008), .B(b[12]), .ZN(n1593) );
  XNOR2_X1 U1919 ( .A(n2308), .B(b[18]), .ZN(n1687) );
  XNOR2_X1 U1920 ( .A(n2315), .B(b[20]), .ZN(n1710) );
  XNOR2_X1 U1921 ( .A(n1945), .B(b[12]), .ZN(n1618) );
  XNOR2_X1 U1922 ( .A(n2289), .B(b[2]), .ZN(n1578) );
  XNOR2_X1 U1923 ( .A(n2278), .B(b[2]), .ZN(n1528) );
  XNOR2_X1 U1924 ( .A(n2284), .B(b[10]), .ZN(n1545) );
  XNOR2_X1 U1925 ( .A(n2320), .B(b[20]), .ZN(n1735) );
  XNOR2_X1 U1926 ( .A(n2025), .B(b[18]), .ZN(n1637) );
  XNOR2_X1 U1927 ( .A(n2289), .B(b[22]), .ZN(n1558) );
  XNOR2_X1 U1928 ( .A(n2025), .B(b[22]), .ZN(n1633) );
  XNOR2_X1 U1929 ( .A(n2305), .B(b[22]), .ZN(n1658) );
  XNOR2_X1 U1930 ( .A(n2031), .B(b[10]), .ZN(n1620) );
  XNOR2_X1 U1931 ( .A(n2284), .B(b[18]), .ZN(n1537) );
  XNOR2_X1 U1932 ( .A(n2314), .B(b[12]), .ZN(n1718) );
  XNOR2_X1 U1933 ( .A(n2304), .B(b[2]), .ZN(n1678) );
  XNOR2_X1 U1934 ( .A(n2289), .B(b[10]), .ZN(n1570) );
  XNOR2_X1 U1935 ( .A(n2025), .B(b[2]), .ZN(n1653) );
  XNOR2_X1 U1936 ( .A(n2001), .B(b[10]), .ZN(n1670) );
  XNOR2_X1 U1937 ( .A(n2278), .B(b[18]), .ZN(n1512) );
  XNOR2_X1 U1938 ( .A(n2165), .B(b[12]), .ZN(n1493) );
  XNOR2_X1 U1939 ( .A(n2030), .B(b[20]), .ZN(n1610) );
  XNOR2_X1 U1940 ( .A(n2165), .B(b[10]), .ZN(n1495) );
  XNOR2_X1 U1941 ( .A(n2308), .B(b[20]), .ZN(n1685) );
  XNOR2_X1 U1942 ( .A(n2319), .B(b[10]), .ZN(n1745) );
  XNOR2_X1 U1943 ( .A(n2290), .B(b[18]), .ZN(n1562) );
  XNOR2_X1 U1944 ( .A(n2002), .B(b[20]), .ZN(n1660) );
  XNOR2_X1 U1945 ( .A(n2285), .B(b[22]), .ZN(n1533) );
  XNOR2_X1 U1946 ( .A(n2030), .B(b[18]), .ZN(n1612) );
  XNOR2_X1 U1947 ( .A(n2284), .B(b[12]), .ZN(n1543) );
  XNOR2_X1 U1948 ( .A(n2300), .B(b[20]), .ZN(n1635) );
  XNOR2_X1 U1949 ( .A(n2278), .B(b[12]), .ZN(n1518) );
  XNOR2_X1 U1950 ( .A(n2278), .B(b[10]), .ZN(n1520) );
  XNOR2_X1 U1951 ( .A(n2017), .B(b[2]), .ZN(n1728) );
  XNOR2_X1 U1952 ( .A(n2279), .B(b[22]), .ZN(n1508) );
  XNOR2_X1 U1953 ( .A(n2165), .B(b[20]), .ZN(n1485) );
  XNOR2_X1 U1954 ( .A(n2289), .B(b[20]), .ZN(n1560) );
  XNOR2_X1 U1955 ( .A(n2165), .B(b[18]), .ZN(n1487) );
  XNOR2_X1 U1956 ( .A(n2319), .B(b[2]), .ZN(n1753) );
  XNOR2_X1 U1957 ( .A(n2279), .B(b[20]), .ZN(n1510) );
  XNOR2_X1 U1958 ( .A(n2017), .B(b[10]), .ZN(n1720) );
  XNOR2_X1 U1959 ( .A(n2285), .B(b[20]), .ZN(n1535) );
  XNOR2_X1 U1960 ( .A(n2323), .B(b[16]), .ZN(n1764) );
  XNOR2_X1 U1961 ( .A(n2322), .B(b[8]), .ZN(n1772) );
  XNOR2_X1 U1962 ( .A(n2322), .B(b[6]), .ZN(n1774) );
  XNOR2_X1 U1963 ( .A(n2322), .B(b[4]), .ZN(n1776) );
  XNOR2_X1 U1964 ( .A(n2308), .B(b[8]), .ZN(n1697) );
  XNOR2_X1 U1965 ( .A(n2014), .B(b[8]), .ZN(n1597) );
  XNOR2_X1 U1966 ( .A(n2278), .B(b[4]), .ZN(n1526) );
  XNOR2_X1 U1967 ( .A(n2284), .B(b[4]), .ZN(n1551) );
  XNOR2_X1 U1968 ( .A(n2299), .B(b[4]), .ZN(n1651) );
  XNOR2_X1 U1969 ( .A(n2030), .B(b[8]), .ZN(n1622) );
  XNOR2_X1 U1970 ( .A(n2165), .B(b[6]), .ZN(n1499) );
  XNOR2_X1 U1971 ( .A(n2029), .B(b[6]), .ZN(n1624) );
  XNOR2_X1 U1972 ( .A(n2165), .B(b[8]), .ZN(n1497) );
  XNOR2_X1 U1973 ( .A(n2165), .B(b[4]), .ZN(n1501) );
  XNOR2_X1 U1974 ( .A(n1993), .B(b[6]), .ZN(n1699) );
  XNOR2_X1 U1975 ( .A(n2289), .B(b[6]), .ZN(n1574) );
  XNOR2_X1 U1976 ( .A(n2290), .B(b[8]), .ZN(n1572) );
  XNOR2_X1 U1977 ( .A(n2313), .B(b[6]), .ZN(n1724) );
  XNOR2_X1 U1978 ( .A(n2278), .B(b[6]), .ZN(n1524) );
  XNOR2_X1 U1979 ( .A(n2002), .B(b[6]), .ZN(n1674) );
  XNOR2_X1 U1980 ( .A(n2284), .B(b[8]), .ZN(n1547) );
  XNOR2_X1 U1981 ( .A(n2284), .B(b[6]), .ZN(n1549) );
  XNOR2_X1 U1982 ( .A(n2299), .B(b[6]), .ZN(n1649) );
  XNOR2_X1 U1983 ( .A(n2296), .B(b[16]), .ZN(n1614) );
  XNOR2_X1 U1984 ( .A(n2308), .B(b[4]), .ZN(n1701) );
  XNOR2_X1 U1985 ( .A(n1994), .B(b[16]), .ZN(n1689) );
  XNOR2_X1 U1986 ( .A(n2024), .B(b[16]), .ZN(n1639) );
  XNOR2_X1 U1987 ( .A(n2008), .B(b[4]), .ZN(n1601) );
  XNOR2_X1 U1988 ( .A(n1944), .B(b[4]), .ZN(n1626) );
  XNOR2_X1 U1989 ( .A(n2304), .B(b[8]), .ZN(n1672) );
  XNOR2_X1 U1990 ( .A(n2001), .B(b[16]), .ZN(n1664) );
  XNOR2_X1 U1991 ( .A(n2285), .B(b[16]), .ZN(n1539) );
  XNOR2_X1 U1992 ( .A(n2278), .B(b[8]), .ZN(n1522) );
  XNOR2_X1 U1993 ( .A(n2165), .B(b[16]), .ZN(n1489) );
  XNOR2_X1 U1994 ( .A(n2320), .B(b[16]), .ZN(n1739) );
  XNOR2_X1 U1995 ( .A(n2319), .B(b[8]), .ZN(n1747) );
  XNOR2_X1 U1996 ( .A(n2290), .B(b[16]), .ZN(n1564) );
  XNOR2_X1 U1997 ( .A(n2319), .B(b[6]), .ZN(n1749) );
  XNOR2_X1 U1998 ( .A(n2304), .B(b[4]), .ZN(n1676) );
  XNOR2_X1 U1999 ( .A(n2017), .B(b[4]), .ZN(n1726) );
  XNOR2_X1 U2000 ( .A(n2319), .B(b[4]), .ZN(n1751) );
  XNOR2_X1 U2001 ( .A(n2017), .B(b[8]), .ZN(n1722) );
  XNOR2_X1 U2002 ( .A(n2279), .B(b[16]), .ZN(n1514) );
  XNOR2_X1 U2003 ( .A(b[23]), .B(n2318), .ZN(n1732) );
  XNOR2_X1 U2004 ( .A(n1993), .B(b[14]), .ZN(n1691) );
  XNOR2_X1 U2005 ( .A(b[23]), .B(n2313), .ZN(n1707) );
  XNOR2_X1 U2006 ( .A(b[23]), .B(n2300), .ZN(n1632) );
  XNOR2_X1 U2007 ( .A(b[23]), .B(n1953), .ZN(n1557) );
  XNOR2_X1 U2008 ( .A(b[23]), .B(n2277), .ZN(n1507) );
  XNOR2_X1 U2009 ( .A(n2322), .B(b[14]), .ZN(n1766) );
  XNOR2_X1 U2010 ( .A(n2294), .B(b[14]), .ZN(n1591) );
  XNOR2_X1 U2011 ( .A(b[7]), .B(n2313), .ZN(n1723) );
  XNOR2_X1 U2012 ( .A(b[7]), .B(n2275), .ZN(n1498) );
  XNOR2_X1 U2013 ( .A(b[3]), .B(n2275), .ZN(n1502) );
  XNOR2_X1 U2014 ( .A(b[3]), .B(n1951), .ZN(n1577) );
  XNOR2_X1 U2015 ( .A(b[7]), .B(n1951), .ZN(n1573) );
  XNOR2_X1 U2016 ( .A(b[7]), .B(n2300), .ZN(n1648) );
  XNOR2_X1 U2017 ( .A(b[7]), .B(n2318), .ZN(n1748) );
  XNOR2_X1 U2018 ( .A(b[3]), .B(n2318), .ZN(n1752) );
  XNOR2_X1 U2019 ( .A(b[3]), .B(n2301), .ZN(n1652) );
  XNOR2_X1 U2020 ( .A(b[3]), .B(n2314), .ZN(n1727) );
  XOR2_X1 U2021 ( .A(a[2]), .B(a[1]), .Z(n2146) );
  XOR2_X1 U2022 ( .A(a[6]), .B(a[5]), .Z(n2147) );
  XNOR2_X1 U2023 ( .A(b[5]), .B(n2025), .ZN(n1650) );
  XNOR2_X1 U2024 ( .A(b[5]), .B(n1990), .ZN(n1500) );
  XNOR2_X1 U2025 ( .A(b[9]), .B(n1952), .ZN(n1571) );
  XNOR2_X1 U2026 ( .A(b[1]), .B(n1953), .ZN(n1579) );
  XNOR2_X1 U2027 ( .A(b[5]), .B(n2314), .ZN(n1725) );
  XNOR2_X1 U2028 ( .A(b[1]), .B(n2024), .ZN(n1654) );
  XNOR2_X1 U2029 ( .A(b[9]), .B(n2275), .ZN(n1496) );
  XNOR2_X1 U2030 ( .A(b[1]), .B(n2318), .ZN(n1754) );
  XNOR2_X1 U2031 ( .A(b[5]), .B(n2318), .ZN(n1750) );
  XNOR2_X1 U2032 ( .A(b[9]), .B(n2318), .ZN(n1746) );
  XNOR2_X1 U2033 ( .A(b[1]), .B(n2314), .ZN(n1729) );
  XNOR2_X1 U2034 ( .A(b[9]), .B(n2314), .ZN(n1721) );
  XNOR2_X1 U2035 ( .A(a[14]), .B(n2175), .ZN(n2150) );
  XNOR2_X1 U2036 ( .A(b[13]), .B(n1989), .ZN(n1492) );
  XNOR2_X1 U2037 ( .A(b[17]), .B(n1989), .ZN(n1488) );
  XNOR2_X1 U2038 ( .A(b[11]), .B(n1990), .ZN(n1494) );
  XNOR2_X1 U2039 ( .A(b[15]), .B(n1990), .ZN(n1490) );
  XNOR2_X1 U2040 ( .A(b[19]), .B(n2275), .ZN(n1486) );
  XNOR2_X1 U2041 ( .A(b[21]), .B(n1989), .ZN(n1484) );
  XNOR2_X1 U2042 ( .A(n2165), .B(b[14]), .ZN(n1491) );
  XNOR2_X1 U2043 ( .A(n1944), .B(b[14]), .ZN(n1616) );
  XNOR2_X1 U2044 ( .A(n2304), .B(b[14]), .ZN(n1666) );
  XNOR2_X1 U2045 ( .A(n2301), .B(b[14]), .ZN(n1641) );
  XNOR2_X1 U2046 ( .A(n2319), .B(b[14]), .ZN(n1741) );
  XNOR2_X1 U2047 ( .A(n2314), .B(b[14]), .ZN(n1716) );
  XNOR2_X1 U2048 ( .A(n2278), .B(b[14]), .ZN(n1516) );
  XNOR2_X1 U2049 ( .A(n2284), .B(b[14]), .ZN(n1541) );
  XNOR2_X1 U2050 ( .A(n2289), .B(b[14]), .ZN(n1566) );
  XNOR2_X1 U2051 ( .A(a[2]), .B(n1935), .ZN(n2152) );
  XNOR2_X1 U2052 ( .A(a[6]), .B(n2310), .ZN(n2153) );
  NOR2_X1 U2053 ( .A1(n2156), .A2(n2158), .ZN(n2155) );
  XNOR2_X1 U2054 ( .A(a[4]), .B(a[5]), .ZN(n2156) );
  OAI21_X1 U2055 ( .B1(a[0]), .B2(n2144), .A(n2327), .ZN(n1458) );
  INV_X1 U2056 ( .A(n1757), .ZN(n2327) );
  INV_X1 U2057 ( .A(n267), .ZN(n2260) );
  INV_X1 U2058 ( .A(a[23]), .ZN(n2276) );
  INV_X1 U2059 ( .A(a[0]), .ZN(n251) );
  XNOR2_X1 U2060 ( .A(n2165), .B(b[22]), .ZN(n1483) );
  XNOR2_X1 U2061 ( .A(b[23]), .B(n1990), .ZN(n1482) );
  INV_X1 U2062 ( .A(n2155), .ZN(n2249) );
  OAI21_X1 U2063 ( .B1(n2154), .B2(n2201), .A(n2337), .ZN(n1218) );
  INV_X1 U2064 ( .A(n2032), .ZN(n667) );
  INV_X1 U2065 ( .A(n2151), .ZN(n2239) );
  INV_X1 U2066 ( .A(n2154), .ZN(n2241) );
  XOR2_X1 U2067 ( .A(n912), .B(n910), .Z(n2171) );
  XOR2_X1 U2068 ( .A(n914), .B(n2171), .Z(n887) );
  NAND2_X1 U2069 ( .A1(n914), .A2(n912), .ZN(n2172) );
  NAND2_X1 U2070 ( .A1(n914), .A2(n910), .ZN(n2173) );
  NAND2_X1 U2071 ( .A1(n912), .A2(n910), .ZN(n2174) );
  NAND3_X1 U2072 ( .A1(n2172), .A2(n2173), .A3(n2174), .ZN(n886) );
  INV_X1 U2073 ( .A(n520), .ZN(n670) );
  OAI21_X1 U2074 ( .B1(n2151), .B2(n2010), .A(n2338), .ZN(n1194) );
  OAI21_X1 U2075 ( .B1(n2149), .B2(n2216), .A(n2332), .ZN(n1338) );
  NAND2_X1 U2076 ( .A1(n1284), .A2(n1372), .ZN(n2176) );
  NAND2_X1 U2077 ( .A1(n1284), .A2(n1438), .ZN(n2177) );
  NAND2_X1 U2078 ( .A1(n1372), .A2(n1438), .ZN(n2178) );
  NAND3_X1 U2079 ( .A1(n2176), .A2(n2177), .A3(n2178), .ZN(n996) );
  XNOR2_X1 U2080 ( .A(n2289), .B(b[4]), .ZN(n1576) );
  INV_X1 U2081 ( .A(n552), .ZN(n554) );
  OR2_X1 U2082 ( .A1(n896), .A2(n1940), .ZN(n2180) );
  NOR2_X1 U2083 ( .A1(n877), .A2(n896), .ZN(n531) );
  OAI21_X1 U2084 ( .B1(n628), .B2(n626), .A(n627), .ZN(n625) );
  OAI22_X1 U2085 ( .A1(n1981), .A2(n1772), .B1(n1771), .B2(n1985), .ZN(n1473)
         );
  OAI22_X1 U2086 ( .A1(n2060), .A2(n1777), .B1(n1776), .B2(n1984), .ZN(n1478)
         );
  OAI22_X1 U2087 ( .A1(n2061), .A2(n1776), .B1(n1775), .B2(n1985), .ZN(n1477)
         );
  OAI22_X1 U2088 ( .A1(n2061), .A2(n1780), .B1(n1779), .B2(n1985), .ZN(n1481)
         );
  OAI22_X1 U2089 ( .A1(n2252), .A2(n1775), .B1(n1774), .B2(n1984), .ZN(n1476)
         );
  OAI22_X1 U2090 ( .A1(n1981), .A2(n1769), .B1(n1768), .B2(n1984), .ZN(n1470)
         );
  OAI22_X1 U2091 ( .A1(n2061), .A2(n1771), .B1(n1770), .B2(n1984), .ZN(n1472)
         );
  OAI22_X1 U2092 ( .A1(n1980), .A2(n1779), .B1(n1778), .B2(n1984), .ZN(n1480)
         );
  OAI22_X1 U2093 ( .A1(n2060), .A2(n1774), .B1(n1773), .B2(n1985), .ZN(n1475)
         );
  OAI22_X1 U2094 ( .A1(n1981), .A2(n1773), .B1(n1772), .B2(n1985), .ZN(n1474)
         );
  OAI22_X1 U2095 ( .A1(n1980), .A2(n1778), .B1(n1777), .B2(n1984), .ZN(n1479)
         );
  OAI22_X1 U2096 ( .A1(n2061), .A2(n1770), .B1(n1769), .B2(n1984), .ZN(n1471)
         );
  XNOR2_X1 U2097 ( .A(b[23]), .B(n2283), .ZN(n1532) );
  XNOR2_X1 U2098 ( .A(b[7]), .B(n2283), .ZN(n1548) );
  XNOR2_X1 U2099 ( .A(b[9]), .B(n2283), .ZN(n1546) );
  XNOR2_X1 U2100 ( .A(b[3]), .B(n2283), .ZN(n1552) );
  XNOR2_X1 U2101 ( .A(b[1]), .B(n2283), .ZN(n1554) );
  XNOR2_X1 U2102 ( .A(b[5]), .B(n2283), .ZN(n1550) );
  XNOR2_X1 U2103 ( .A(b[7]), .B(n2277), .ZN(n1523) );
  XNOR2_X1 U2104 ( .A(b[5]), .B(n2277), .ZN(n1525) );
  XNOR2_X1 U2105 ( .A(b[3]), .B(n2277), .ZN(n1527) );
  XNOR2_X1 U2106 ( .A(b[1]), .B(n2277), .ZN(n1529) );
  XNOR2_X1 U2107 ( .A(b[9]), .B(n2277), .ZN(n1521) );
  NOR2_X1 U2108 ( .A1(n1085), .A2(n1098), .ZN(n592) );
  NAND2_X1 U2109 ( .A1(n1085), .A2(n1098), .ZN(n593) );
  XNOR2_X1 U2110 ( .A(b[3]), .B(n2001), .ZN(n1677) );
  XNOR2_X1 U2111 ( .A(b[9]), .B(n2002), .ZN(n1671) );
  XNOR2_X1 U2112 ( .A(b[23]), .B(n2305), .ZN(n1657) );
  XNOR2_X1 U2113 ( .A(b[7]), .B(n2304), .ZN(n1673) );
  XNOR2_X1 U2114 ( .A(b[5]), .B(n2002), .ZN(n1675) );
  XNOR2_X1 U2115 ( .A(b[1]), .B(n2001), .ZN(n1679) );
  OR2_X1 U2116 ( .A1(n963), .A2(n982), .ZN(n2182) );
  XOR2_X1 U2117 ( .A(n873), .B(n888), .Z(n2183) );
  XOR2_X1 U2118 ( .A(n886), .B(n2183), .Z(n863) );
  NAND2_X1 U2119 ( .A1(n886), .A2(n873), .ZN(n2184) );
  NAND2_X1 U2120 ( .A1(n886), .A2(n888), .ZN(n2185) );
  NAND2_X1 U2121 ( .A1(n873), .A2(n888), .ZN(n2186) );
  NAND3_X1 U2122 ( .A1(n2184), .A2(n2185), .A3(n2186), .ZN(n862) );
  CLKBUF_X1 U2123 ( .A(n535), .Z(n2187) );
  XOR2_X1 U2124 ( .A(n1416), .B(n1328), .Z(n2188) );
  XOR2_X1 U2125 ( .A(n2188), .B(n1306), .Z(n995) );
  NAND2_X1 U2126 ( .A1(n1306), .A2(n1416), .ZN(n2189) );
  NAND2_X1 U2127 ( .A1(n1306), .A2(n1328), .ZN(n2190) );
  NAND2_X1 U2128 ( .A1(n1416), .A2(n1328), .ZN(n2191) );
  NAND3_X1 U2129 ( .A1(n2189), .A2(n2190), .A3(n2191), .ZN(n994) );
  XNOR2_X1 U2130 ( .A(b[5]), .B(n1945), .ZN(n1625) );
  XNOR2_X1 U2131 ( .A(b[1]), .B(n1945), .ZN(n1629) );
  XNOR2_X1 U2132 ( .A(b[9]), .B(n2029), .ZN(n1621) );
  XNOR2_X1 U2133 ( .A(b[7]), .B(n2029), .ZN(n1623) );
  XNOR2_X1 U2134 ( .A(b[3]), .B(n1945), .ZN(n1627) );
  XNOR2_X1 U2135 ( .A(b[23]), .B(n2031), .ZN(n1607) );
  NOR2_X1 U2136 ( .A1(n558), .A2(n563), .ZN(n552) );
  NOR2_X1 U2137 ( .A1(n963), .A2(n982), .ZN(n558) );
  OAI21_X1 U2138 ( .B1(n2179), .B2(n2260), .A(n2335), .ZN(n1266) );
  NAND2_X1 U2139 ( .A1(n921), .A2(n942), .ZN(n2192) );
  NAND2_X1 U2140 ( .A1(n921), .A2(n923), .ZN(n2193) );
  NAND2_X1 U2141 ( .A1(n942), .A2(n923), .ZN(n2194) );
  NAND3_X1 U2142 ( .A1(n2192), .A2(n2193), .A3(n2194), .ZN(n918) );
  XNOR2_X1 U2143 ( .A(b[3]), .B(n2008), .ZN(n1602) );
  XNOR2_X1 U2144 ( .A(b[23]), .B(n2008), .ZN(n1582) );
  XNOR2_X1 U2145 ( .A(b[5]), .B(n2008), .ZN(n1600) );
  XNOR2_X1 U2146 ( .A(b[9]), .B(n2014), .ZN(n1596) );
  XNOR2_X1 U2147 ( .A(b[1]), .B(n2014), .ZN(n1604) );
  NOR2_X1 U2148 ( .A1(n919), .A2(n940), .ZN(n2195) );
  NAND2_X1 U2149 ( .A1(n670), .A2(n2092), .ZN(n319) );
  INV_X1 U2150 ( .A(n521), .ZN(n519) );
  NAND2_X1 U2151 ( .A1(n857), .A2(n876), .ZN(n521) );
  NOR2_X1 U2152 ( .A1(n2265), .A2(n2326), .ZN(n1385) );
  NOR2_X1 U2153 ( .A1(n2270), .A2(n2326), .ZN(n1433) );
  NOR2_X1 U2154 ( .A1(n1931), .A2(n2326), .ZN(n1361) );
  NOR2_X1 U2155 ( .A1(n1946), .A2(n2326), .ZN(n1241) );
  NOR2_X1 U2156 ( .A1(n2256), .A2(n2326), .ZN(n1265) );
  NOR2_X1 U2157 ( .A1(n2267), .A2(n2326), .ZN(n1409) );
  NOR2_X1 U2158 ( .A1(n2262), .A2(n2326), .ZN(n1313) );
  NOR2_X1 U2159 ( .A1(n2023), .A2(n2326), .ZN(n1337) );
  NOR2_X1 U2160 ( .A1(n2259), .A2(n2326), .ZN(n1289) );
  NAND2_X1 U2161 ( .A1(n2319), .A2(n2326), .ZN(n1756) );
  NAND2_X1 U2162 ( .A1(n2017), .A2(n2326), .ZN(n1731) );
  NOR2_X1 U2163 ( .A1(n2272), .A2(n2326), .ZN(n1457) );
  NAND2_X1 U2164 ( .A1(n2001), .A2(n2326), .ZN(n1681) );
  NAND2_X1 U2165 ( .A1(n2322), .A2(n2326), .ZN(n1781) );
  NAND2_X1 U2166 ( .A1(n2290), .A2(n2326), .ZN(n1581) );
  NAND2_X1 U2167 ( .A1(n1944), .A2(n2326), .ZN(n1631) );
  NAND2_X1 U2168 ( .A1(n2284), .A2(n2326), .ZN(n1556) );
  NAND2_X1 U2169 ( .A1(n1993), .A2(n2326), .ZN(n1706) );
  NAND2_X1 U2170 ( .A1(n2278), .A2(n2326), .ZN(n1531) );
  XNOR2_X1 U2171 ( .A(n2290), .B(n2016), .ZN(n1580) );
  XNOR2_X1 U2172 ( .A(n2315), .B(n2016), .ZN(n1730) );
  XNOR2_X1 U2173 ( .A(n2030), .B(n2016), .ZN(n1630) );
  XNOR2_X1 U2174 ( .A(n1994), .B(n2016), .ZN(n1705) );
  NAND2_X1 U2175 ( .A1(n2024), .A2(n2326), .ZN(n1656) );
  XNOR2_X1 U2176 ( .A(n2025), .B(n2016), .ZN(n1655) );
  XNOR2_X1 U2177 ( .A(n2323), .B(n2016), .ZN(n1780) );
  NAND2_X1 U2178 ( .A1(n2008), .A2(n2326), .ZN(n1606) );
  XNOR2_X1 U2179 ( .A(n2285), .B(n2016), .ZN(n1555) );
  NAND2_X1 U2180 ( .A1(n2165), .A2(n2326), .ZN(n1506) );
  XNOR2_X1 U2181 ( .A(n2002), .B(n2016), .ZN(n1680) );
  XNOR2_X1 U2182 ( .A(n2320), .B(n2016), .ZN(n1755) );
  XNOR2_X1 U2183 ( .A(n2008), .B(n2016), .ZN(n1605) );
  XNOR2_X1 U2184 ( .A(n2279), .B(n2016), .ZN(n1530) );
  OAI22_X1 U2185 ( .A1(n2060), .A2(n2324), .B1(n1781), .B2(n1984), .ZN(n1193)
         );
  OAI22_X1 U2186 ( .A1(n2060), .A2(n1764), .B1(n1763), .B2(n1985), .ZN(n1465)
         );
  OAI22_X1 U2187 ( .A1(n2252), .A2(n1768), .B1(n1767), .B2(n1984), .ZN(n1469)
         );
  OAI22_X1 U2188 ( .A1(n2061), .A2(n1760), .B1(n1759), .B2(n2274), .ZN(n1461)
         );
  OAI22_X1 U2189 ( .A1(n1980), .A2(n1767), .B1(n1766), .B2(n1985), .ZN(n1468)
         );
  OAI22_X1 U2190 ( .A1(n2252), .A2(n1759), .B1(n1758), .B2(n2274), .ZN(n1460)
         );
  OAI22_X1 U2191 ( .A1(n2060), .A2(n1763), .B1(n1762), .B2(n1984), .ZN(n1464)
         );
  OAI22_X1 U2192 ( .A1(n1980), .A2(n1765), .B1(n1764), .B2(n1985), .ZN(n1466)
         );
  OAI22_X1 U2193 ( .A1(n2252), .A2(n1766), .B1(n1765), .B2(n1984), .ZN(n1467)
         );
  OAI22_X1 U2194 ( .A1(n1981), .A2(n1758), .B1(n1757), .B2(n2274), .ZN(n1459)
         );
  OAI22_X1 U2195 ( .A1(n2253), .A2(n1762), .B1(n1761), .B2(n2274), .ZN(n1463)
         );
  XNOR2_X1 U2196 ( .A(b[23]), .B(n2059), .ZN(n1757) );
  NAND2_X1 U2197 ( .A1(n2043), .A2(n461), .ZN(n313) );
  INV_X1 U2198 ( .A(n461), .ZN(n459) );
  OAI22_X1 U2199 ( .A1(n1948), .A2(n1538), .B1(n2256), .B2(n1537), .ZN(n1247)
         );
  NOR2_X1 U2200 ( .A1(n2034), .A2(n534), .ZN(n525) );
  OR2_X1 U2201 ( .A1(n473), .A2(n460), .ZN(n456) );
  XNOR2_X1 U2202 ( .A(b[5]), .B(n2309), .ZN(n1700) );
  XNOR2_X1 U2203 ( .A(b[1]), .B(n2309), .ZN(n1704) );
  XNOR2_X1 U2204 ( .A(b[7]), .B(n1994), .ZN(n1698) );
  XNOR2_X1 U2205 ( .A(b[3]), .B(n1994), .ZN(n1702) );
  XNOR2_X1 U2206 ( .A(b[9]), .B(n2309), .ZN(n1696) );
  XNOR2_X1 U2207 ( .A(b[23]), .B(n2308), .ZN(n1682) );
  OAI22_X1 U2208 ( .A1(n1948), .A2(n1534), .B1(n2256), .B2(n1533), .ZN(n1243)
         );
  OAI22_X1 U2209 ( .A1(n1934), .A2(n1536), .B1(n2021), .B2(n1535), .ZN(n1245)
         );
  OAI22_X1 U2210 ( .A1(n1934), .A2(n1542), .B1(n2256), .B2(n1541), .ZN(n1251)
         );
  OAI22_X1 U2211 ( .A1(n1934), .A2(n1540), .B1(n2021), .B2(n1539), .ZN(n1249)
         );
  NAND2_X1 U2212 ( .A1(n842), .A2(n827), .ZN(n2198) );
  NAND2_X1 U2213 ( .A1(n842), .A2(n844), .ZN(n2199) );
  NAND2_X1 U2214 ( .A1(n827), .A2(n844), .ZN(n2200) );
  NAND3_X1 U2215 ( .A1(n2198), .A2(n2199), .A3(n2200), .ZN(n822) );
  INV_X1 U2216 ( .A(n2286), .ZN(n2282) );
  XOR2_X1 U2217 ( .A(n1053), .B(n1062), .Z(n2202) );
  NAND2_X1 U2218 ( .A1(n2051), .A2(n1053), .ZN(n2203) );
  NAND2_X1 U2219 ( .A1(n1060), .A2(n1062), .ZN(n2204) );
  NAND2_X1 U2220 ( .A1(n1053), .A2(n1062), .ZN(n2205) );
  NAND3_X1 U2221 ( .A1(n2203), .A2(n2204), .A3(n2205), .ZN(n1042) );
  INV_X1 U2222 ( .A(n2158), .ZN(n2269) );
  INV_X1 U2223 ( .A(n2155), .ZN(n2248) );
  NAND2_X1 U2224 ( .A1(n818), .A2(n1296), .ZN(n2207) );
  NAND2_X1 U2225 ( .A1(n818), .A2(n1274), .ZN(n2208) );
  NAND2_X1 U2226 ( .A1(n1296), .A2(n1274), .ZN(n2209) );
  NAND3_X1 U2227 ( .A1(n2207), .A2(n2208), .A3(n2209), .ZN(n796) );
  NAND2_X1 U2228 ( .A1(n2000), .A2(n1417), .ZN(n2210) );
  NAND2_X1 U2229 ( .A1(n1417), .A2(n2019), .ZN(n2211) );
  NAND2_X1 U2230 ( .A1(n2000), .A2(n2019), .ZN(n2212) );
  NAND3_X1 U2231 ( .A1(n2210), .A2(n2211), .A3(n2212), .ZN(n1014) );
  INV_X1 U2232 ( .A(n555), .ZN(n2213) );
  OAI22_X1 U2233 ( .A1(n2253), .A2(n1761), .B1(n1760), .B2(n2274), .ZN(n1462)
         );
  XNOR2_X1 U2234 ( .A(n2315), .B(b[16]), .ZN(n1714) );
  NAND2_X1 U2235 ( .A1(n919), .A2(n940), .ZN(n543) );
  NOR2_X1 U2236 ( .A1(n919), .A2(n940), .ZN(n542) );
  OAI21_X1 U2237 ( .B1(n2039), .B2(n2157), .A(n2333), .ZN(n1314) );
  INV_X1 U2238 ( .A(n874), .ZN(n875) );
  OAI22_X1 U2239 ( .A1(n2170), .A2(n1513), .B1(n1946), .B2(n1512), .ZN(n1223)
         );
  OAI22_X1 U2240 ( .A1(n2169), .A2(n1515), .B1(n1946), .B2(n1514), .ZN(n1225)
         );
  OAI22_X1 U2241 ( .A1(n2170), .A2(n1511), .B1(n1946), .B2(n1510), .ZN(n1221)
         );
  OAI22_X1 U2242 ( .A1(n2169), .A2(n1509), .B1(n1946), .B2(n1508), .ZN(n1219)
         );
  OAI22_X1 U2243 ( .A1(n2169), .A2(n1517), .B1(n1946), .B2(n1516), .ZN(n1227)
         );
  OR2_X1 U2244 ( .A1(n919), .A2(n940), .ZN(n2214) );
  INV_X1 U2245 ( .A(n802), .ZN(n803) );
  AOI21_X1 U2246 ( .B1(n595), .B2(n609), .A(n596), .ZN(n594) );
  NOR2_X1 U2247 ( .A1(n1003), .A2(n1020), .ZN(n569) );
  INV_X1 U2248 ( .A(n2251), .ZN(n2215) );
  INV_X1 U2249 ( .A(n2044), .ZN(n2267) );
  OAI21_X1 U2250 ( .B1(n600), .B2(n597), .A(n598), .ZN(n596) );
  OAI21_X1 U2251 ( .B1(n1999), .B2(n2147), .A(n2330), .ZN(n1386) );
  INV_X1 U2252 ( .A(n2260), .ZN(n2257) );
  NOR2_X1 U2253 ( .A1(n821), .A2(n838), .ZN(n502) );
  NAND2_X1 U2254 ( .A1(n2104), .A2(n1326), .ZN(n2217) );
  NAND2_X1 U2255 ( .A1(n961), .A2(n1392), .ZN(n2218) );
  NAND2_X1 U2256 ( .A1(n1326), .A2(n1392), .ZN(n2219) );
  NAND3_X1 U2257 ( .A1(n2217), .A2(n2218), .A3(n2219), .ZN(n952) );
  OR2_X1 U2258 ( .A1(n2048), .A2(n1505), .ZN(n2220) );
  OR2_X1 U2259 ( .A1(n1504), .A2(n2254), .ZN(n2221) );
  NAND2_X1 U2260 ( .A1(n2220), .A2(n2221), .ZN(n1216) );
  XNOR2_X1 U2261 ( .A(n2165), .B(n2016), .ZN(n1505) );
  XNOR2_X1 U2262 ( .A(b[1]), .B(n1989), .ZN(n1504) );
  OAI21_X1 U2263 ( .B1(n1986), .B2(n1938), .A(n2334), .ZN(n1290) );
  XNOR2_X1 U2264 ( .A(n522), .B(n319), .ZN(product[27]) );
  XNOR2_X1 U2265 ( .A(n515), .B(n318), .ZN(product[28]) );
  XNOR2_X1 U2266 ( .A(n504), .B(n317), .ZN(product[29]) );
  XNOR2_X1 U2267 ( .A(n497), .B(n316), .ZN(product[30]) );
  XNOR2_X1 U2268 ( .A(n486), .B(n315), .ZN(product[31]) );
  XNOR2_X1 U2269 ( .A(n533), .B(n320), .ZN(product[26]) );
  OAI21_X1 U2270 ( .B1(n2155), .B2(n2012), .A(n2329), .ZN(n1410) );
  AOI21_X1 U2271 ( .B1(n359), .B2(n2134), .A(n350), .ZN(n348) );
  AOI21_X1 U2272 ( .B1(n581), .B2(n567), .A(n568), .ZN(n566) );
  INV_X1 U2273 ( .A(n277), .ZN(n2251) );
  OAI21_X1 U2274 ( .B1(n2004), .B2(n1995), .A(n2336), .ZN(n1242) );
  INV_X1 U2275 ( .A(n2066), .ZN(n665) );
  INV_X1 U2276 ( .A(n2251), .ZN(n2250) );
  INV_X1 U2277 ( .A(n2154), .ZN(n2240) );
  NAND2_X1 U2278 ( .A1(n2120), .A2(n418), .ZN(n309) );
  INV_X1 U2279 ( .A(n418), .ZN(n416) );
  NOR2_X1 U2280 ( .A1(n1159), .A2(n1161), .ZN(n626) );
  NAND2_X1 U2281 ( .A1(n1159), .A2(n1161), .ZN(n627) );
  INV_X1 U2282 ( .A(n2196), .ZN(n507) );
  AOI21_X1 U2283 ( .B1(n589), .B2(n2118), .A(n1968), .ZN(n583) );
  NAND2_X1 U2284 ( .A1(n588), .A2(n2118), .ZN(n582) );
  XNOR2_X1 U2285 ( .A(b[19]), .B(n2299), .ZN(n1636) );
  XNOR2_X1 U2286 ( .A(b[21]), .B(n2301), .ZN(n1634) );
  NAND2_X1 U2287 ( .A1(n685), .A2(n688), .ZN(n369) );
  AOI21_X1 U2288 ( .B1(n629), .B2(n635), .A(n630), .ZN(n628) );
  NOR2_X1 U2289 ( .A1(n1175), .A2(n1178), .ZN(n636) );
  NAND2_X1 U2290 ( .A1(n1175), .A2(n1178), .ZN(n637) );
  NOR2_X1 U2291 ( .A1(n897), .A2(n918), .ZN(n534) );
  NAND2_X1 U2292 ( .A1(n1937), .A2(n672), .ZN(n321) );
  NAND2_X1 U2293 ( .A1(n897), .A2(n918), .ZN(n535) );
  NAND2_X1 U2294 ( .A1(n2126), .A2(n2128), .ZN(n571) );
  AOI21_X1 U2295 ( .B1(n2126), .B2(n1957), .A(n1969), .ZN(n572) );
  NOR2_X1 U2296 ( .A1(n1181), .A2(n1192), .ZN(n644) );
  NAND2_X1 U2297 ( .A1(n1181), .A2(n1192), .ZN(n645) );
  INV_X1 U2298 ( .A(n400), .ZN(n398) );
  NAND2_X1 U2299 ( .A1(n400), .A2(n2122), .ZN(n389) );
  NOR2_X1 U2300 ( .A1(n542), .A2(n547), .ZN(n540) );
  NAND2_X1 U2301 ( .A1(n1031), .A2(n1033), .ZN(n2224) );
  NAND2_X1 U2302 ( .A1(n1031), .A2(n1048), .ZN(n2225) );
  NAND2_X1 U2303 ( .A1(n1033), .A2(n1048), .ZN(n2226) );
  NAND3_X1 U2304 ( .A1(n2224), .A2(n2225), .A3(n2226), .ZN(n1026) );
  OAI21_X1 U2305 ( .B1(n566), .B2(n538), .A(n539), .ZN(n2227) );
  OR2_X1 U2306 ( .A1(n2244), .A2(n1647), .ZN(n2228) );
  OR2_X1 U2307 ( .A1(n1646), .A2(n2263), .ZN(n2229) );
  NAND2_X1 U2308 ( .A1(n2228), .A2(n2229), .ZN(n1352) );
  XNOR2_X1 U2309 ( .A(n2024), .B(b[8]), .ZN(n1647) );
  XNOR2_X1 U2310 ( .A(b[9]), .B(n2299), .ZN(n1646) );
  INV_X1 U2311 ( .A(n490), .ZN(n492) );
  OAI21_X1 U2312 ( .B1(n503), .B2(n495), .A(n496), .ZN(n490) );
  INV_X1 U2313 ( .A(n383), .ZN(n381) );
  AOI21_X1 U2314 ( .B1(n383), .B2(n2181), .A(n376), .ZN(n372) );
  OAI21_X1 U2315 ( .B1(n390), .B2(n384), .A(n387), .ZN(n383) );
  NAND2_X1 U2316 ( .A1(n1099), .A2(n1110), .ZN(n598) );
  AOI21_X1 U2317 ( .B1(n2043), .B2(n472), .A(n459), .ZN(n457) );
  INV_X1 U2318 ( .A(n2146), .ZN(n2271) );
  OAI21_X1 U2319 ( .B1(n1998), .B2(n1942), .A(n2328), .ZN(n1434) );
  AOI21_X1 U2320 ( .B1(n2040), .B2(n2009), .A(n2105), .ZN(n2230) );
  OAI22_X1 U2321 ( .A1(n1997), .A2(n1620), .B1(n1619), .B2(n2023), .ZN(n1326)
         );
  OAI22_X1 U2322 ( .A1(n2022), .A2(n1626), .B1(n1625), .B2(n2023), .ZN(n1332)
         );
  OAI22_X1 U2323 ( .A1(n1997), .A2(n1621), .B1(n2023), .B2(n1620), .ZN(n1327)
         );
  OAI22_X1 U2324 ( .A1(n2022), .A2(n1625), .B1(n2023), .B2(n1624), .ZN(n1331)
         );
  OAI22_X1 U2325 ( .A1(n2022), .A2(n1629), .B1(n2023), .B2(n1628), .ZN(n1335)
         );
  NAND2_X1 U2326 ( .A1(n2076), .A2(n996), .ZN(n2231) );
  NAND2_X1 U2327 ( .A1(n2076), .A2(n1217), .ZN(n2232) );
  NAND2_X1 U2328 ( .A1(n996), .A2(n1217), .ZN(n2233) );
  NAND3_X1 U2329 ( .A1(n2231), .A2(n2232), .A3(n2233), .ZN(n972) );
  INV_X1 U2330 ( .A(n508), .ZN(n2234) );
  NOR2_X1 U2331 ( .A1(n2254), .A2(n2326), .ZN(n1217) );
  XNOR2_X1 U2332 ( .A(n2014), .B(b[6]), .ZN(n1599) );
  XNOR2_X1 U2333 ( .A(b[7]), .B(n2014), .ZN(n1598) );
  NAND2_X1 U2334 ( .A1(n2127), .A2(n2123), .ZN(n599) );
  INV_X1 U2335 ( .A(n502), .ZN(n668) );
  INV_X1 U2336 ( .A(n439), .ZN(n445) );
  OAI21_X1 U2337 ( .B1(n421), .B2(n402), .A(n405), .ZN(n401) );
  XNOR2_X1 U2338 ( .A(b[3]), .B(n2059), .ZN(n1777) );
  XNOR2_X1 U2339 ( .A(b[7]), .B(n2059), .ZN(n1773) );
  XNOR2_X1 U2340 ( .A(b[1]), .B(n2058), .ZN(n1779) );
  XNOR2_X1 U2341 ( .A(b[5]), .B(n2058), .ZN(n1775) );
  XNOR2_X1 U2342 ( .A(b[9]), .B(n2058), .ZN(n1771) );
  INV_X1 U2343 ( .A(n420), .ZN(n422) );
  NOR2_X1 U2344 ( .A1(n420), .A2(n347), .ZN(n345) );
  NOR2_X1 U2345 ( .A1(n336), .A2(n334), .ZN(n332) );
  NAND2_X1 U2346 ( .A1(n709), .A2(n716), .ZN(n409) );
  OAI21_X1 U2347 ( .B1(n631), .B2(n634), .A(n632), .ZN(n630) );
  NAND2_X1 U2348 ( .A1(n540), .A2(n552), .ZN(n538) );
  NOR2_X1 U2349 ( .A1(n571), .A2(n2091), .ZN(n567) );
  NOR2_X1 U2350 ( .A1(n1071), .A2(n1084), .ZN(n590) );
  OAI21_X1 U2351 ( .B1(n590), .B2(n593), .A(n591), .ZN(n589) );
  NOR2_X1 U2352 ( .A1(n590), .A2(n592), .ZN(n588) );
  NAND2_X1 U2353 ( .A1(n2011), .A2(n670), .ZN(n516) );
  INV_X1 U2354 ( .A(n534), .ZN(n672) );
  AOI21_X1 U2355 ( .B1(n526), .B2(n511), .A(n512), .ZN(n506) );
  NOR2_X1 U2356 ( .A1(n520), .A2(n513), .ZN(n511) );
  OAI21_X1 U2357 ( .B1(n531), .B2(n535), .A(n532), .ZN(n526) );
  NOR2_X1 U2358 ( .A1(n857), .A2(n876), .ZN(n520) );
  OAI21_X1 U2359 ( .B1(n572), .B2(n569), .A(n570), .ZN(n568) );
  INV_X1 U2360 ( .A(n474), .ZN(n472) );
  NOR2_X1 U2361 ( .A1(n554), .A2(n2090), .ZN(n545) );
  OAI21_X1 U2362 ( .B1(n555), .B2(n2090), .A(n550), .ZN(n546) );
  NAND2_X1 U2363 ( .A1(n941), .A2(n962), .ZN(n550) );
  OAI21_X1 U2364 ( .B1(n564), .B2(n558), .A(n559), .ZN(n553) );
  INV_X1 U2365 ( .A(n2230), .ZN(n508) );
  NAND2_X1 U2366 ( .A1(n839), .A2(n856), .ZN(n514) );
  NAND2_X1 U2367 ( .A1(n983), .A2(n1002), .ZN(n564) );
  OAI22_X1 U2368 ( .A1(n2036), .A2(n1671), .B1(n2266), .B2(n1670), .ZN(n1375)
         );
  OAI22_X1 U2369 ( .A1(n2035), .A2(n1672), .B1(n1671), .B2(n2266), .ZN(n1376)
         );
  OAI22_X1 U2370 ( .A1(n2035), .A2(n1670), .B1(n1669), .B2(n2266), .ZN(n1374)
         );
  OAI22_X1 U2371 ( .A1(n2245), .A2(n1676), .B1(n1675), .B2(n2265), .ZN(n1380)
         );
  OAI22_X1 U2372 ( .A1(n2036), .A2(n1669), .B1(n2265), .B2(n1668), .ZN(n1373)
         );
  OAI22_X1 U2373 ( .A1(n2036), .A2(n1677), .B1(n2266), .B2(n1676), .ZN(n1381)
         );
  OAI22_X1 U2374 ( .A1(n2036), .A2(n1679), .B1(n2265), .B2(n1678), .ZN(n1383)
         );
  OAI22_X1 U2375 ( .A1(n2245), .A2(n1675), .B1(n2265), .B2(n1674), .ZN(n1379)
         );
  OAI22_X1 U2376 ( .A1(n2036), .A2(n1674), .B1(n1673), .B2(n2265), .ZN(n1378)
         );
  OAI22_X1 U2377 ( .A1(n2036), .A2(n1673), .B1(n2265), .B2(n1672), .ZN(n1377)
         );
  XNOR2_X1 U2378 ( .A(b[15]), .B(n2308), .ZN(n1690) );
  XNOR2_X1 U2379 ( .A(b[17]), .B(n2309), .ZN(n1688) );
  XNOR2_X1 U2380 ( .A(b[21]), .B(n1994), .ZN(n1684) );
  XNOR2_X1 U2381 ( .A(b[11]), .B(n1994), .ZN(n1694) );
  XNOR2_X1 U2382 ( .A(b[19]), .B(n2309), .ZN(n1686) );
  XNOR2_X1 U2383 ( .A(b[13]), .B(n1993), .ZN(n1692) );
  NOR2_X1 U2384 ( .A1(n2084), .A2(n480), .ZN(n478) );
  OAI21_X1 U2385 ( .B1(n492), .B2(n480), .A(n481), .ZN(n479) );
  INV_X1 U2386 ( .A(n480), .ZN(n666) );
  NOR2_X1 U2387 ( .A1(n456), .A2(n480), .ZN(n454) );
  NAND2_X1 U2388 ( .A1(n877), .A2(n896), .ZN(n532) );
  XNOR2_X1 U2389 ( .A(b[13]), .B(n2299), .ZN(n1642) );
  XNOR2_X1 U2390 ( .A(b[15]), .B(n2301), .ZN(n1640) );
  XNOR2_X1 U2391 ( .A(b[11]), .B(n2301), .ZN(n1644) );
  XNOR2_X1 U2392 ( .A(b[17]), .B(n2300), .ZN(n1638) );
  OAI22_X1 U2393 ( .A1(n1997), .A2(n1627), .B1(n2023), .B2(n1626), .ZN(n1333)
         );
  OAI21_X1 U2394 ( .B1(n594), .B2(n582), .A(n583), .ZN(n581) );
  NOR2_X1 U2395 ( .A1(n1171), .A2(n1174), .ZN(n633) );
  NAND2_X1 U2396 ( .A1(n1171), .A2(n1174), .ZN(n634) );
  AOI21_X1 U2397 ( .B1(n508), .B2(n478), .A(n479), .ZN(n477) );
  AOI21_X1 U2398 ( .B1(n508), .B2(n465), .A(n466), .ZN(n464) );
  AOI21_X1 U2399 ( .B1(n508), .B2(n668), .A(n501), .ZN(n499) );
  AOI21_X1 U2400 ( .B1(n508), .B2(n2078), .A(n2079), .ZN(n488) );
  OAI22_X1 U2401 ( .A1(n2168), .A2(n1484), .B1(n2255), .B2(n1483), .ZN(n1195)
         );
  OAI22_X1 U2402 ( .A1(n2168), .A2(n1488), .B1(n2255), .B2(n1487), .ZN(n1199)
         );
  OAI22_X1 U2403 ( .A1(n2167), .A2(n1490), .B1(n2255), .B2(n1489), .ZN(n1201)
         );
  OAI22_X1 U2404 ( .A1(n2167), .A2(n1486), .B1(n2254), .B2(n1485), .ZN(n1197)
         );
  OAI22_X1 U2405 ( .A1(n2166), .A2(n1492), .B1(n2255), .B2(n1491), .ZN(n1203)
         );
  XNOR2_X1 U2406 ( .A(b[11]), .B(n2277), .ZN(n1519) );
  XNOR2_X1 U2407 ( .A(b[17]), .B(n2277), .ZN(n1513) );
  XNOR2_X1 U2408 ( .A(b[13]), .B(n2277), .ZN(n1517) );
  XNOR2_X1 U2409 ( .A(b[21]), .B(n2277), .ZN(n1509) );
  XNOR2_X1 U2410 ( .A(b[19]), .B(n2277), .ZN(n1511) );
  XNOR2_X1 U2411 ( .A(b[15]), .B(n2277), .ZN(n1515) );
  AOI21_X1 U2412 ( .B1(n565), .B2(n1975), .A(n2213), .ZN(n551) );
  INV_X1 U2413 ( .A(n553), .ZN(n555) );
  AOI21_X1 U2414 ( .B1(n553), .B2(n540), .A(n541), .ZN(n539) );
  OAI22_X1 U2415 ( .A1(n1997), .A2(n1624), .B1(n1623), .B2(n2023), .ZN(n1330)
         );
  OAI22_X1 U2416 ( .A1(n2022), .A2(n1622), .B1(n1621), .B2(n2023), .ZN(n1328)
         );
  OAI22_X1 U2417 ( .A1(n1997), .A2(n1619), .B1(n2023), .B2(n1618), .ZN(n1325)
         );
  OAI22_X1 U2418 ( .A1(n2022), .A2(n1623), .B1(n2023), .B2(n1622), .ZN(n1329)
         );
  INV_X1 U2419 ( .A(n428), .ZN(n661) );
  OAI21_X1 U2420 ( .B1(n428), .B2(n436), .A(n429), .ZN(n427) );
  NAND2_X1 U2421 ( .A1(n727), .A2(n736), .ZN(n429) );
  INV_X1 U2422 ( .A(n772), .ZN(n773) );
  AOI21_X1 U2423 ( .B1(n333), .B2(n2136), .A(n2137), .ZN(n327) );
  OAI21_X1 U2424 ( .B1(n337), .B2(n334), .A(n335), .ZN(n333) );
  NAND2_X1 U2425 ( .A1(n717), .A2(n726), .ZN(n418) );
  INV_X1 U2426 ( .A(n746), .ZN(n747) );
  INV_X1 U2427 ( .A(n2227), .ZN(n536) );
  NAND2_X1 U2428 ( .A1(n1165), .A2(n1170), .ZN(n632) );
  INV_X1 U2429 ( .A(n2075), .ZN(n565) );
  XNOR2_X1 U2430 ( .A(b[19]), .B(n2031), .ZN(n1611) );
  XNOR2_X1 U2431 ( .A(b[17]), .B(n2296), .ZN(n1613) );
  XNOR2_X1 U2432 ( .A(b[21]), .B(n1944), .ZN(n1609) );
  XNOR2_X1 U2433 ( .A(b[11]), .B(n1945), .ZN(n1619) );
  XNOR2_X1 U2434 ( .A(b[13]), .B(n1944), .ZN(n1617) );
  XNOR2_X1 U2435 ( .A(b[15]), .B(n2296), .ZN(n1615) );
  NAND2_X1 U2436 ( .A1(n2227), .A2(n450), .ZN(n2235) );
  INV_X1 U2437 ( .A(n451), .ZN(n2236) );
  OAI22_X1 U2438 ( .A1(n2223), .A2(n1733), .B1(n1732), .B2(n2272), .ZN(n2237)
         );
  NOR2_X1 U2439 ( .A1(n505), .A2(n452), .ZN(n450) );
  NAND2_X1 U2440 ( .A1(n478), .A2(n507), .ZN(n476) );
  NAND2_X1 U2441 ( .A1(n465), .A2(n507), .ZN(n463) );
  NAND2_X1 U2442 ( .A1(n507), .A2(n2078), .ZN(n487) );
  NAND2_X1 U2443 ( .A1(n507), .A2(n668), .ZN(n498) );
  OAI22_X1 U2444 ( .A1(n2005), .A2(n1570), .B1(n1569), .B2(n2259), .ZN(n1278)
         );
  OAI22_X1 U2445 ( .A1(n2138), .A2(n1575), .B1(n1992), .B2(n1574), .ZN(n1283)
         );
  OAI22_X1 U2446 ( .A1(n2138), .A2(n1571), .B1(n2259), .B2(n1570), .ZN(n1279)
         );
  OAI22_X1 U2447 ( .A1(n1569), .A2(n2138), .B1(n2259), .B2(n1568), .ZN(n1277)
         );
  OAI22_X1 U2448 ( .A1(n2138), .A2(n1573), .B1(n1992), .B2(n1572), .ZN(n1281)
         );
  OAI22_X1 U2449 ( .A1(n2005), .A2(n1580), .B1(n1579), .B2(n2259), .ZN(n1288)
         );
  OAI22_X1 U2450 ( .A1(n1579), .A2(n2138), .B1(n1992), .B2(n1578), .ZN(n1287)
         );
  OAI22_X1 U2451 ( .A1(n2138), .A2(n1578), .B1(n1577), .B2(n1992), .ZN(n1286)
         );
  OAI22_X1 U2452 ( .A1(n2138), .A2(n1577), .B1(n2259), .B2(n1576), .ZN(n1285)
         );
  OAI22_X1 U2453 ( .A1(n2138), .A2(n1572), .B1(n1571), .B2(n2259), .ZN(n1280)
         );
  OAI22_X1 U2454 ( .A1(n2138), .A2(n1574), .B1(n1573), .B2(n2259), .ZN(n1282)
         );
  NAND2_X1 U2455 ( .A1(n382), .A2(n2181), .ZN(n371) );
  NOR2_X1 U2456 ( .A1(n737), .A2(n748), .ZN(n435) );
  OAI21_X1 U2457 ( .B1(n2195), .B2(n550), .A(n543), .ZN(n541) );
  OAI22_X1 U2458 ( .A1(n1948), .A2(n1535), .B1(n1534), .B2(n2021), .ZN(n1244)
         );
  OAI22_X1 U2459 ( .A1(n1934), .A2(n1537), .B1(n1536), .B2(n2021), .ZN(n1246)
         );
  OAI22_X1 U2460 ( .A1(n1934), .A2(n1543), .B1(n1542), .B2(n2256), .ZN(n1252)
         );
  OAI22_X1 U2461 ( .A1(n1934), .A2(n1533), .B1(n1532), .B2(n2256), .ZN(n692)
         );
  OAI22_X1 U2462 ( .A1(n1948), .A2(n1539), .B1(n1538), .B2(n2256), .ZN(n1248)
         );
  OAI22_X1 U2463 ( .A1(n1934), .A2(n1982), .B1(n1556), .B2(n2021), .ZN(n1184)
         );
  OAI22_X1 U2464 ( .A1(n1948), .A2(n1541), .B1(n1540), .B2(n2021), .ZN(n1250)
         );
  INV_X1 U2465 ( .A(n401), .ZN(n399) );
  AOI21_X1 U2466 ( .B1(n401), .B2(n2122), .A(n394), .ZN(n390) );
  NAND2_X1 U2467 ( .A1(n749), .A2(n760), .ZN(n439) );
  NOR2_X1 U2468 ( .A1(n749), .A2(n760), .ZN(n438) );
  INV_X1 U2469 ( .A(n345), .ZN(n343) );
  NAND2_X1 U2470 ( .A1(n345), .A2(n2135), .ZN(n336) );
  NAND2_X1 U2471 ( .A1(n694), .A2(n689), .ZN(n378) );
  INV_X1 U2472 ( .A(n706), .ZN(n707) );
  XNOR2_X1 U2473 ( .A(n462), .B(n313), .ZN(product[33]) );
  NAND2_X1 U2474 ( .A1(n805), .A2(n820), .ZN(n496) );
  OAI22_X1 U2475 ( .A1(n2169), .A2(n1508), .B1(n1507), .B2(n1946), .ZN(n682)
         );
  OAI22_X1 U2476 ( .A1(n2169), .A2(n1518), .B1(n1517), .B2(n1946), .ZN(n1228)
         );
  OAI22_X1 U2477 ( .A1(n2170), .A2(n1514), .B1(n1513), .B2(n1946), .ZN(n1224)
         );
  XNOR2_X1 U2478 ( .A(n1237), .B(n1215), .ZN(n939) );
  OAI22_X1 U2479 ( .A1(n2169), .A2(n1510), .B1(n1509), .B2(n1946), .ZN(n1220)
         );
  OR2_X1 U2480 ( .A1(n1215), .A2(n1237), .ZN(n938) );
  OAI22_X1 U2481 ( .A1(n2169), .A2(n1512), .B1(n1511), .B2(n1946), .ZN(n1222)
         );
  OAI22_X1 U2482 ( .A1(n2169), .A2(n1516), .B1(n1515), .B2(n1946), .ZN(n1226)
         );
  XNOR2_X1 U2483 ( .A(n437), .B(n311), .ZN(product[35]) );
  XNOR2_X1 U2484 ( .A(n430), .B(n310), .ZN(product[36]) );
  NAND2_X1 U2485 ( .A1(n1071), .A2(n1084), .ZN(n591) );
  OAI22_X1 U2486 ( .A1(n2243), .A2(n1648), .B1(n2263), .B2(n1647), .ZN(n1353)
         );
  OAI22_X1 U2487 ( .A1(n2243), .A2(n1652), .B1(n1931), .B2(n1651), .ZN(n1357)
         );
  OAI22_X1 U2488 ( .A1(n2243), .A2(n1649), .B1(n1648), .B2(n2263), .ZN(n1354)
         );
  OAI22_X1 U2489 ( .A1(n2243), .A2(n1653), .B1(n1652), .B2(n2163), .ZN(n1358)
         );
  OAI22_X1 U2490 ( .A1(n2243), .A2(n1645), .B1(n1644), .B2(n2263), .ZN(n1350)
         );
  OAI22_X1 U2491 ( .A1(n2243), .A2(n1654), .B1(n1931), .B2(n1653), .ZN(n1359)
         );
  OAI22_X1 U2492 ( .A1(n2244), .A2(n1644), .B1(n2263), .B2(n1643), .ZN(n1349)
         );
  OAI22_X1 U2493 ( .A1(n2243), .A2(n1650), .B1(n2263), .B2(n1649), .ZN(n1355)
         );
  OAI22_X1 U2494 ( .A1(n2243), .A2(n1655), .B1(n1654), .B2(n2163), .ZN(n1360)
         );
  OAI22_X1 U2495 ( .A1(n2244), .A2(n1651), .B1(n1650), .B2(n2263), .ZN(n1356)
         );
  OAI22_X1 U2496 ( .A1(n2244), .A2(n1646), .B1(n2263), .B2(n1645), .ZN(n1351)
         );
  XNOR2_X1 U2497 ( .A(n419), .B(n309), .ZN(product[37]) );
  OAI22_X1 U2498 ( .A1(n1941), .A2(n1695), .B1(n1694), .B2(n2268), .ZN(n1398)
         );
  OAI22_X1 U2499 ( .A1(n2247), .A2(n1704), .B1(n2268), .B2(n1703), .ZN(n1407)
         );
  OAI22_X1 U2500 ( .A1(n1941), .A2(n1701), .B1(n1700), .B2(n2268), .ZN(n1404)
         );
  OAI22_X1 U2501 ( .A1(n1941), .A2(n1702), .B1(n2267), .B2(n1701), .ZN(n1405)
         );
  OAI22_X1 U2502 ( .A1(n1955), .A2(n1698), .B1(n2268), .B2(n1697), .ZN(n1401)
         );
  OAI22_X1 U2503 ( .A1(n1941), .A2(n1694), .B1(n2268), .B2(n1693), .ZN(n1397)
         );
  OAI22_X1 U2504 ( .A1(n1941), .A2(n1696), .B1(n2268), .B2(n1695), .ZN(n1399)
         );
  OAI22_X1 U2505 ( .A1(n1941), .A2(n1700), .B1(n2268), .B2(n1699), .ZN(n1403)
         );
  OAI22_X1 U2506 ( .A1(n1955), .A2(n1699), .B1(n1698), .B2(n2267), .ZN(n1402)
         );
  OAI22_X1 U2507 ( .A1(n1955), .A2(n1705), .B1(n1704), .B2(n2267), .ZN(n1408)
         );
  OAI22_X1 U2508 ( .A1(n1955), .A2(n1703), .B1(n1702), .B2(n2267), .ZN(n1406)
         );
  OAI22_X1 U2509 ( .A1(n1955), .A2(n1697), .B1(n1696), .B2(n2267), .ZN(n1400)
         );
  XNOR2_X1 U2510 ( .A(n410), .B(n308), .ZN(product[38]) );
  NAND2_X1 U2511 ( .A1(n761), .A2(n774), .ZN(n461) );
  NOR2_X1 U2512 ( .A1(n2006), .A2(n774), .ZN(n460) );
  OAI22_X1 U2513 ( .A1(n2162), .A2(n2316), .B1(n1731), .B2(n2270), .ZN(n1191)
         );
  OAI22_X1 U2514 ( .A1(n2162), .A2(n1718), .B1(n1717), .B2(n2097), .ZN(n1420)
         );
  OAI22_X1 U2515 ( .A1(n2161), .A2(n1711), .B1(n2270), .B2(n1710), .ZN(n1413)
         );
  OAI22_X1 U2516 ( .A1(n2248), .A2(n1708), .B1(n1707), .B2(n2270), .ZN(n874)
         );
  OAI22_X1 U2517 ( .A1(n2162), .A2(n1713), .B1(n2097), .B2(n1712), .ZN(n1415)
         );
  OAI22_X1 U2518 ( .A1(n2162), .A2(n1717), .B1(n2096), .B2(n1716), .ZN(n1419)
         );
  OAI22_X1 U2519 ( .A1(n2162), .A2(n1716), .B1(n1715), .B2(n2097), .ZN(n1418)
         );
  OAI22_X1 U2520 ( .A1(n2248), .A2(n1709), .B1(n2096), .B2(n1708), .ZN(n1411)
         );
  OAI22_X1 U2521 ( .A1(n2248), .A2(n1710), .B1(n1709), .B2(n2095), .ZN(n1412)
         );
  OAI22_X1 U2522 ( .A1(n2248), .A2(n1712), .B1(n1711), .B2(n2270), .ZN(n1414)
         );
  XNOR2_X1 U2523 ( .A(b[21]), .B(n2318), .ZN(n1734) );
  XNOR2_X1 U2524 ( .A(b[11]), .B(n2318), .ZN(n1744) );
  XNOR2_X1 U2525 ( .A(b[15]), .B(n2318), .ZN(n1740) );
  XNOR2_X1 U2526 ( .A(b[17]), .B(n2318), .ZN(n1738) );
  XNOR2_X1 U2527 ( .A(b[19]), .B(n2318), .ZN(n1736) );
  XNOR2_X1 U2528 ( .A(b[13]), .B(n2318), .ZN(n1742) );
  OAI22_X1 U2529 ( .A1(n2248), .A2(n1714), .B1(n1713), .B2(n2095), .ZN(n1416)
         );
  XNOR2_X1 U2530 ( .A(b[17]), .B(n2322), .ZN(n1763) );
  XNOR2_X1 U2531 ( .A(b[13]), .B(n2323), .ZN(n1767) );
  XNOR2_X1 U2532 ( .A(b[21]), .B(n2322), .ZN(n1759) );
  XNOR2_X1 U2533 ( .A(b[15]), .B(n2323), .ZN(n1765) );
  XNOR2_X1 U2534 ( .A(b[11]), .B(n2323), .ZN(n1769) );
  XNOR2_X1 U2535 ( .A(b[19]), .B(n2323), .ZN(n1761) );
  OAI22_X1 U2536 ( .A1(n2167), .A2(n1483), .B1(n1482), .B2(n2254), .ZN(n676)
         );
  OAI22_X1 U2537 ( .A1(n2167), .A2(n1485), .B1(n1484), .B2(n2254), .ZN(n1196)
         );
  OAI22_X1 U2538 ( .A1(n2167), .A2(n1491), .B1(n1490), .B2(n2255), .ZN(n1202)
         );
  OAI22_X1 U2539 ( .A1(n2168), .A2(n1487), .B1(n1486), .B2(n2254), .ZN(n1198)
         );
  OAI22_X1 U2540 ( .A1(n2168), .A2(n1497), .B1(n1496), .B2(n2255), .ZN(n1208)
         );
  OAI22_X1 U2541 ( .A1(n2168), .A2(n1496), .B1(n2254), .B2(n1495), .ZN(n1207)
         );
  OAI22_X1 U2542 ( .A1(n2167), .A2(n1494), .B1(n2255), .B2(n1493), .ZN(n1205)
         );
  OAI22_X1 U2543 ( .A1(n2168), .A2(n1495), .B1(n1494), .B2(n2254), .ZN(n1206)
         );
  OAI22_X1 U2544 ( .A1(n2047), .A2(n1502), .B1(n2254), .B2(n1501), .ZN(n1213)
         );
  OAI22_X1 U2545 ( .A1(n2166), .A2(n1501), .B1(n1500), .B2(n2255), .ZN(n1212)
         );
  OAI22_X1 U2546 ( .A1(n2167), .A2(n1489), .B1(n1488), .B2(n2254), .ZN(n1200)
         );
  OAI22_X1 U2547 ( .A1(n2168), .A2(n1493), .B1(n1492), .B2(n2255), .ZN(n1204)
         );
  OAI22_X1 U2548 ( .A1(n2048), .A2(n1500), .B1(n2254), .B2(n1499), .ZN(n1211)
         );
  OAI22_X1 U2549 ( .A1(n2048), .A2(n1503), .B1(n1502), .B2(n2254), .ZN(n1214)
         );
  OAI22_X1 U2550 ( .A1(n2276), .A2(n2238), .B1(n1506), .B2(n2255), .ZN(n1182)
         );
  OAI22_X1 U2551 ( .A1(n2238), .A2(n1504), .B1(n2255), .B2(n1503), .ZN(n1215)
         );
  OAI22_X1 U2552 ( .A1(n2047), .A2(n1498), .B1(n2255), .B2(n1497), .ZN(n1209)
         );
  INV_X1 U2553 ( .A(n2040), .ZN(n524) );
  AOI21_X1 U2554 ( .B1(n2040), .B2(n670), .A(n519), .ZN(n517) );
  OAI22_X1 U2555 ( .A1(n2035), .A2(n1661), .B1(n2266), .B2(n1660), .ZN(n1365)
         );
  OAI22_X1 U2556 ( .A1(n2035), .A2(n1660), .B1(n1659), .B2(n2266), .ZN(n1364)
         );
  OAI22_X1 U2557 ( .A1(n2245), .A2(n1663), .B1(n2265), .B2(n1662), .ZN(n1367)
         );
  OAI22_X1 U2558 ( .A1(n2245), .A2(n2306), .B1(n1681), .B2(n2266), .ZN(n1189)
         );
  OAI22_X1 U2559 ( .A1(n2245), .A2(n1664), .B1(n1663), .B2(n2266), .ZN(n1368)
         );
  OAI22_X1 U2560 ( .A1(n2035), .A2(n1665), .B1(n2265), .B2(n1664), .ZN(n1369)
         );
  OAI22_X1 U2561 ( .A1(n2245), .A2(n1658), .B1(n1657), .B2(n2266), .ZN(n802)
         );
  OAI22_X1 U2562 ( .A1(n2246), .A2(n1667), .B1(n2266), .B2(n1666), .ZN(n1371)
         );
  OAI22_X1 U2563 ( .A1(n2246), .A2(n1662), .B1(n1661), .B2(n2266), .ZN(n1366)
         );
  OAI22_X1 U2564 ( .A1(n2036), .A2(n1666), .B1(n1665), .B2(n2266), .ZN(n1370)
         );
  OAI22_X1 U2565 ( .A1(n2035), .A2(n1659), .B1(n2265), .B2(n1658), .ZN(n1363)
         );
  OAI22_X1 U2566 ( .A1(n2245), .A2(n1680), .B1(n1679), .B2(n2266), .ZN(n1384)
         );
  OAI22_X1 U2567 ( .A1(n2035), .A2(n1678), .B1(n1677), .B2(n2265), .ZN(n1382)
         );
  OAI22_X1 U2568 ( .A1(n2246), .A2(n1668), .B1(n1667), .B2(n2265), .ZN(n1372)
         );
  XNOR2_X1 U2569 ( .A(n397), .B(n307), .ZN(product[39]) );
  NOR2_X1 U2570 ( .A1(n775), .A2(n788), .ZN(n473) );
  NAND2_X1 U2571 ( .A1(n775), .A2(n788), .ZN(n474) );
  INV_X1 U2572 ( .A(n1954), .ZN(n837) );
  NAND2_X1 U2573 ( .A1(n356), .A2(n2134), .ZN(n347) );
  NAND2_X1 U2574 ( .A1(n332), .A2(n2136), .ZN(n326) );
  OAI21_X1 U2575 ( .B1(n2038), .B2(n521), .A(n514), .ZN(n512) );
  XNOR2_X1 U2576 ( .A(n388), .B(n306), .ZN(product[40]) );
  OAI22_X1 U2577 ( .A1(n2028), .A2(n1593), .B1(n1592), .B2(n2262), .ZN(n1300)
         );
  OAI22_X1 U2578 ( .A1(n2028), .A2(n1589), .B1(n1588), .B2(n2262), .ZN(n1296)
         );
  OAI22_X1 U2579 ( .A1(n2028), .A2(n1587), .B1(n1586), .B2(n2262), .ZN(n1294)
         );
  OAI22_X1 U2580 ( .A1(n2027), .A2(n1591), .B1(n1590), .B2(n2262), .ZN(n1298)
         );
  OAI22_X1 U2581 ( .A1(n2028), .A2(n1583), .B1(n1582), .B2(n2261), .ZN(n724)
         );
  OAI22_X1 U2582 ( .A1(n2028), .A2(n1585), .B1(n1584), .B2(n2262), .ZN(n1292)
         );
  OAI22_X1 U2583 ( .A1(n2027), .A2(n2295), .B1(n1606), .B2(n2261), .ZN(n1186)
         );
  XNOR2_X1 U2584 ( .A(n379), .B(n305), .ZN(product[41]) );
  OAI22_X1 U2585 ( .A1(n2223), .A2(n2321), .B1(n1756), .B2(n2272), .ZN(n1192)
         );
  OAI22_X1 U2586 ( .A1(n2223), .A2(n1738), .B1(n2271), .B2(n1737), .ZN(n1439)
         );
  OAI22_X1 U2587 ( .A1(n2223), .A2(n1741), .B1(n1740), .B2(n2272), .ZN(n1442)
         );
  INV_X1 U2588 ( .A(n916), .ZN(n917) );
  OAI22_X1 U2589 ( .A1(n2223), .A2(n1740), .B1(n2271), .B2(n1739), .ZN(n1441)
         );
  OAI22_X1 U2590 ( .A1(n2223), .A2(n1739), .B1(n1738), .B2(n2271), .ZN(n1440)
         );
  OAI22_X1 U2591 ( .A1(n2223), .A2(n1734), .B1(n2272), .B2(n1733), .ZN(n1435)
         );
  OAI22_X1 U2592 ( .A1(n2223), .A2(n1736), .B1(n2271), .B2(n1735), .ZN(n1437)
         );
  OAI22_X1 U2593 ( .A1(n2223), .A2(n1742), .B1(n2272), .B2(n1741), .ZN(n1443)
         );
  OAI22_X1 U2594 ( .A1(n2215), .A2(n1735), .B1(n1734), .B2(n2271), .ZN(n1436)
         );
  OAI22_X1 U2595 ( .A1(n2215), .A2(n1737), .B1(n1736), .B2(n2272), .ZN(n1438)
         );
  OAI22_X1 U2596 ( .A1(n2250), .A2(n1743), .B1(n1742), .B2(n2271), .ZN(n1444)
         );
  OAI22_X1 U2597 ( .A1(n2250), .A2(n1733), .B1(n1732), .B2(n2272), .ZN(n916)
         );
  XNOR2_X1 U2598 ( .A(n353), .B(n303), .ZN(product[43]) );
  OAI22_X1 U2599 ( .A1(n2223), .A2(n1753), .B1(n1752), .B2(n2271), .ZN(n1454)
         );
  OAI22_X1 U2600 ( .A1(n2223), .A2(n1747), .B1(n1746), .B2(n2272), .ZN(n1448)
         );
  OAI22_X1 U2601 ( .A1(n2223), .A2(n1750), .B1(n2272), .B2(n1749), .ZN(n1451)
         );
  OAI22_X1 U2602 ( .A1(n2223), .A2(n1749), .B1(n1748), .B2(n2271), .ZN(n1450)
         );
  OAI22_X1 U2603 ( .A1(n2223), .A2(n1745), .B1(n1744), .B2(n2271), .ZN(n1446)
         );
  OAI22_X1 U2604 ( .A1(n2223), .A2(n1748), .B1(n2272), .B2(n1747), .ZN(n1449)
         );
  OAI22_X1 U2605 ( .A1(n2223), .A2(n1744), .B1(n2272), .B2(n1743), .ZN(n1445)
         );
  OAI22_X1 U2606 ( .A1(n2215), .A2(n1746), .B1(n2271), .B2(n1745), .ZN(n1447)
         );
  OAI22_X1 U2607 ( .A1(n2223), .A2(n1754), .B1(n2271), .B2(n1753), .ZN(n1455)
         );
  OAI22_X1 U2608 ( .A1(n2223), .A2(n1752), .B1(n2271), .B2(n1751), .ZN(n1453)
         );
  OAI22_X1 U2609 ( .A1(n2215), .A2(n1751), .B1(n1750), .B2(n2272), .ZN(n1452)
         );
  OAI22_X1 U2610 ( .A1(n2250), .A2(n1755), .B1(n1754), .B2(n2271), .ZN(n1456)
         );
  INV_X1 U2611 ( .A(n346), .ZN(n344) );
  AOI21_X1 U2612 ( .B1(n346), .B2(n2135), .A(n339), .ZN(n337) );
  OAI22_X1 U2613 ( .A1(n1997), .A2(n1613), .B1(n2023), .B2(n1612), .ZN(n1319)
         );
  OAI22_X1 U2614 ( .A1(n1997), .A2(n1612), .B1(n1611), .B2(n2023), .ZN(n1318)
         );
  OAI22_X1 U2615 ( .A1(n1997), .A2(n1610), .B1(n1609), .B2(n2023), .ZN(n1316)
         );
  OAI22_X1 U2616 ( .A1(n1997), .A2(n1611), .B1(n2023), .B2(n1610), .ZN(n1317)
         );
  OAI22_X1 U2617 ( .A1(n2022), .A2(n1617), .B1(n2023), .B2(n1616), .ZN(n1323)
         );
  OAI22_X1 U2618 ( .A1(n1997), .A2(n1615), .B1(n2023), .B2(n1614), .ZN(n1321)
         );
  OAI22_X1 U2619 ( .A1(n2041), .A2(n1630), .B1(n1629), .B2(n2023), .ZN(n1336)
         );
  OAI22_X1 U2620 ( .A1(n2041), .A2(n1943), .B1(n1631), .B2(n2023), .ZN(n1187)
         );
  OAI22_X1 U2621 ( .A1(n2022), .A2(n1618), .B1(n1617), .B2(n2023), .ZN(n1324)
         );
  OAI22_X1 U2622 ( .A1(n2022), .A2(n1609), .B1(n2023), .B2(n1608), .ZN(n1315)
         );
  OAI22_X1 U2623 ( .A1(n1997), .A2(n1614), .B1(n1613), .B2(n2023), .ZN(n1320)
         );
  OAI22_X1 U2624 ( .A1(n2022), .A2(n1616), .B1(n1615), .B2(n2023), .ZN(n1322)
         );
  OAI22_X1 U2625 ( .A1(n2022), .A2(n1628), .B1(n1627), .B2(n2023), .ZN(n1334)
         );
  OAI22_X1 U2626 ( .A1(n2022), .A2(n1608), .B1(n1607), .B2(n2023), .ZN(n746)
         );
  XNOR2_X1 U2627 ( .A(n370), .B(n304), .ZN(product[42]) );
  INV_X1 U2628 ( .A(n421), .ZN(n423) );
  OAI21_X1 U2629 ( .B1(n421), .B2(n347), .A(n348), .ZN(n346) );
  OAI22_X1 U2630 ( .A1(n2243), .A2(n1637), .B1(n1636), .B2(n2163), .ZN(n1342)
         );
  OAI22_X1 U2631 ( .A1(n2243), .A2(n1636), .B1(n1931), .B2(n1635), .ZN(n1341)
         );
  OAI22_X1 U2632 ( .A1(n2243), .A2(n1634), .B1(n2263), .B2(n1633), .ZN(n1339)
         );
  OAI22_X1 U2633 ( .A1(n2243), .A2(n1635), .B1(n1634), .B2(n2163), .ZN(n1340)
         );
  OAI22_X1 U2634 ( .A1(n2244), .A2(n1639), .B1(n1638), .B2(n2163), .ZN(n1344)
         );
  OAI22_X1 U2635 ( .A1(n2243), .A2(n1640), .B1(n2263), .B2(n1639), .ZN(n1345)
         );
  OAI22_X1 U2636 ( .A1(n2244), .A2(n1638), .B1(n2263), .B2(n1637), .ZN(n1343)
         );
  OAI22_X1 U2637 ( .A1(n2243), .A2(n1642), .B1(n2263), .B2(n1641), .ZN(n1347)
         );
  OAI22_X1 U2638 ( .A1(n2244), .A2(n1641), .B1(n1640), .B2(n2163), .ZN(n1346)
         );
  OAI22_X1 U2639 ( .A1(n2243), .A2(n1633), .B1(n1632), .B2(n2163), .ZN(n772)
         );
  OAI22_X1 U2640 ( .A1(n2243), .A2(n2303), .B1(n1656), .B2(n2163), .ZN(n1188)
         );
  OAI22_X1 U2641 ( .A1(n2244), .A2(n1643), .B1(n1642), .B2(n2163), .ZN(n1348)
         );
  XNOR2_X1 U2642 ( .A(b[17]), .B(n2304), .ZN(n1663) );
  XNOR2_X1 U2643 ( .A(b[11]), .B(n2304), .ZN(n1669) );
  XNOR2_X1 U2644 ( .A(b[19]), .B(n2305), .ZN(n1661) );
  XNOR2_X1 U2645 ( .A(b[15]), .B(n2305), .ZN(n1665) );
  XNOR2_X1 U2646 ( .A(b[21]), .B(n2001), .ZN(n1659) );
  XNOR2_X1 U2647 ( .A(b[13]), .B(n2002), .ZN(n1667) );
  OAI22_X1 U2648 ( .A1(n1948), .A2(n1544), .B1(n2021), .B2(n1543), .ZN(n1253)
         );
  OAI22_X1 U2649 ( .A1(n1546), .A2(n1948), .B1(n2021), .B2(n1545), .ZN(n1255)
         );
  OAI22_X1 U2650 ( .A1(n1948), .A2(n1552), .B1(n2256), .B2(n1551), .ZN(n1261)
         );
  OAI22_X1 U2651 ( .A1(n1934), .A2(n1549), .B1(n1548), .B2(n2256), .ZN(n1258)
         );
  OAI22_X1 U2652 ( .A1(n1948), .A2(n1548), .B1(n2021), .B2(n1547), .ZN(n1257)
         );
  OAI22_X1 U2653 ( .A1(n1934), .A2(n1555), .B1(n1554), .B2(n2021), .ZN(n1264)
         );
  OAI22_X1 U2654 ( .A1(n1934), .A2(n1547), .B1(n1546), .B2(n2021), .ZN(n1256)
         );
  OAI22_X1 U2655 ( .A1(n1948), .A2(n1545), .B1(n1544), .B2(n2020), .ZN(n1254)
         );
  OAI22_X1 U2656 ( .A1(n1934), .A2(n1550), .B1(n2256), .B2(n1549), .ZN(n1259)
         );
  OAI22_X1 U2657 ( .A1(n1934), .A2(n1554), .B1(n2256), .B2(n1553), .ZN(n1263)
         );
  OAI22_X1 U2658 ( .A1(n1948), .A2(n1551), .B1(n2020), .B2(n1550), .ZN(n1260)
         );
  OAI22_X1 U2659 ( .A1(n1948), .A2(n1553), .B1(n2020), .B2(n1552), .ZN(n1262)
         );
  XNOR2_X1 U2660 ( .A(b[15]), .B(n1952), .ZN(n1565) );
  XNOR2_X1 U2661 ( .A(b[21]), .B(n1952), .ZN(n1559) );
  XNOR2_X1 U2662 ( .A(b[17]), .B(n1952), .ZN(n1563) );
  XNOR2_X1 U2663 ( .A(b[11]), .B(n1953), .ZN(n1569) );
  XNOR2_X1 U2664 ( .A(b[13]), .B(n1952), .ZN(n1567) );
  XNOR2_X1 U2665 ( .A(b[19]), .B(n1953), .ZN(n1561) );
  AOI21_X1 U2666 ( .B1(n454), .B2(n490), .A(n455), .ZN(n453) );
  NAND2_X1 U2667 ( .A1(n454), .A2(n489), .ZN(n452) );
  NAND2_X1 U2668 ( .A1(n525), .A2(n511), .ZN(n505) );
  OAI22_X1 U2669 ( .A1(n2170), .A2(n1522), .B1(n1521), .B2(n1946), .ZN(n1232)
         );
  OAI22_X1 U2670 ( .A1(n2170), .A2(n1521), .B1(n1946), .B2(n1520), .ZN(n1231)
         );
  OAI22_X1 U2671 ( .A1(n2169), .A2(n1519), .B1(n1946), .B2(n1518), .ZN(n1229)
         );
  OAI22_X1 U2672 ( .A1(n2170), .A2(n1520), .B1(n1519), .B2(n1946), .ZN(n1230)
         );
  OAI22_X1 U2673 ( .A1(n2240), .A2(n1525), .B1(n1946), .B2(n1524), .ZN(n1235)
         );
  XNOR2_X1 U2674 ( .A(b[19]), .B(n2282), .ZN(n1536) );
  OAI22_X1 U2675 ( .A1(n2240), .A2(n1524), .B1(n1523), .B2(n1946), .ZN(n1234)
         );
  OAI22_X1 U2676 ( .A1(n2170), .A2(n1523), .B1(n1946), .B2(n1522), .ZN(n1233)
         );
  OAI22_X1 U2677 ( .A1(n2240), .A2(n1529), .B1(n1946), .B2(n1528), .ZN(n1239)
         );
  OAI22_X1 U2678 ( .A1(n2240), .A2(n1526), .B1(n1525), .B2(n1946), .ZN(n1236)
         );
  XNOR2_X1 U2679 ( .A(b[21]), .B(n2282), .ZN(n1534) );
  OAI22_X1 U2680 ( .A1(n2240), .A2(n1528), .B1(n1527), .B2(n1946), .ZN(n1238)
         );
  OAI22_X1 U2681 ( .A1(n2240), .A2(n1530), .B1(n1529), .B2(n1946), .ZN(n1240)
         );
  OAI22_X1 U2682 ( .A1(n2240), .A2(n1527), .B1(n1946), .B2(n1526), .ZN(n1237)
         );
  XNOR2_X1 U2683 ( .A(b[13]), .B(n2282), .ZN(n1542) );
  XNOR2_X1 U2684 ( .A(b[17]), .B(n2282), .ZN(n1538) );
  XNOR2_X1 U2685 ( .A(b[11]), .B(n2282), .ZN(n1544) );
  XNOR2_X1 U2686 ( .A(b[15]), .B(n2282), .ZN(n1540) );
  XNOR2_X1 U2687 ( .A(n342), .B(n302), .ZN(product[44]) );
  OAI22_X1 U2688 ( .A1(n1987), .A2(n1602), .B1(n2261), .B2(n1601), .ZN(n1309)
         );
  OAI22_X1 U2689 ( .A1(n1988), .A2(n1600), .B1(n2261), .B2(n1599), .ZN(n1307)
         );
  OAI22_X1 U2690 ( .A1(n1988), .A2(n1601), .B1(n1600), .B2(n2261), .ZN(n1308)
         );
  OAI22_X1 U2691 ( .A1(n1987), .A2(n1594), .B1(n2262), .B2(n1593), .ZN(n1301)
         );
  OAI22_X1 U2692 ( .A1(n1988), .A2(n1596), .B1(n2262), .B2(n1595), .ZN(n1303)
         );
  OAI22_X1 U2693 ( .A1(n1987), .A2(n1598), .B1(n2262), .B2(n1597), .ZN(n1305)
         );
  OAI22_X1 U2694 ( .A1(n1988), .A2(n1597), .B1(n1596), .B2(n2261), .ZN(n1304)
         );
  OAI22_X1 U2695 ( .A1(n1987), .A2(n1603), .B1(n1602), .B2(n2262), .ZN(n1310)
         );
  OAI22_X1 U2696 ( .A1(n1987), .A2(n1595), .B1(n1594), .B2(n2262), .ZN(n1302)
         );
  OAI22_X1 U2697 ( .A1(n1987), .A2(n1604), .B1(n2261), .B2(n1603), .ZN(n1311)
         );
  OAI22_X1 U2698 ( .A1(n1988), .A2(n1605), .B1(n1604), .B2(n2261), .ZN(n1312)
         );
  OAI21_X1 U2699 ( .B1(n506), .B2(n452), .A(n453), .ZN(n451) );
  XNOR2_X1 U2700 ( .A(n475), .B(n314), .ZN(product[32]) );
  XOR2_X1 U2701 ( .A(n1978), .B(n321), .Z(product[25]) );
  OAI21_X1 U2702 ( .B1(n1978), .B2(n516), .A(n517), .ZN(n515) );
  OAI21_X1 U2703 ( .B1(n1977), .B2(n2033), .A(n524), .ZN(n522) );
  OAI21_X1 U2704 ( .B1(n1976), .B2(n476), .A(n477), .ZN(n475) );
  OAI21_X1 U2705 ( .B1(n1977), .B2(n2018), .A(n2187), .ZN(n533) );
  OAI21_X1 U2706 ( .B1(n1977), .B2(n463), .A(n464), .ZN(n462) );
  OAI21_X1 U2707 ( .B1(n1978), .B2(n487), .A(n488), .ZN(n486) );
  OAI21_X1 U2708 ( .B1(n1976), .B2(n498), .A(n499), .ZN(n497) );
  OAI21_X1 U2709 ( .B1(n1976), .B2(n2196), .A(n2234), .ZN(n504) );
  OAI22_X1 U2710 ( .A1(n2162), .A2(n1727), .B1(n2096), .B2(n1726), .ZN(n1429)
         );
  OAI22_X1 U2711 ( .A1(n2162), .A2(n1720), .B1(n1719), .B2(n2270), .ZN(n1422)
         );
  OAI22_X1 U2712 ( .A1(n2162), .A2(n1721), .B1(n2096), .B2(n1720), .ZN(n1423)
         );
  OAI22_X1 U2713 ( .A1(n2162), .A2(n1726), .B1(n1725), .B2(n2270), .ZN(n1428)
         );
  OAI22_X1 U2714 ( .A1(n2162), .A2(n1730), .B1(n1729), .B2(n2097), .ZN(n1432)
         );
  OAI22_X1 U2715 ( .A1(n2162), .A2(n1725), .B1(n2270), .B2(n1724), .ZN(n1427)
         );
  OAI22_X1 U2716 ( .A1(n2162), .A2(n1723), .B1(n2096), .B2(n1722), .ZN(n1425)
         );
  OAI22_X1 U2717 ( .A1(n2162), .A2(n1728), .B1(n1727), .B2(n2096), .ZN(n1430)
         );
  OAI22_X1 U2718 ( .A1(n2162), .A2(n1722), .B1(n1721), .B2(n2270), .ZN(n1424)
         );
  OAI22_X1 U2719 ( .A1(n2162), .A2(n1729), .B1(n2097), .B2(n1728), .ZN(n1431)
         );
  OAI22_X1 U2720 ( .A1(n2161), .A2(n1724), .B1(n1723), .B2(n2096), .ZN(n1426)
         );
  INV_X1 U2721 ( .A(n325), .ZN(product[47]) );
  AOI21_X1 U2722 ( .B1(n423), .B2(n356), .A(n359), .ZN(n355) );
  NAND2_X1 U2723 ( .A1(n422), .A2(n356), .ZN(n354) );
  OAI22_X1 U2724 ( .A1(n2242), .A2(n1563), .B1(n1992), .B2(n1562), .ZN(n1271)
         );
  OAI22_X1 U2725 ( .A1(n2242), .A2(n1567), .B1(n1992), .B2(n1566), .ZN(n1275)
         );
  OAI22_X1 U2726 ( .A1(n2117), .A2(n1566), .B1(n1565), .B2(n2259), .ZN(n1274)
         );
  OAI22_X1 U2727 ( .A1(n2117), .A2(n1561), .B1(n1992), .B2(n1560), .ZN(n1269)
         );
  OAI22_X1 U2728 ( .A1(n2117), .A2(n1564), .B1(n1563), .B2(n1992), .ZN(n1272)
         );
  OAI22_X1 U2729 ( .A1(n2116), .A2(n1560), .B1(n1559), .B2(n2259), .ZN(n1268)
         );
  OAI22_X1 U2730 ( .A1(n2116), .A2(n1565), .B1(n1992), .B2(n1564), .ZN(n1273)
         );
  OAI22_X1 U2731 ( .A1(n2116), .A2(n2292), .B1(n1581), .B2(n2259), .ZN(n1185)
         );
  OAI22_X1 U2732 ( .A1(n2117), .A2(n1559), .B1(n1992), .B2(n1558), .ZN(n1267)
         );
  OAI22_X1 U2733 ( .A1(n2242), .A2(n1562), .B1(n1561), .B2(n1992), .ZN(n1270)
         );
  OAI22_X1 U2734 ( .A1(n2242), .A2(n1568), .B1(n1567), .B2(n1992), .ZN(n1276)
         );
  XNOR2_X1 U2735 ( .A(b[17]), .B(n2293), .ZN(n1588) );
  XNOR2_X1 U2736 ( .A(b[15]), .B(n2293), .ZN(n1590) );
  XNOR2_X1 U2737 ( .A(b[13]), .B(n2293), .ZN(n1592) );
  OAI22_X1 U2738 ( .A1(n2116), .A2(n1558), .B1(n1557), .B2(n1992), .ZN(n706)
         );
  XNOR2_X1 U2739 ( .A(b[19]), .B(n2293), .ZN(n1586) );
  XNOR2_X1 U2740 ( .A(b[21]), .B(n2293), .ZN(n1584) );
  XNOR2_X1 U2741 ( .A(b[11]), .B(n2293), .ZN(n1594) );
  XNOR2_X1 U2742 ( .A(a[16]), .B(a[15]), .ZN(n267) );
  OAI21_X1 U2743 ( .B1(n326), .B2(n301), .A(n327), .ZN(n325) );
  NAND2_X1 U2744 ( .A1(n665), .A2(n474), .ZN(n314) );
  OAI21_X1 U2745 ( .B1(n2222), .B2(n431), .A(n432), .ZN(n430) );
  OAI21_X1 U2746 ( .B1(n301), .B2(n420), .A(n421), .ZN(n419) );
  OAI21_X1 U2747 ( .B1(n301), .B2(n438), .A(n439), .ZN(n437) );
  OAI21_X1 U2748 ( .B1(n2222), .B2(n411), .A(n412), .ZN(n410) );
  OAI21_X1 U2749 ( .B1(n301), .B2(n354), .A(n355), .ZN(n353) );
  OAI21_X1 U2750 ( .B1(n2222), .B2(n371), .A(n372), .ZN(n370) );
  OAI21_X1 U2751 ( .B1(n301), .B2(n380), .A(n381), .ZN(n379) );
  OAI21_X1 U2752 ( .B1(n301), .B2(n343), .A(n344), .ZN(n342) );
  OAI21_X1 U2753 ( .B1(n2222), .B2(n398), .A(n399), .ZN(n397) );
  OAI21_X1 U2754 ( .B1(n2222), .B2(n389), .A(n390), .ZN(n388) );
  AOI21_X1 U2755 ( .B1(n665), .B2(n483), .A(n472), .ZN(n468) );
  NAND2_X1 U2756 ( .A1(n666), .A2(n665), .ZN(n467) );
  OAI22_X1 U2757 ( .A1(n1941), .A2(n1691), .B1(n1690), .B2(n2268), .ZN(n1394)
         );
  OAI22_X1 U2758 ( .A1(n1941), .A2(n1686), .B1(n2267), .B2(n1685), .ZN(n1389)
         );
  OAI22_X1 U2759 ( .A1(n2247), .A2(n1689), .B1(n1688), .B2(n2267), .ZN(n1392)
         );
  OAI22_X1 U2760 ( .A1(n1941), .A2(n1690), .B1(n2268), .B2(n1689), .ZN(n1393)
         );
  OAI22_X1 U2761 ( .A1(n1941), .A2(n1687), .B1(n1686), .B2(n2268), .ZN(n1390)
         );
  OAI22_X1 U2762 ( .A1(n1941), .A2(n1692), .B1(n2267), .B2(n1691), .ZN(n1395)
         );
  OAI22_X1 U2763 ( .A1(n1941), .A2(n1685), .B1(n1684), .B2(n2267), .ZN(n1388)
         );
  OAI22_X1 U2764 ( .A1(n2247), .A2(n1688), .B1(n2268), .B2(n1687), .ZN(n1391)
         );
  OAI22_X1 U2765 ( .A1(n1955), .A2(n1684), .B1(n2267), .B2(n1683), .ZN(n1387)
         );
  OAI22_X1 U2766 ( .A1(n1941), .A2(n2311), .B1(n1706), .B2(n2267), .ZN(n1190)
         );
  OAI22_X1 U2767 ( .A1(n2247), .A2(n1693), .B1(n1692), .B2(n2268), .ZN(n1396)
         );
  XNOR2_X1 U2768 ( .A(b[13]), .B(n2314), .ZN(n1717) );
  XNOR2_X1 U2769 ( .A(b[21]), .B(n2313), .ZN(n1709) );
  XNOR2_X1 U2770 ( .A(b[15]), .B(n2314), .ZN(n1715) );
  XNOR2_X1 U2771 ( .A(b[11]), .B(n2314), .ZN(n1719) );
  XNOR2_X1 U2772 ( .A(b[19]), .B(n2313), .ZN(n1711) );
  XNOR2_X1 U2773 ( .A(b[17]), .B(n2313), .ZN(n1713) );
  INV_X1 U2774 ( .A(n1938), .ZN(n2262) );
  INV_X1 U2775 ( .A(n2197), .ZN(n2266) );
  INV_X1 U2776 ( .A(n2158), .ZN(n2270) );
  INV_X1 U2777 ( .A(n2281), .ZN(n2279) );
  INV_X1 U2778 ( .A(a[21]), .ZN(n2280) );
  INV_X1 U2779 ( .A(a[21]), .ZN(n2281) );
  INV_X1 U2780 ( .A(n2287), .ZN(n2285) );
  INV_X1 U2781 ( .A(a[19]), .ZN(n2286) );
  INV_X1 U2782 ( .A(a[19]), .ZN(n2287) );
  INV_X1 U2783 ( .A(n2292), .ZN(n2290) );
  INV_X1 U2784 ( .A(a[17]), .ZN(n2291) );
  INV_X1 U2785 ( .A(a[17]), .ZN(n2292) );
  INV_X1 U2786 ( .A(a[15]), .ZN(n2295) );
  INV_X1 U2787 ( .A(n2298), .ZN(n2297) );
  INV_X1 U2788 ( .A(a[13]), .ZN(n2298) );
  INV_X1 U2789 ( .A(n2303), .ZN(n2301) );
  INV_X1 U2790 ( .A(a[11]), .ZN(n2302) );
  INV_X1 U2791 ( .A(a[11]), .ZN(n2303) );
  INV_X1 U2792 ( .A(n2307), .ZN(n2305) );
  INV_X1 U2793 ( .A(a[9]), .ZN(n2306) );
  INV_X1 U2794 ( .A(a[9]), .ZN(n2307) );
  INV_X1 U2795 ( .A(a[7]), .ZN(n2311) );
  INV_X1 U2796 ( .A(a[7]), .ZN(n2312) );
  INV_X1 U2797 ( .A(n2316), .ZN(n2315) );
  INV_X1 U2798 ( .A(a[5]), .ZN(n2316) );
  INV_X1 U2799 ( .A(a[5]), .ZN(n2317) );
  INV_X1 U2800 ( .A(n2321), .ZN(n2320) );
  INV_X1 U2801 ( .A(a[3]), .ZN(n2321) );
  INV_X1 U2802 ( .A(n2325), .ZN(n2323) );
  INV_X1 U2803 ( .A(a[1]), .ZN(n2324) );
  INV_X1 U2804 ( .A(a[1]), .ZN(n2325) );
endmodule


module iir_filter_DW_mult_tc_1 ( a, b, product );
  input [23:0] a;
  input [23:0] b;
  output [47:0] product;
  wire   n251, n257, n277, n281, n287, n295, n297, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n325, n326, n327, n332, n333, n334,
         n335, n336, n337, n339, n341, n342, n344, n345, n346, n347, n348,
         n350, n352, n353, n354, n355, n356, n359, n360, n361, n362, n363,
         n364, n365, n367, n369, n370, n371, n372, n376, n378, n379, n380,
         n381, n382, n383, n384, n387, n388, n389, n390, n394, n396, n397,
         n398, n399, n400, n401, n402, n405, n407, n409, n410, n411, n412,
         n416, n418, n419, n420, n421, n422, n423, n426, n427, n428, n429,
         n430, n431, n432, n434, n435, n436, n437, n438, n439, n445, n451,
         n452, n453, n454, n455, n456, n457, n459, n461, n462, n463, n464,
         n465, n466, n467, n468, n474, n475, n476, n477, n478, n479, n480,
         n481, n483, n486, n487, n488, n489, n490, n492, n495, n496, n497,
         n498, n499, n501, n502, n503, n504, n505, n506, n507, n508, n511,
         n512, n513, n514, n515, n516, n517, n519, n520, n521, n522, n523,
         n524, n525, n526, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n550, n551,
         n552, n553, n554, n555, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n581, n582, n583,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n609, n610, n611, n620, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n643, n644,
         n645, n646, n657, n661, n662, n663, n666, n667, n668, n669, n670,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1806, n1807, n1810, n1811, n1814, n1817, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294;

  FA_X1 U546 ( .A(n1195), .B(n682), .CI(n1218), .CO(n678), .S(n679) );
  FA_X1 U547 ( .A(n683), .B(n1196), .CI(n686), .CO(n680), .S(n681) );
  FA_X1 U549 ( .A(n690), .B(n1242), .CI(n687), .CO(n684), .S(n685) );
  FA_X1 U550 ( .A(n1219), .B(n692), .CI(n1197), .CO(n686), .S(n687) );
  FA_X1 U551 ( .A(n691), .B(n698), .CI(n696), .CO(n688), .S(n689) );
  FA_X1 U552 ( .A(n1198), .B(n1220), .CI(n693), .CO(n690), .S(n691) );
  FA_X1 U554 ( .A(n702), .B(n699), .CI(n697), .CO(n694), .S(n695) );
  FA_X1 U555 ( .A(n1266), .B(n1243), .CI(n704), .CO(n696), .S(n697) );
  FA_X1 U556 ( .A(n1221), .B(n1199), .CI(n706), .CO(n698), .S(n699) );
  FA_X1 U557 ( .A(n710), .B(n712), .CI(n703), .CO(n700), .S(n701) );
  FA_X1 U558 ( .A(n714), .B(n1244), .CI(n705), .CO(n702), .S(n703) );
  FA_X1 U559 ( .A(n1222), .B(n1200), .CI(n707), .CO(n704), .S(n705) );
  FA_X1 U561 ( .A(n718), .B(n713), .CI(n711), .CO(n708), .S(n709) );
  FA_X1 U562 ( .A(n715), .B(n722), .CI(n720), .CO(n710), .S(n711) );
  FA_X1 U563 ( .A(n1245), .B(n1223), .CI(n1290), .CO(n712), .S(n713) );
  FA_X1 U564 ( .A(n1267), .B(n1201), .CI(n724), .CO(n714), .S(n715) );
  FA_X1 U565 ( .A(n728), .B(n721), .CI(n719), .CO(n716), .S(n717) );
  FA_X1 U566 ( .A(n723), .B(n732), .CI(n730), .CO(n718), .S(n719) );
  FA_X1 U567 ( .A(n1202), .B(n1246), .CI(n734), .CO(n720), .S(n721) );
  FA_X1 U568 ( .A(n1268), .B(n1224), .CI(n725), .CO(n722), .S(n723) );
  FA_X1 U570 ( .A(n738), .B(n731), .CI(n729), .CO(n726), .S(n727) );
  FA_X1 U571 ( .A(n735), .B(n733), .CI(n740), .CO(n728), .S(n729) );
  FA_X1 U572 ( .A(n744), .B(n1314), .CI(n742), .CO(n730), .S(n731) );
  FA_X1 U573 ( .A(n1225), .B(n1291), .CI(n1269), .CO(n732), .S(n733) );
  FA_X1 U574 ( .A(n746), .B(n1247), .CI(n1203), .CO(n734), .S(n735) );
  FA_X1 U575 ( .A(n750), .B(n741), .CI(n739), .CO(n736), .S(n737) );
  FA_X1 U576 ( .A(n754), .B(n745), .CI(n752), .CO(n738), .S(n739) );
  FA_X1 U577 ( .A(n756), .B(n758), .CI(n743), .CO(n740), .S(n741) );
  FA_X1 U578 ( .A(n1226), .B(n1204), .CI(n1270), .CO(n742), .S(n743) );
  FA_X1 U579 ( .A(n1292), .B(n1248), .CI(n747), .CO(n744), .S(n745) );
  FA_X1 U581 ( .A(n762), .B(n753), .CI(n751), .CO(n748), .S(n749) );
  FA_X1 U582 ( .A(n755), .B(n766), .CI(n764), .CO(n750), .S(n751) );
  FA_X1 U583 ( .A(n757), .B(n768), .CI(n759), .CO(n752), .S(n753) );
  FA_X1 U584 ( .A(n1338), .B(n1271), .CI(n770), .CO(n754), .S(n755) );
  FA_X1 U585 ( .A(n1249), .B(n1293), .CI(n1315), .CO(n756), .S(n757) );
  FA_X1 U586 ( .A(n772), .B(n1205), .CI(n1227), .CO(n758), .S(n759) );
  FA_X1 U587 ( .A(n776), .B(n765), .CI(n763), .CO(n760), .S(n761) );
  FA_X1 U588 ( .A(n767), .B(n780), .CI(n778), .CO(n762), .S(n763) );
  FA_X1 U589 ( .A(n771), .B(n769), .CI(n782), .CO(n764), .S(n765) );
  FA_X1 U590 ( .A(n786), .B(n1228), .CI(n784), .CO(n766), .S(n767) );
  FA_X1 U591 ( .A(n1294), .B(n1206), .CI(n1272), .CO(n768), .S(n769) );
  FA_X1 U592 ( .A(n1316), .B(n1250), .CI(n773), .CO(n770), .S(n771) );
  FA_X1 U594 ( .A(n790), .B(n779), .CI(n777), .CO(n774), .S(n775) );
  FA_X1 U595 ( .A(n781), .B(n794), .CI(n792), .CO(n776), .S(n777) );
  FA_X1 U596 ( .A(n783), .B(n787), .CI(n796), .CO(n778), .S(n779) );
  FA_X1 U597 ( .A(n798), .B(n800), .CI(n785), .CO(n780), .S(n781) );
  FA_X1 U598 ( .A(n1339), .B(n1229), .CI(n1362), .CO(n782), .S(n783) );
  FA_X1 U599 ( .A(n1273), .B(n1317), .CI(n1295), .CO(n784), .S(n785) );
  FA_X1 U600 ( .A(n802), .B(n1207), .CI(n1251), .CO(n786), .S(n787) );
  FA_X1 U601 ( .A(n806), .B(n793), .CI(n791), .CO(n788), .S(n789) );
  FA_X1 U603 ( .A(n797), .B(n801), .CI(n812), .CO(n792), .S(n793) );
  FA_X1 U604 ( .A(n814), .B(n816), .CI(n799), .CO(n794), .S(n795) );
  FA_X1 U606 ( .A(n1208), .B(n1318), .CI(n1230), .CO(n798), .S(n799) );
  FA_X1 U607 ( .A(n1340), .B(n1252), .CI(n803), .CO(n800), .S(n801) );
  FA_X1 U609 ( .A(n822), .B(n809), .CI(n807), .CO(n804), .S(n805) );
  FA_X1 U610 ( .A(n811), .B(n826), .CI(n824), .CO(n806), .S(n807) );
  FA_X1 U611 ( .A(n828), .B(n819), .CI(n813), .CO(n808), .S(n809) );
  FA_X1 U612 ( .A(n815), .B(n832), .CI(n817), .CO(n810), .S(n811) );
  FA_X1 U613 ( .A(n830), .B(n1386), .CI(n834), .CO(n812), .S(n813) );
  FA_X1 U614 ( .A(n1319), .B(n1253), .CI(n1341), .CO(n814), .S(n815) );
  FA_X1 U615 ( .A(n1231), .B(n1297), .CI(n1275), .CO(n816), .S(n817) );
  FA_X1 U616 ( .A(n2189), .B(n1209), .CI(n1363), .CO(n818), .S(n819) );
  FA_X1 U617 ( .A(n840), .B(n825), .CI(n823), .CO(n820), .S(n821) );
  FA_X1 U619 ( .A(n846), .B(n848), .CI(n829), .CO(n824), .S(n825) );
  FA_X1 U620 ( .A(n835), .B(n831), .CI(n833), .CO(n826), .S(n827) );
  FA_X1 U621 ( .A(n850), .B(n854), .CI(n852), .CO(n828), .S(n829) );
  FA_X1 U622 ( .A(n1254), .B(n1320), .CI(n1298), .CO(n830), .S(n831) );
  FA_X1 U623 ( .A(n1232), .B(n1364), .CI(n1342), .CO(n832), .S(n833) );
  FA_X1 U624 ( .A(n1276), .B(n1210), .CI(n837), .CO(n834), .S(n835) );
  FA_X1 U626 ( .A(n858), .B(n843), .CI(n841), .CO(n838), .S(n839) );
  FA_X1 U627 ( .A(n845), .B(n847), .CI(n860), .CO(n840), .S(n841) );
  FA_X1 U628 ( .A(n864), .B(n849), .CI(n862), .CO(n842), .S(n843) );
  FA_X1 U629 ( .A(n855), .B(n853), .CI(n866), .CO(n844), .S(n845) );
  FA_X1 U631 ( .A(n1410), .B(n1365), .CI(n872), .CO(n848), .S(n849) );
  FA_X1 U632 ( .A(n1343), .B(n1277), .CI(n1299), .CO(n850), .S(n851) );
  FA_X1 U633 ( .A(n1255), .B(n1321), .CI(n874), .CO(n852), .S(n853) );
  FA_X1 U634 ( .A(n1387), .B(n1233), .CI(n1211), .CO(n854), .S(n855) );
  FA_X1 U637 ( .A(n867), .B(n884), .CI(n865), .CO(n860), .S(n861) );
  FA_X1 U639 ( .A(n869), .B(n890), .CI(n871), .CO(n864), .S(n865) );
  FA_X1 U640 ( .A(n894), .B(n1300), .CI(n892), .CO(n866), .S(n867) );
  FA_X1 U641 ( .A(n1256), .B(n1234), .CI(n1322), .CO(n868), .S(n869) );
  FA_X1 U642 ( .A(n1344), .B(n1366), .CI(n1212), .CO(n870), .S(n871) );
  FA_X1 U643 ( .A(n1388), .B(n1278), .CI(n875), .CO(n872), .S(n873) );
  FA_X1 U645 ( .A(n898), .B(n881), .CI(n1937), .CO(n876), .S(n877) );
  FA_X1 U646 ( .A(n883), .B(n885), .CI(n900), .CO(n878), .S(n879) );
  FA_X1 U648 ( .A(n906), .B(n893), .CI(n889), .CO(n882), .S(n883) );
  FA_X1 U649 ( .A(n891), .B(n908), .CI(n895), .CO(n884), .S(n885) );
  FA_X1 U651 ( .A(n1367), .B(n1389), .CI(n1434), .CO(n888), .S(n889) );
  FA_X1 U652 ( .A(n1257), .B(n1345), .CI(n1301), .CO(n890), .S(n891) );
  FA_X1 U653 ( .A(n1279), .B(n1323), .CI(n2198), .CO(n892), .S(n893) );
  FA_X1 U654 ( .A(n1411), .B(n1235), .CI(n1213), .CO(n894), .S(n895) );
  FA_X1 U656 ( .A(n903), .B(n924), .CI(n922), .CO(n898), .S(n899) );
  FA_X1 U657 ( .A(n907), .B(n926), .CI(n905), .CO(n900), .S(n901) );
  FA_X1 U658 ( .A(n909), .B(n930), .CI(n928), .CO(n902), .S(n903) );
  FA_X1 U659 ( .A(n913), .B(n911), .CI(n915), .CO(n904), .S(n905) );
  FA_X1 U660 ( .A(n932), .B(n936), .CI(n934), .CO(n906), .S(n907) );
  FA_X1 U661 ( .A(n1368), .B(n1390), .CI(n938), .CO(n908), .S(n909) );
  FA_X1 U662 ( .A(n1324), .B(n1346), .CI(n1280), .CO(n910), .S(n911) );
  FA_X1 U663 ( .A(n1412), .B(n1258), .CI(n1236), .CO(n912), .S(n913) );
  FA_X1 U664 ( .A(n1302), .B(n1214), .CI(n917), .CO(n914), .S(n915) );
  FA_X1 U667 ( .A(n925), .B(n927), .CI(n944), .CO(n920), .S(n921) );
  FA_X1 U668 ( .A(n929), .B(n948), .CI(n946), .CO(n922), .S(n923) );
  FA_X1 U669 ( .A(n950), .B(n935), .CI(n931), .CO(n924), .S(n925) );
  FA_X1 U670 ( .A(n937), .B(n933), .CI(n952), .CO(n926), .S(n927) );
  FA_X1 U671 ( .A(n954), .B(n958), .CI(n956), .CO(n928), .S(n929) );
  FA_X1 U672 ( .A(n1458), .B(n960), .CI(n939), .CO(n930), .S(n931) );
  FA_X1 U673 ( .A(n1325), .B(n1413), .CI(n1435), .CO(n932), .S(n933) );
  FA_X1 U674 ( .A(n1281), .B(n1369), .CI(n1391), .CO(n934), .S(n935) );
  FA_X1 U675 ( .A(n1303), .B(n1347), .CI(n1259), .CO(n936), .S(n937) );
  FA_X1 U678 ( .A(n964), .B(n945), .CI(n943), .CO(n940), .S(n941) );
  FA_X1 U679 ( .A(n947), .B(n949), .CI(n966), .CO(n942), .S(n943) );
  FA_X1 U680 ( .A(n951), .B(n970), .CI(n968), .CO(n944), .S(n945) );
  FA_X1 U682 ( .A(n955), .B(n974), .CI(n957), .CO(n948), .S(n949) );
  FA_X1 U683 ( .A(n976), .B(n980), .CI(n978), .CO(n950), .S(n951) );
  FA_X1 U685 ( .A(n1282), .B(n1414), .CI(n1304), .CO(n954), .S(n955) );
  FA_X1 U686 ( .A(n1459), .B(n1370), .CI(n1436), .CO(n956), .S(n957) );
  FA_X1 U687 ( .A(n1260), .B(n1182), .CI(n1348), .CO(n958), .S(n959) );
  HA_X1 U688 ( .A(n1216), .B(n1238), .CO(n960), .S(n961) );
  FA_X1 U689 ( .A(n984), .B(n967), .CI(n965), .CO(n962), .S(n963) );
  FA_X1 U690 ( .A(n969), .B(n971), .CI(n986), .CO(n964), .S(n965) );
  FA_X1 U691 ( .A(n973), .B(n990), .CI(n988), .CO(n966), .S(n967) );
  FA_X1 U692 ( .A(n975), .B(n981), .CI(n992), .CO(n968), .S(n969) );
  FA_X1 U693 ( .A(n977), .B(n998), .CI(n979), .CO(n970), .S(n971) );
  FA_X1 U695 ( .A(n1393), .B(n1415), .CI(n1000), .CO(n974), .S(n975) );
  FA_X1 U696 ( .A(n1305), .B(n1437), .CI(n1327), .CO(n976), .S(n977) );
  FA_X1 U697 ( .A(n1460), .B(n1371), .CI(n1283), .CO(n978), .S(n979) );
  FA_X1 U698 ( .A(n1239), .B(n1349), .CI(n1261), .CO(n980), .S(n981) );
  FA_X1 U699 ( .A(n1004), .B(n987), .CI(n985), .CO(n982), .S(n983) );
  FA_X1 U700 ( .A(n989), .B(n991), .CI(n1006), .CO(n984), .S(n985) );
  FA_X1 U701 ( .A(n993), .B(n1010), .CI(n1008), .CO(n986), .S(n987) );
  FA_X1 U702 ( .A(n999), .B(n997), .CI(n1012), .CO(n988), .S(n989) );
  FA_X1 U703 ( .A(n1014), .B(n1016), .CI(n995), .CO(n990), .S(n991) );
  FA_X1 U704 ( .A(n1001), .B(n1394), .CI(n1018), .CO(n992), .S(n993) );
  FA_X1 U707 ( .A(n1461), .B(n1350), .CI(n1183), .CO(n998), .S(n999) );
  HA_X1 U708 ( .A(n1240), .B(n1262), .CO(n1000), .S(n1001) );
  FA_X1 U709 ( .A(n1022), .B(n1007), .CI(n1005), .CO(n1002), .S(n1003) );
  FA_X1 U710 ( .A(n1009), .B(n1011), .CI(n1024), .CO(n1004), .S(n1005) );
  FA_X1 U711 ( .A(n1013), .B(n1028), .CI(n1026), .CO(n1006), .S(n1007) );
  FA_X1 U712 ( .A(n1019), .B(n1015), .CI(n1017), .CO(n1008), .S(n1009) );
  FA_X1 U713 ( .A(n1030), .B(n1034), .CI(n1241), .CO(n1010), .S(n1011) );
  FA_X1 U714 ( .A(n1036), .B(n1439), .CI(n1032), .CO(n1012), .S(n1013) );
  FA_X1 U715 ( .A(n1395), .B(n1462), .CI(n1417), .CO(n1014), .S(n1015) );
  FA_X1 U716 ( .A(n1307), .B(n1373), .CI(n1329), .CO(n1016), .S(n1017) );
  FA_X1 U717 ( .A(n1263), .B(n1351), .CI(n1285), .CO(n1018), .S(n1019) );
  FA_X1 U719 ( .A(n1027), .B(n1044), .CI(n1042), .CO(n1022), .S(n1023) );
  FA_X1 U720 ( .A(n1046), .B(n1035), .CI(n1029), .CO(n1024), .S(n1025) );
  FA_X1 U721 ( .A(n1031), .B(n1048), .CI(n1033), .CO(n1026), .S(n1027) );
  FA_X1 U722 ( .A(n1052), .B(n1037), .CI(n1050), .CO(n1028), .S(n1029) );
  FA_X1 U723 ( .A(n1352), .B(n1440), .CI(n1418), .CO(n1030), .S(n1031) );
  FA_X1 U724 ( .A(n1463), .B(n1330), .CI(n1396), .CO(n1032), .S(n1033) );
  FA_X1 U725 ( .A(n1184), .B(n1374), .CI(n1308), .CO(n1034), .S(n1035) );
  HA_X1 U726 ( .A(n1264), .B(n1286), .CO(n1036), .S(n1037) );
  FA_X1 U727 ( .A(n1056), .B(n1043), .CI(n1041), .CO(n1038), .S(n1039) );
  FA_X1 U728 ( .A(n1058), .B(n1047), .CI(n1045), .CO(n1040), .S(n1041) );
  FA_X1 U729 ( .A(n1062), .B(n1053), .CI(n1060), .CO(n1042), .S(n1043) );
  FA_X1 U730 ( .A(n1049), .B(n1265), .CI(n1051), .CO(n1044), .S(n1045) );
  FA_X1 U731 ( .A(n1064), .B(n1068), .CI(n1066), .CO(n1046), .S(n1047) );
  FA_X1 U732 ( .A(n1397), .B(n1419), .CI(n1441), .CO(n1048), .S(n1049) );
  FA_X1 U733 ( .A(n1331), .B(n1353), .CI(n1375), .CO(n1050), .S(n1051) );
  FA_X1 U734 ( .A(n1287), .B(n1464), .CI(n1309), .CO(n1052), .S(n1053) );
  FA_X1 U735 ( .A(n1072), .B(n1059), .CI(n1057), .CO(n1054), .S(n1055) );
  FA_X1 U736 ( .A(n1074), .B(n1063), .CI(n1061), .CO(n1056), .S(n1057) );
  FA_X1 U737 ( .A(n1067), .B(n1065), .CI(n1076), .CO(n1058), .S(n1059) );
  FA_X1 U738 ( .A(n1080), .B(n1082), .CI(n1078), .CO(n1060), .S(n1061) );
  FA_X1 U739 ( .A(n1398), .B(n1420), .CI(n1069), .CO(n1062), .S(n1063) );
  FA_X1 U740 ( .A(n1442), .B(n1354), .CI(n1332), .CO(n1064), .S(n1065) );
  FA_X1 U741 ( .A(n1465), .B(n1376), .CI(n1185), .CO(n1066), .S(n1067) );
  HA_X1 U742 ( .A(n1288), .B(n1310), .CO(n1068), .S(n1069) );
  FA_X1 U743 ( .A(n1086), .B(n1075), .CI(n1073), .CO(n1070), .S(n1071) );
  FA_X1 U744 ( .A(n1088), .B(n1090), .CI(n1077), .CO(n1072), .S(n1073) );
  FA_X1 U745 ( .A(n1083), .B(n1081), .CI(n1079), .CO(n1074), .S(n1075) );
  FA_X1 U746 ( .A(n1289), .B(n1094), .CI(n1092), .CO(n1076), .S(n1077) );
  FA_X1 U747 ( .A(n1399), .B(n1421), .CI(n1096), .CO(n1078), .S(n1079) );
  FA_X1 U748 ( .A(n1355), .B(n1443), .CI(n1377), .CO(n1080), .S(n1081) );
  FA_X1 U749 ( .A(n1311), .B(n1466), .CI(n1333), .CO(n1082), .S(n1083) );
  FA_X1 U750 ( .A(n1100), .B(n1089), .CI(n1087), .CO(n1084), .S(n1085) );
  FA_X1 U751 ( .A(n1102), .B(n1104), .CI(n1091), .CO(n1086), .S(n1087) );
  FA_X1 U752 ( .A(n1093), .B(n1106), .CI(n1095), .CO(n1088), .S(n1089) );
  FA_X1 U753 ( .A(n1097), .B(n1422), .CI(n1108), .CO(n1090), .S(n1091) );
  FA_X1 U754 ( .A(n1356), .B(n1444), .CI(n1378), .CO(n1092), .S(n1093) );
  FA_X1 U755 ( .A(n1467), .B(n1400), .CI(n1186), .CO(n1094), .S(n1095) );
  HA_X1 U756 ( .A(n1334), .B(n1312), .CO(n1096), .S(n1097) );
  FA_X1 U757 ( .A(n1103), .B(n1112), .CI(n1101), .CO(n1098), .S(n1099) );
  FA_X1 U758 ( .A(n1114), .B(n1109), .CI(n1105), .CO(n1100), .S(n1101) );
  FA_X1 U759 ( .A(n1313), .B(n1116), .CI(n1107), .CO(n1102), .S(n1103) );
  FA_X1 U760 ( .A(n1120), .B(n1423), .CI(n1118), .CO(n1104), .S(n1105) );
  FA_X1 U761 ( .A(n1379), .B(n1445), .CI(n1401), .CO(n1106), .S(n1107) );
  FA_X1 U762 ( .A(n1335), .B(n1468), .CI(n1357), .CO(n1108), .S(n1109) );
  FA_X1 U763 ( .A(n1124), .B(n1115), .CI(n1113), .CO(n1110), .S(n1111) );
  FA_X1 U764 ( .A(n1119), .B(n1117), .CI(n1126), .CO(n1112), .S(n1113) );
  FA_X1 U765 ( .A(n1130), .B(n1121), .CI(n1128), .CO(n1114), .S(n1115) );
  FA_X1 U766 ( .A(n1424), .B(n1469), .CI(n1446), .CO(n1116), .S(n1117) );
  FA_X1 U767 ( .A(n1380), .B(n1402), .CI(n1187), .CO(n1118), .S(n1119) );
  HA_X1 U768 ( .A(n1336), .B(n1358), .CO(n1120), .S(n1121) );
  FA_X1 U769 ( .A(n1127), .B(n1134), .CI(n1125), .CO(n1122), .S(n1123) );
  FA_X1 U770 ( .A(n1131), .B(n1129), .CI(n1136), .CO(n1124), .S(n1125) );
  FA_X1 U771 ( .A(n1138), .B(n1140), .CI(n1337), .CO(n1126), .S(n1127) );
  FA_X1 U772 ( .A(n1403), .B(n1447), .CI(n1425), .CO(n1128), .S(n1129) );
  FA_X1 U773 ( .A(n1359), .B(n1470), .CI(n1381), .CO(n1130), .S(n1131) );
  FA_X1 U774 ( .A(n1144), .B(n1137), .CI(n1135), .CO(n1132), .S(n1133) );
  FA_X1 U775 ( .A(n1146), .B(n1148), .CI(n1139), .CO(n1134), .S(n1135) );
  FA_X1 U776 ( .A(n1404), .B(n1448), .CI(n1141), .CO(n1136), .S(n1137) );
  FA_X1 U777 ( .A(n1471), .B(n1426), .CI(n1188), .CO(n1138), .S(n1139) );
  HA_X1 U778 ( .A(n1360), .B(n1382), .CO(n1140), .S(n1141) );
  FA_X1 U779 ( .A(n1152), .B(n1147), .CI(n1145), .CO(n1142), .S(n1143) );
  FA_X1 U780 ( .A(n1361), .B(n1154), .CI(n1149), .CO(n1144), .S(n1145) );
  FA_X1 U781 ( .A(n1427), .B(n1449), .CI(n1156), .CO(n1146), .S(n1147) );
  FA_X1 U782 ( .A(n1383), .B(n1472), .CI(n1405), .CO(n1148), .S(n1149) );
  FA_X1 U783 ( .A(n1160), .B(n1155), .CI(n1153), .CO(n1150), .S(n1151) );
  FA_X1 U784 ( .A(n1157), .B(n1473), .CI(n1162), .CO(n1152), .S(n1153) );
  FA_X1 U785 ( .A(n1450), .B(n1428), .CI(n1189), .CO(n1154), .S(n1155) );
  HA_X1 U786 ( .A(n1384), .B(n1406), .CO(n1156), .S(n1157) );
  FA_X1 U787 ( .A(n1163), .B(n1385), .CI(n1164), .CO(n1158), .S(n1159) );
  FA_X1 U788 ( .A(n1168), .B(n1429), .CI(n1166), .CO(n1160), .S(n1161) );
  FA_X1 U789 ( .A(n1451), .B(n1474), .CI(n1407), .CO(n1162), .S(n1163) );
  FA_X1 U790 ( .A(n1172), .B(n1169), .CI(n1167), .CO(n1164), .S(n1165) );
  FA_X1 U791 ( .A(n1452), .B(n1475), .CI(n1190), .CO(n1166), .S(n1167) );
  HA_X1 U792 ( .A(n1408), .B(n1430), .CO(n1168), .S(n1169) );
  FA_X1 U793 ( .A(n1409), .B(n1176), .CI(n1173), .CO(n1170), .S(n1171) );
  FA_X1 U794 ( .A(n1476), .B(n1453), .CI(n1431), .CO(n1172), .S(n1173) );
  FA_X1 U795 ( .A(n1191), .B(n1454), .CI(n1177), .CO(n1174), .S(n1175) );
  HA_X1 U796 ( .A(n1432), .B(n1477), .CO(n1176), .S(n1177) );
  FA_X1 U797 ( .A(n1455), .B(n1478), .CI(n1180), .CO(n1178), .S(n1179) );
  HA_X1 U798 ( .A(n1456), .B(n1479), .CO(n1180), .S(n1181) );
  OR2_X2 U1448 ( .A1(n2134), .A2(n2128), .ZN(n1929) );
  OR2_X1 U1449 ( .A1(n2134), .A2(n2128), .ZN(n1987) );
  INV_X1 U1450 ( .A(n2128), .ZN(n2222) );
  CLKBUF_X1 U1451 ( .A(n287), .Z(n2180) );
  BUF_X1 U1452 ( .A(n550), .Z(n1930) );
  OAI21_X1 U1453 ( .B1(n535), .B2(n2071), .A(n2050), .ZN(n1931) );
  CLKBUF_X1 U1454 ( .A(n532), .Z(n2050) );
  CLKBUF_X1 U1455 ( .A(n552), .Z(n1932) );
  BUF_X1 U1456 ( .A(n1284), .Z(n1933) );
  XNOR2_X1 U1457 ( .A(n1934), .B(n994), .ZN(n973) );
  XNOR2_X1 U1458 ( .A(n996), .B(n1217), .ZN(n1934) );
  BUF_X1 U1459 ( .A(n2022), .Z(n2146) );
  INV_X1 U1460 ( .A(n2251), .ZN(n2249) );
  INV_X1 U1461 ( .A(n2135), .ZN(n2004) );
  CLKBUF_X1 U1462 ( .A(a[16]), .Z(n1935) );
  INV_X1 U1463 ( .A(a[1]), .ZN(n1936) );
  FA_X1 U1464 ( .A(n883), .B(n885), .CI(n900), .S(n1937) );
  XOR2_X1 U1465 ( .A(n870), .B(n868), .Z(n1938) );
  XOR2_X1 U1466 ( .A(n851), .B(n1938), .Z(n847) );
  NAND2_X1 U1467 ( .A1(n851), .A2(n870), .ZN(n1939) );
  NAND2_X1 U1468 ( .A1(n851), .A2(n868), .ZN(n1940) );
  NAND2_X1 U1469 ( .A1(n870), .A2(n868), .ZN(n1941) );
  NAND3_X1 U1470 ( .A1(n1939), .A2(n1940), .A3(n1941), .ZN(n846) );
  INV_X2 U1471 ( .A(n1968), .ZN(n2238) );
  INV_X2 U1472 ( .A(n2244), .ZN(n2241) );
  INV_X2 U1473 ( .A(n2126), .ZN(n2169) );
  INV_X1 U1474 ( .A(n2175), .ZN(n1942) );
  OR2_X1 U1475 ( .A1(n1614), .A2(n1999), .ZN(n1943) );
  OR2_X1 U1476 ( .A1(n1613), .A2(n2143), .ZN(n1944) );
  NAND2_X1 U1477 ( .A1(n1943), .A2(n1944), .ZN(n1320) );
  INV_X1 U1478 ( .A(n2175), .ZN(n2225) );
  BUF_X2 U1479 ( .A(n2091), .Z(n2142) );
  CLKBUF_X3 U1480 ( .A(n281), .Z(n2193) );
  XNOR2_X1 U1481 ( .A(a[8]), .B(a[7]), .ZN(n2093) );
  INV_X1 U1482 ( .A(a[19]), .ZN(n1946) );
  INV_X1 U1483 ( .A(a[19]), .ZN(n1945) );
  INV_X1 U1484 ( .A(n2032), .ZN(n2192) );
  INV_X1 U1485 ( .A(n2137), .ZN(n2069) );
  NOR2_X1 U1486 ( .A1(n821), .A2(n838), .ZN(n502) );
  OAI21_X1 U1487 ( .B1(n572), .B2(n569), .A(n570), .ZN(n568) );
  OR2_X1 U1488 ( .A1(n709), .A2(n716), .ZN(n2115) );
  AND2_X1 U1489 ( .A1(n1193), .A2(n1481), .ZN(n1947) );
  OR2_X1 U1490 ( .A1(n1457), .A2(n1480), .ZN(n1948) );
  OR2_X1 U1491 ( .A1(n1179), .A2(n1433), .ZN(n1949) );
  AND2_X1 U1492 ( .A1(n1123), .A2(n1132), .ZN(n1950) );
  AND2_X1 U1493 ( .A1(n1143), .A2(n1150), .ZN(n1951) );
  AND2_X1 U1494 ( .A1(n1151), .A2(n1158), .ZN(n1952) );
  OR2_X1 U1495 ( .A1(n694), .A2(n689), .ZN(n1953) );
  AND2_X1 U1496 ( .A1(n1457), .A2(n1480), .ZN(n1954) );
  AND2_X1 U1497 ( .A1(n1179), .A2(n1433), .ZN(n1955) );
  AND2_X1 U1498 ( .A1(n1039), .A2(n1054), .ZN(n1956) );
  AND2_X1 U1499 ( .A1(n1111), .A2(n1122), .ZN(n1957) );
  AND2_X1 U1500 ( .A1(n1133), .A2(n1142), .ZN(n1958) );
  AND2_X1 U1501 ( .A1(n1055), .A2(n1070), .ZN(n1959) );
  OR2_X1 U1502 ( .A1(n1151), .A2(n1158), .ZN(n1960) );
  XNOR2_X1 U1503 ( .A(n551), .B(n1961), .ZN(product[23]) );
  AND2_X1 U1504 ( .A1(n674), .A2(n1930), .ZN(n1961) );
  XNOR2_X1 U1505 ( .A(n560), .B(n1962), .ZN(product[22]) );
  AND2_X1 U1506 ( .A1(n675), .A2(n559), .ZN(n1962) );
  XNOR2_X1 U1507 ( .A(n544), .B(n1963), .ZN(product[24]) );
  AND2_X1 U1508 ( .A1(n673), .A2(n543), .ZN(n1963) );
  CLKBUF_X1 U1509 ( .A(n2224), .Z(n1964) );
  CLKBUF_X3 U1510 ( .A(n2224), .Z(n1965) );
  INV_X1 U1511 ( .A(n2158), .ZN(n2224) );
  XNOR2_X1 U1512 ( .A(n2007), .B(n1966), .ZN(product[34]) );
  AND2_X1 U1513 ( .A1(n663), .A2(n439), .ZN(n1966) );
  BUF_X2 U1514 ( .A(n2246), .Z(n1997) );
  BUF_X1 U1515 ( .A(n2202), .Z(n2007) );
  INV_X2 U1516 ( .A(n2255), .ZN(n2254) );
  AND2_X1 U1517 ( .A1(n2106), .A2(n2022), .ZN(n2136) );
  INV_X1 U1518 ( .A(n2022), .ZN(n2178) );
  INV_X1 U1519 ( .A(n2264), .ZN(n1967) );
  INV_X1 U1520 ( .A(a[21]), .ZN(n1968) );
  XNOR2_X1 U1521 ( .A(a[10]), .B(n2016), .ZN(n2106) );
  CLKBUF_X1 U1522 ( .A(n902), .Z(n1969) );
  CLKBUF_X1 U1523 ( .A(n2142), .Z(n1970) );
  CLKBUF_X1 U1524 ( .A(n2173), .Z(n1971) );
  BUF_X2 U1525 ( .A(n2173), .Z(n1973) );
  CLKBUF_X3 U1526 ( .A(n2173), .Z(n1972) );
  BUF_X1 U1527 ( .A(n297), .Z(n2173) );
  INV_X1 U1528 ( .A(n2158), .ZN(n1974) );
  INV_X1 U1529 ( .A(n2013), .ZN(n2158) );
  XNOR2_X1 U1530 ( .A(n1975), .B(n1985), .ZN(n995) );
  XNOR2_X1 U1531 ( .A(n1416), .B(n1328), .ZN(n1975) );
  INV_X1 U1532 ( .A(n2251), .ZN(n1977) );
  INV_X1 U1533 ( .A(n2251), .ZN(n1976) );
  XNOR2_X1 U1534 ( .A(n1978), .B(n953), .ZN(n947) );
  XNOR2_X1 U1535 ( .A(n972), .B(n959), .ZN(n1978) );
  AOI21_X1 U1536 ( .B1(n581), .B2(n567), .A(n568), .ZN(n1980) );
  AOI21_X1 U1537 ( .B1(n581), .B2(n567), .A(n568), .ZN(n1979) );
  AOI21_X1 U1538 ( .B1(n581), .B2(n567), .A(n568), .ZN(n566) );
  BUF_X2 U1539 ( .A(n2145), .Z(n1981) );
  XNOR2_X1 U1540 ( .A(a[14]), .B(n2251), .ZN(n1810) );
  NOR2_X1 U1541 ( .A1(n513), .A2(n520), .ZN(n1982) );
  INV_X1 U1542 ( .A(b[0]), .ZN(n1984) );
  INV_X1 U1543 ( .A(b[0]), .ZN(n1983) );
  INV_X1 U1544 ( .A(b[0]), .ZN(n2282) );
  BUF_X1 U1545 ( .A(n1306), .Z(n1985) );
  INV_X2 U1546 ( .A(n2127), .ZN(n1986) );
  INV_X1 U1547 ( .A(n2127), .ZN(n2221) );
  OR2_X1 U1548 ( .A1(n2134), .A2(n2128), .ZN(n2040) );
  CLKBUF_X1 U1549 ( .A(n2255), .Z(n1988) );
  INV_X2 U1550 ( .A(n2126), .ZN(n2209) );
  INV_X1 U1551 ( .A(n2259), .ZN(n1990) );
  INV_X1 U1552 ( .A(n2259), .ZN(n1989) );
  NOR2_X1 U1553 ( .A1(n505), .A2(n452), .ZN(n2188) );
  BUF_X1 U1554 ( .A(n536), .Z(n1991) );
  BUF_X1 U1555 ( .A(n536), .Z(n1993) );
  BUF_X1 U1556 ( .A(n536), .Z(n1992) );
  INV_X1 U1557 ( .A(n2048), .ZN(n1994) );
  INV_X1 U1558 ( .A(n1976), .ZN(n1995) );
  CLKBUF_X1 U1559 ( .A(n2246), .Z(n1996) );
  BUF_X2 U1560 ( .A(n2246), .Z(n1998) );
  INV_X1 U1561 ( .A(n2136), .ZN(n2015) );
  NAND2_X2 U1562 ( .A1(n1811), .A2(n2142), .ZN(n1999) );
  CLKBUF_X1 U1563 ( .A(n2013), .Z(n2000) );
  INV_X1 U1564 ( .A(n2030), .ZN(n2127) );
  XOR2_X1 U1565 ( .A(a[6]), .B(a[7]), .Z(n1814) );
  XOR2_X1 U1566 ( .A(a[2]), .B(a[1]), .Z(n2129) );
  INV_X1 U1567 ( .A(a[1]), .ZN(n2281) );
  INV_X1 U1568 ( .A(n2039), .ZN(n2001) );
  XNOR2_X1 U1569 ( .A(a[20]), .B(a[19]), .ZN(n2095) );
  BUF_X2 U1570 ( .A(n2229), .Z(n2002) );
  INV_X1 U1571 ( .A(n2230), .ZN(n2229) );
  INV_X1 U1572 ( .A(n2135), .ZN(n2003) );
  INV_X1 U1573 ( .A(n2135), .ZN(n2211) );
  BUF_X1 U1574 ( .A(n251), .Z(n2006) );
  CLKBUF_X3 U1575 ( .A(n251), .Z(n2005) );
  CLKBUF_X1 U1576 ( .A(n251), .Z(n2234) );
  XNOR2_X1 U1577 ( .A(a[22]), .B(n2237), .ZN(n1806) );
  BUF_X2 U1578 ( .A(n2225), .Z(n2143) );
  FA_X1 U1579 ( .A(n898), .B(n881), .CI(n879), .S(n2008) );
  INV_X1 U1580 ( .A(n2223), .ZN(n2009) );
  AND2_X2 U1581 ( .A1(n2010), .A2(n2012), .ZN(n2126) );
  XNOR2_X1 U1582 ( .A(a[18]), .B(n1946), .ZN(n2010) );
  CLKBUF_X3 U1583 ( .A(n2095), .Z(n2038) );
  INV_X1 U1584 ( .A(n2275), .ZN(n2011) );
  INV_X2 U1585 ( .A(n2277), .ZN(n2275) );
  INV_X2 U1586 ( .A(n2230), .ZN(n2228) );
  XNOR2_X1 U1587 ( .A(a[18]), .B(a[17]), .ZN(n2012) );
  INV_X2 U1588 ( .A(n2086), .ZN(n2089) );
  XNOR2_X1 U1589 ( .A(a[14]), .B(a[13]), .ZN(n2013) );
  AND2_X1 U1590 ( .A1(n775), .A2(n788), .ZN(n2036) );
  INV_X1 U1591 ( .A(n2269), .ZN(n2265) );
  NOR2_X1 U1592 ( .A1(n897), .A2(n918), .ZN(n534) );
  INV_X1 U1593 ( .A(n2036), .ZN(n474) );
  INV_X1 U1594 ( .A(n2136), .ZN(n2014) );
  INV_X1 U1595 ( .A(a[11]), .ZN(n2016) );
  OR2_X1 U1596 ( .A1(n2213), .A2(n1642), .ZN(n2017) );
  OR2_X1 U1597 ( .A1(n2226), .A2(n1641), .ZN(n2018) );
  NAND2_X1 U1598 ( .A1(n2017), .A2(n2018), .ZN(n1347) );
  INV_X1 U1599 ( .A(n2136), .ZN(n2213) );
  BUF_X2 U1600 ( .A(n287), .Z(n2177) );
  NOR2_X1 U1601 ( .A1(n941), .A2(n962), .ZN(n2019) );
  NOR2_X1 U1602 ( .A1(n962), .A2(n941), .ZN(n547) );
  INV_X1 U1603 ( .A(n2251), .ZN(n2250) );
  OR2_X2 U1604 ( .A1(n775), .A2(n788), .ZN(n2034) );
  NOR2_X2 U1605 ( .A1(n963), .A2(n982), .ZN(n558) );
  INV_X1 U1606 ( .A(n2259), .ZN(n2256) );
  CLKBUF_X1 U1607 ( .A(n2093), .Z(n2145) );
  CLKBUF_X1 U1608 ( .A(n2008), .Z(n2020) );
  XNOR2_X1 U1609 ( .A(a[0]), .B(n2281), .ZN(n1817) );
  XOR2_X1 U1610 ( .A(a[8]), .B(n2264), .Z(n2131) );
  INV_X1 U1611 ( .A(n2264), .ZN(n2261) );
  BUF_X4 U1612 ( .A(a[23]), .Z(n2021) );
  CLKBUF_X1 U1613 ( .A(n2155), .Z(n2071) );
  XNOR2_X1 U1614 ( .A(a[10]), .B(a[9]), .ZN(n2022) );
  INV_X2 U1615 ( .A(n2178), .ZN(n2226) );
  XOR2_X1 U1616 ( .A(n1326), .B(n1392), .Z(n2023) );
  XOR2_X1 U1617 ( .A(n2023), .B(n961), .Z(n953) );
  NAND2_X1 U1618 ( .A1(n1326), .A2(n1392), .ZN(n2024) );
  NAND2_X1 U1619 ( .A1(n1326), .A2(n961), .ZN(n2025) );
  NAND2_X1 U1620 ( .A1(n1392), .A2(n961), .ZN(n2026) );
  NAND3_X1 U1621 ( .A1(n2024), .A2(n2025), .A3(n2026), .ZN(n952) );
  NAND2_X1 U1622 ( .A1(n972), .A2(n959), .ZN(n2027) );
  NAND2_X1 U1623 ( .A1(n972), .A2(n953), .ZN(n2028) );
  NAND2_X1 U1624 ( .A1(n959), .A2(n953), .ZN(n2029) );
  NAND3_X1 U1625 ( .A1(n2027), .A2(n2028), .A3(n2029), .ZN(n946) );
  XNOR2_X1 U1626 ( .A(a[22]), .B(a[21]), .ZN(n2030) );
  CLKBUF_X1 U1627 ( .A(n1215), .Z(n2035) );
  XNOR2_X1 U1628 ( .A(a[20]), .B(n2240), .ZN(n1807) );
  NAND3_X1 U1629 ( .A1(n2073), .A2(n2074), .A3(n2075), .ZN(n2031) );
  XNOR2_X1 U1630 ( .A(a[4]), .B(a[3]), .ZN(n2032) );
  INV_X2 U1631 ( .A(n2192), .ZN(n2231) );
  CLKBUF_X3 U1632 ( .A(n2032), .Z(n2141) );
  NOR2_X1 U1633 ( .A1(n542), .A2(n547), .ZN(n2033) );
  AND2_X2 U1634 ( .A1(n1817), .A2(n2234), .ZN(n2138) );
  INV_X2 U1635 ( .A(n2137), .ZN(n2217) );
  INV_X1 U1636 ( .A(n2091), .ZN(n2175) );
  XOR2_X1 U1637 ( .A(a[15]), .B(a[16]), .Z(n2128) );
  INV_X1 U1638 ( .A(n2186), .ZN(n2037) );
  XOR2_X1 U1639 ( .A(n1935), .B(n2248), .Z(n2134) );
  INV_X1 U1640 ( .A(n1929), .ZN(n2133) );
  INV_X1 U1641 ( .A(n2126), .ZN(n2208) );
  INV_X2 U1642 ( .A(n2138), .ZN(n2219) );
  INV_X1 U1643 ( .A(n2093), .ZN(n2186) );
  XOR2_X1 U1644 ( .A(a[20]), .B(a[19]), .Z(n2039) );
  NAND2_X1 U1645 ( .A1(n1416), .A2(n1328), .ZN(n2041) );
  NAND2_X1 U1646 ( .A1(n1416), .A2(n1306), .ZN(n2042) );
  NAND2_X1 U1647 ( .A1(n1328), .A2(n1306), .ZN(n2043) );
  NAND3_X1 U1648 ( .A1(n2041), .A2(n2042), .A3(n2043), .ZN(n994) );
  NAND2_X1 U1649 ( .A1(n996), .A2(n1217), .ZN(n2044) );
  NAND2_X1 U1650 ( .A1(n996), .A2(n994), .ZN(n2045) );
  NAND2_X1 U1651 ( .A1(n1217), .A2(n994), .ZN(n2046) );
  NAND3_X1 U1652 ( .A1(n2044), .A2(n2045), .A3(n2046), .ZN(n972) );
  INV_X1 U1653 ( .A(n2137), .ZN(n2216) );
  INV_X1 U1654 ( .A(n2232), .ZN(n2047) );
  INV_X1 U1655 ( .A(n2047), .ZN(n2048) );
  INV_X2 U1656 ( .A(n2047), .ZN(n2049) );
  AOI21_X1 U1657 ( .B1(n540), .B2(n553), .A(n541), .ZN(n2051) );
  NOR2_X1 U1658 ( .A1(n531), .A2(n534), .ZN(n2052) );
  NOR2_X1 U1659 ( .A1(n531), .A2(n534), .ZN(n525) );
  INV_X1 U1660 ( .A(n2218), .ZN(n2190) );
  INV_X1 U1661 ( .A(n555), .ZN(n2053) );
  INV_X2 U1662 ( .A(n2138), .ZN(n2220) );
  OAI21_X1 U1663 ( .B1(n538), .B2(n1979), .A(n539), .ZN(n2054) );
  INV_X1 U1664 ( .A(n2096), .ZN(n2055) );
  OR2_X1 U1665 ( .A1(n2214), .A2(n1683), .ZN(n2056) );
  OR2_X1 U1666 ( .A1(n1682), .A2(n2229), .ZN(n2057) );
  NAND2_X1 U1667 ( .A1(n2056), .A2(n2057), .ZN(n836) );
  BUF_X1 U1668 ( .A(n836), .Z(n2189) );
  XOR2_X1 U1669 ( .A(n844), .B(n827), .Z(n2058) );
  XOR2_X1 U1670 ( .A(n842), .B(n2058), .Z(n823) );
  NAND2_X1 U1671 ( .A1(n842), .A2(n844), .ZN(n2059) );
  NAND2_X1 U1672 ( .A1(n842), .A2(n827), .ZN(n2060) );
  NAND2_X1 U1673 ( .A1(n844), .A2(n827), .ZN(n2061) );
  NAND3_X1 U1674 ( .A1(n2059), .A2(n2060), .A3(n2061), .ZN(n822) );
  OR2_X2 U1675 ( .A1(n2131), .A2(n2132), .ZN(n2063) );
  OR2_X2 U1676 ( .A1(n2131), .A2(n2132), .ZN(n2062) );
  OR2_X1 U1677 ( .A1(n2131), .A2(n2132), .ZN(n2070) );
  INV_X1 U1678 ( .A(n2218), .ZN(n2191) );
  XOR2_X1 U1679 ( .A(b[9]), .B(n1988), .Z(n1621) );
  INV_X2 U1680 ( .A(n2255), .ZN(n2253) );
  NAND3_X1 U1681 ( .A1(n2081), .A2(n2080), .A3(n2079), .ZN(n2064) );
  XOR2_X1 U1682 ( .A(n795), .B(n810), .Z(n2065) );
  XOR2_X1 U1683 ( .A(n808), .B(n2065), .Z(n791) );
  NAND2_X1 U1684 ( .A1(n808), .A2(n795), .ZN(n2066) );
  NAND2_X1 U1685 ( .A1(n808), .A2(n810), .ZN(n2067) );
  NAND2_X1 U1686 ( .A1(n795), .A2(n810), .ZN(n2068) );
  NAND3_X1 U1687 ( .A1(n2066), .A2(n2067), .A3(n2068), .ZN(n790) );
  INV_X1 U1688 ( .A(n2063), .ZN(n2130) );
  AND2_X2 U1689 ( .A1(n2105), .A2(n2032), .ZN(n2137) );
  INV_X1 U1690 ( .A(n1945), .ZN(n2243) );
  INV_X1 U1691 ( .A(n2237), .ZN(n2236) );
  XOR2_X1 U1692 ( .A(n887), .B(n904), .Z(n2072) );
  XOR2_X1 U1693 ( .A(n1969), .B(n2072), .Z(n881) );
  NAND2_X1 U1694 ( .A1(n902), .A2(n887), .ZN(n2073) );
  NAND2_X1 U1695 ( .A1(n902), .A2(n904), .ZN(n2074) );
  NAND2_X1 U1696 ( .A1(n887), .A2(n904), .ZN(n2075) );
  NAND3_X1 U1697 ( .A1(n2073), .A2(n2074), .A3(n2075), .ZN(n880) );
  INV_X1 U1698 ( .A(n2279), .ZN(n2076) );
  INV_X2 U1699 ( .A(n1936), .ZN(n2279) );
  CLKBUF_X1 U1700 ( .A(n489), .Z(n2156) );
  CLKBUF_X1 U1701 ( .A(n1982), .Z(n2077) );
  XNOR2_X1 U1702 ( .A(a[12]), .B(n2255), .ZN(n1811) );
  XOR2_X1 U1703 ( .A(n910), .B(n912), .Z(n2078) );
  XOR2_X1 U1704 ( .A(n2078), .B(n914), .Z(n887) );
  NAND2_X1 U1705 ( .A1(n910), .A2(n912), .ZN(n2079) );
  NAND2_X1 U1706 ( .A1(n910), .A2(n914), .ZN(n2080) );
  NAND2_X1 U1707 ( .A1(n912), .A2(n914), .ZN(n2081) );
  NAND3_X1 U1708 ( .A1(n2079), .A2(n2080), .A3(n2081), .ZN(n886) );
  XOR2_X1 U1709 ( .A(n888), .B(n873), .Z(n2082) );
  XOR2_X1 U1710 ( .A(n2082), .B(n886), .Z(n863) );
  NAND2_X1 U1711 ( .A1(n888), .A2(n873), .ZN(n2083) );
  NAND2_X1 U1712 ( .A1(n888), .A2(n2064), .ZN(n2084) );
  NAND2_X1 U1713 ( .A1(n873), .A2(n886), .ZN(n2085) );
  NAND3_X1 U1714 ( .A1(n2083), .A2(n2084), .A3(n2085), .ZN(n862) );
  INV_X1 U1715 ( .A(n2012), .ZN(n2086) );
  INV_X1 U1716 ( .A(n2086), .ZN(n2087) );
  INV_X1 U1717 ( .A(n2086), .ZN(n2088) );
  CLKBUF_X1 U1718 ( .A(n503), .Z(n2090) );
  XNOR2_X1 U1719 ( .A(a[11]), .B(a[12]), .ZN(n2091) );
  BUF_X1 U1720 ( .A(n2225), .Z(n2144) );
  NOR2_X1 U1721 ( .A1(n805), .A2(n820), .ZN(n2092) );
  NOR2_X1 U1722 ( .A1(n805), .A2(n820), .ZN(n495) );
  INV_X2 U1723 ( .A(n2186), .ZN(n2227) );
  CLKBUF_X1 U1724 ( .A(n512), .Z(n2094) );
  INV_X1 U1725 ( .A(n2248), .ZN(n2246) );
  CLKBUF_X3 U1726 ( .A(n295), .Z(n2187) );
  BUF_X2 U1727 ( .A(n277), .Z(n2195) );
  AND2_X2 U1728 ( .A1(n1810), .A2(n2000), .ZN(n2135) );
  INV_X1 U1729 ( .A(n2215), .ZN(n2096) );
  OAI21_X1 U1730 ( .B1(n535), .B2(n2071), .A(n2050), .ZN(n2097) );
  CLKBUF_X1 U1731 ( .A(n2187), .Z(n2098) );
  XOR2_X1 U1732 ( .A(n1296), .B(n1274), .Z(n2099) );
  XOR2_X1 U1733 ( .A(n818), .B(n2099), .Z(n797) );
  NAND2_X1 U1734 ( .A1(n818), .A2(n1296), .ZN(n2100) );
  NAND2_X1 U1735 ( .A1(n818), .A2(n1274), .ZN(n2101) );
  NAND2_X1 U1736 ( .A1(n1296), .A2(n1274), .ZN(n2102) );
  NAND3_X1 U1737 ( .A1(n2100), .A2(n2101), .A3(n2102), .ZN(n796) );
  INV_X1 U1738 ( .A(n2244), .ZN(n2242) );
  OAI21_X1 U1739 ( .B1(n538), .B2(n566), .A(n2051), .ZN(n537) );
  NOR2_X1 U1740 ( .A1(n695), .A2(n700), .ZN(n384) );
  NAND2_X1 U1741 ( .A1(n695), .A2(n700), .ZN(n387) );
  OR2_X1 U1742 ( .A1(n1143), .A2(n1150), .ZN(n2103) );
  XNOR2_X1 U1743 ( .A(n1933), .B(n2104), .ZN(n997) );
  XNOR2_X1 U1744 ( .A(n1372), .B(n1438), .ZN(n2104) );
  XOR2_X1 U1745 ( .A(a[4]), .B(a[5]), .Z(n2105) );
  INV_X1 U1746 ( .A(n537), .ZN(n536) );
  NOR2_X1 U1747 ( .A1(n2157), .A2(n467), .ZN(n465) );
  INV_X1 U1748 ( .A(n552), .ZN(n554) );
  NOR2_X1 U1749 ( .A1(n558), .A2(n563), .ZN(n552) );
  NAND2_X1 U1750 ( .A1(n662), .A2(n436), .ZN(n311) );
  OAI21_X1 U1751 ( .B1(n492), .B2(n467), .A(n468), .ZN(n466) );
  INV_X1 U1752 ( .A(n481), .ZN(n483) );
  INV_X1 U1753 ( .A(n521), .ZN(n519) );
  INV_X1 U1754 ( .A(n1980), .ZN(n565) );
  INV_X1 U1755 ( .A(n435), .ZN(n662) );
  NOR2_X1 U1756 ( .A1(n420), .A2(n402), .ZN(n400) );
  NAND2_X1 U1757 ( .A1(n666), .A2(n481), .ZN(n315) );
  NAND2_X1 U1758 ( .A1(n667), .A2(n496), .ZN(n316) );
  NAND2_X1 U1759 ( .A1(n669), .A2(n514), .ZN(n318) );
  NAND2_X1 U1760 ( .A1(n670), .A2(n521), .ZN(n319) );
  AOI21_X1 U1761 ( .B1(n565), .B2(n561), .A(n562), .ZN(n560) );
  AOI21_X1 U1762 ( .B1(n565), .B2(n545), .A(n546), .ZN(n544) );
  AOI21_X1 U1763 ( .B1(n662), .B2(n445), .A(n434), .ZN(n432) );
  INV_X1 U1764 ( .A(n436), .ZN(n434) );
  INV_X1 U1765 ( .A(n439), .ZN(n445) );
  INV_X1 U1766 ( .A(n520), .ZN(n670) );
  NOR2_X1 U1767 ( .A1(n402), .A2(n360), .ZN(n356) );
  INV_X1 U1768 ( .A(n563), .ZN(n561) );
  INV_X1 U1769 ( .A(n564), .ZN(n562) );
  INV_X1 U1770 ( .A(n438), .ZN(n663) );
  INV_X1 U1771 ( .A(n383), .ZN(n381) );
  NOR2_X1 U1772 ( .A1(n384), .A2(n364), .ZN(n362) );
  AOI21_X1 U1773 ( .B1(n426), .B2(n445), .A(n427), .ZN(n421) );
  NOR2_X1 U1774 ( .A1(n737), .A2(n748), .ZN(n435) );
  NOR2_X1 U1775 ( .A1(n983), .A2(n1002), .ZN(n563) );
  NAND2_X1 U1776 ( .A1(n657), .A2(n387), .ZN(n306) );
  NAND2_X1 U1777 ( .A1(n2115), .A2(n409), .ZN(n308) );
  NAND2_X1 U1778 ( .A1(n422), .A2(n2117), .ZN(n411) );
  INV_X1 U1779 ( .A(n382), .ZN(n380) );
  NAND2_X1 U1780 ( .A1(n2116), .A2(n396), .ZN(n307) );
  NAND2_X1 U1781 ( .A1(n2117), .A2(n418), .ZN(n309) );
  NAND2_X1 U1782 ( .A1(n661), .A2(n429), .ZN(n310) );
  INV_X1 U1783 ( .A(n428), .ZN(n661) );
  AOI21_X1 U1784 ( .B1(n401), .B2(n2116), .A(n394), .ZN(n390) );
  AND2_X1 U1785 ( .A1(n1021), .A2(n1038), .ZN(n2107) );
  NAND2_X1 U1786 ( .A1(n789), .A2(n804), .ZN(n481) );
  NAND2_X1 U1787 ( .A1(n857), .A2(n876), .ZN(n521) );
  NOR2_X1 U1788 ( .A1(n857), .A2(n876), .ZN(n520) );
  NOR2_X1 U1789 ( .A1(n435), .A2(n428), .ZN(n426) );
  NAND2_X1 U1790 ( .A1(n737), .A2(n748), .ZN(n436) );
  INV_X1 U1791 ( .A(n418), .ZN(n416) );
  AOI21_X1 U1792 ( .B1(n2115), .B2(n416), .A(n407), .ZN(n405) );
  INV_X1 U1793 ( .A(n409), .ZN(n407) );
  OR2_X1 U1794 ( .A1(n1021), .A2(n1038), .ZN(n2108) );
  OR2_X1 U1795 ( .A1(n761), .A2(n774), .ZN(n2109) );
  AOI21_X1 U1796 ( .B1(n423), .B2(n2117), .A(n416), .ZN(n412) );
  INV_X1 U1797 ( .A(n396), .ZN(n394) );
  XNOR2_X1 U1798 ( .A(n533), .B(n320), .ZN(product[26]) );
  NAND2_X1 U1799 ( .A1(n2117), .A2(n2115), .ZN(n402) );
  NAND2_X1 U1800 ( .A1(n362), .A2(n2116), .ZN(n360) );
  INV_X1 U1801 ( .A(n378), .ZN(n376) );
  OR2_X1 U1802 ( .A1(n1055), .A2(n1070), .ZN(n2110) );
  OR2_X1 U1803 ( .A1(n1039), .A2(n1054), .ZN(n2111) );
  AOI21_X1 U1804 ( .B1(n362), .B2(n394), .A(n363), .ZN(n361) );
  OAI21_X1 U1805 ( .B1(n364), .B2(n387), .A(n365), .ZN(n363) );
  AOI21_X1 U1806 ( .B1(n376), .B2(n2121), .A(n367), .ZN(n365) );
  NOR2_X1 U1807 ( .A1(n633), .A2(n631), .ZN(n629) );
  XNOR2_X1 U1808 ( .A(n921), .B(n2112), .ZN(n919) );
  XNOR2_X1 U1809 ( .A(n942), .B(n923), .ZN(n2112) );
  XNOR2_X1 U1810 ( .A(n899), .B(n2113), .ZN(n897) );
  XNOR2_X1 U1811 ( .A(n920), .B(n901), .ZN(n2113) );
  XNOR2_X1 U1812 ( .A(n2114), .B(n859), .ZN(n857) );
  XNOR2_X1 U1813 ( .A(n878), .B(n861), .ZN(n2114) );
  OR2_X2 U1814 ( .A1(n701), .A2(n708), .ZN(n2116) );
  OR2_X2 U1815 ( .A1(n717), .A2(n726), .ZN(n2117) );
  NAND2_X1 U1816 ( .A1(n2121), .A2(n369), .ZN(n304) );
  NAND2_X1 U1817 ( .A1(n2123), .A2(n341), .ZN(n302) );
  NAND2_X1 U1818 ( .A1(n2122), .A2(n352), .ZN(n303) );
  NOR2_X1 U1819 ( .A1(n1099), .A2(n1110), .ZN(n597) );
  AOI21_X1 U1820 ( .B1(n2119), .B2(n1950), .A(n1957), .ZN(n600) );
  OR2_X1 U1821 ( .A1(n1133), .A2(n1142), .ZN(n2118) );
  AOI21_X1 U1822 ( .B1(n2118), .B2(n1951), .A(n1958), .ZN(n611) );
  AOI21_X1 U1823 ( .B1(n359), .B2(n2122), .A(n350), .ZN(n348) );
  INV_X1 U1824 ( .A(n352), .ZN(n350) );
  AOI21_X1 U1825 ( .B1(n625), .B2(n1960), .A(n1952), .ZN(n620) );
  OAI21_X1 U1826 ( .B1(n628), .B2(n626), .A(n627), .ZN(n625) );
  OR2_X1 U1827 ( .A1(n1111), .A2(n1122), .ZN(n2119) );
  NAND2_X1 U1828 ( .A1(n701), .A2(n708), .ZN(n396) );
  NOR2_X1 U1829 ( .A1(n336), .A2(n334), .ZN(n332) );
  INV_X1 U1830 ( .A(n369), .ZN(n367) );
  NAND2_X1 U1831 ( .A1(n2103), .A2(n2118), .ZN(n610) );
  OR2_X1 U1832 ( .A1(n1123), .A2(n1132), .ZN(n2120) );
  NAND2_X1 U1833 ( .A1(n1099), .A2(n1110), .ZN(n598) );
  CLKBUF_X3 U1834 ( .A(a[21]), .Z(n2140) );
  AOI21_X1 U1835 ( .B1(n1948), .B2(n1947), .A(n1954), .ZN(n646) );
  NOR2_X1 U1836 ( .A1(n1165), .A2(n1170), .ZN(n631) );
  OR2_X2 U1837 ( .A1(n685), .A2(n688), .ZN(n2121) );
  OR2_X1 U1838 ( .A1(n681), .A2(n684), .ZN(n2122) );
  NAND2_X1 U1839 ( .A1(n678), .A2(n677), .ZN(n335) );
  INV_X1 U1840 ( .A(n341), .ZN(n339) );
  AOI21_X1 U1841 ( .B1(n643), .B2(n1949), .A(n1955), .ZN(n638) );
  OAI21_X1 U1842 ( .B1(n646), .B2(n644), .A(n645), .ZN(n643) );
  OR2_X1 U1843 ( .A1(n679), .A2(n680), .ZN(n2123) );
  NAND2_X1 U1844 ( .A1(n681), .A2(n684), .ZN(n352) );
  NAND2_X1 U1845 ( .A1(n679), .A2(n680), .ZN(n341) );
  NOR2_X1 U1846 ( .A1(n1175), .A2(n1178), .ZN(n636) );
  NAND2_X1 U1847 ( .A1(n1175), .A2(n1178), .ZN(n637) );
  INV_X1 U1848 ( .A(n676), .ZN(n677) );
  OR2_X1 U1849 ( .A1(n1194), .A2(n676), .ZN(n2124) );
  NOR2_X1 U1850 ( .A1(n678), .A2(n677), .ZN(n334) );
  AND2_X1 U1851 ( .A1(n1194), .A2(n676), .ZN(n2125) );
  OAI22_X1 U1852 ( .A1(n2220), .A2(n1779), .B1(n1778), .B2(n2005), .ZN(n1480)
         );
  INV_X1 U1853 ( .A(n2269), .ZN(n2267) );
  INV_X1 U1854 ( .A(n2259), .ZN(n2257) );
  INV_X1 U1855 ( .A(n2264), .ZN(n2262) );
  NAND2_X1 U1856 ( .A1(n2274), .A2(n1983), .ZN(n1756) );
  NOR2_X1 U1857 ( .A1(n2049), .A2(n1984), .ZN(n1457) );
  INV_X1 U1858 ( .A(n2129), .ZN(n2232) );
  INV_X1 U1859 ( .A(n2281), .ZN(n2278) );
  OAI21_X1 U1860 ( .B1(n2207), .B2(n2039), .A(n2293), .ZN(n1218) );
  INV_X1 U1861 ( .A(n1507), .ZN(n2293) );
  INV_X1 U1862 ( .A(n682), .ZN(n683) );
  NAND2_X1 U1863 ( .A1(n2270), .A2(n1983), .ZN(n1731) );
  NOR2_X1 U1864 ( .A1(n2141), .A2(n1984), .ZN(n1433) );
  NOR2_X1 U1865 ( .A1(n2002), .A2(n1984), .ZN(n1409) );
  INV_X1 U1866 ( .A(n692), .ZN(n693) );
  INV_X1 U1867 ( .A(n1632), .ZN(n2288) );
  OAI22_X1 U1868 ( .A1(n2220), .A2(n1777), .B1(n1776), .B2(n2235), .ZN(n1478)
         );
  NOR2_X1 U1869 ( .A1(n2037), .A2(n1983), .ZN(n1385) );
  INV_X1 U1870 ( .A(n1532), .ZN(n2292) );
  NAND2_X1 U1871 ( .A1(n2238), .A2(n1983), .ZN(n1531) );
  NAND2_X1 U1872 ( .A1(n2243), .A2(n1984), .ZN(n1556) );
  NAND2_X1 U1873 ( .A1(n2250), .A2(n2282), .ZN(n1606) );
  NAND2_X1 U1874 ( .A1(n1989), .A2(n1983), .ZN(n1656) );
  NAND2_X1 U1875 ( .A1(n2267), .A2(n1983), .ZN(n1706) );
  NAND2_X1 U1876 ( .A1(n1967), .A2(n1983), .ZN(n1681) );
  NAND2_X1 U1877 ( .A1(n2245), .A2(n1984), .ZN(n1581) );
  NOR2_X1 U1878 ( .A1(n1986), .A2(n1984), .ZN(n1217) );
  INV_X1 U1879 ( .A(n1682), .ZN(n2286) );
  NOR2_X1 U1880 ( .A1(n1974), .A2(n1984), .ZN(n1313) );
  OAI22_X1 U1881 ( .A1(n2220), .A2(n1769), .B1(n1768), .B2(n2006), .ZN(n1470)
         );
  OAI22_X1 U1882 ( .A1(n2219), .A2(n1770), .B1(n1769), .B2(n2006), .ZN(n1471)
         );
  OAI22_X1 U1883 ( .A1(n2220), .A2(n1772), .B1(n1771), .B2(n2006), .ZN(n1473)
         );
  OAI22_X1 U1884 ( .A1(n2220), .A2(n1775), .B1(n1774), .B2(n2005), .ZN(n1476)
         );
  NOR2_X1 U1885 ( .A1(n2088), .A2(n1983), .ZN(n1265) );
  NOR2_X1 U1886 ( .A1(n2226), .A2(n1984), .ZN(n1361) );
  OAI22_X1 U1887 ( .A1(n2220), .A2(n1771), .B1(n1770), .B2(n2006), .ZN(n1472)
         );
  OAI22_X1 U1888 ( .A1(n2220), .A2(n1774), .B1(n1773), .B2(n2005), .ZN(n1475)
         );
  NOR2_X1 U1889 ( .A1(n2038), .A2(n1984), .ZN(n1241) );
  INV_X1 U1890 ( .A(n1707), .ZN(n2285) );
  NOR2_X1 U1891 ( .A1(n1942), .A2(n1983), .ZN(n1337) );
  OAI22_X1 U1892 ( .A1(n2220), .A2(n1773), .B1(n1772), .B2(n2006), .ZN(n1474)
         );
  INV_X1 U1893 ( .A(n1557), .ZN(n2291) );
  INV_X1 U1894 ( .A(n1607), .ZN(n2289) );
  NOR2_X1 U1895 ( .A1(n2223), .A2(n1984), .ZN(n1289) );
  CLKBUF_X1 U1896 ( .A(n251), .Z(n2235) );
  OAI22_X1 U1897 ( .A1(n2220), .A2(n1780), .B1(n1779), .B2(n2235), .ZN(n1481)
         );
  NAND2_X1 U1898 ( .A1(n2280), .A2(n1983), .ZN(n1781) );
  INV_X1 U1899 ( .A(n802), .ZN(n803) );
  INV_X1 U1900 ( .A(n724), .ZN(n725) );
  INV_X1 U1901 ( .A(n874), .ZN(n875) );
  INV_X1 U1902 ( .A(n1732), .ZN(n2284) );
  INV_X1 U1903 ( .A(n1582), .ZN(n2290) );
  INV_X1 U1904 ( .A(n1657), .ZN(n2287) );
  INV_X1 U1905 ( .A(n1482), .ZN(n2294) );
  XNOR2_X1 U1906 ( .A(n2278), .B(b[6]), .ZN(n1774) );
  XNOR2_X1 U1907 ( .A(n2279), .B(b[2]), .ZN(n1778) );
  XNOR2_X1 U1908 ( .A(n2279), .B(b[4]), .ZN(n1776) );
  XNOR2_X1 U1909 ( .A(n2140), .B(b[0]), .ZN(n1530) );
  XNOR2_X1 U1910 ( .A(n2279), .B(b[10]), .ZN(n1770) );
  XNOR2_X1 U1911 ( .A(n2278), .B(b[8]), .ZN(n1772) );
  XNOR2_X1 U1912 ( .A(n2278), .B(b[12]), .ZN(n1768) );
  XNOR2_X1 U1913 ( .A(n2276), .B(b[22]), .ZN(n1733) );
  XNOR2_X1 U1914 ( .A(n2279), .B(b[16]), .ZN(n1764) );
  XNOR2_X1 U1915 ( .A(n2238), .B(b[16]), .ZN(n1514) );
  XNOR2_X1 U1916 ( .A(n2250), .B(b[12]), .ZN(n1593) );
  XNOR2_X1 U1917 ( .A(n2243), .B(b[16]), .ZN(n1539) );
  XNOR2_X1 U1918 ( .A(n2253), .B(b[16]), .ZN(n1614) );
  XNOR2_X1 U1919 ( .A(n1998), .B(b[12]), .ZN(n1568) );
  XNOR2_X1 U1920 ( .A(n2241), .B(b[12]), .ZN(n1543) );
  XNOR2_X1 U1921 ( .A(n2140), .B(b[6]), .ZN(n1524) );
  XNOR2_X1 U1922 ( .A(n2238), .B(b[12]), .ZN(n1518) );
  XNOR2_X1 U1923 ( .A(n2254), .B(b[12]), .ZN(n1618) );
  XNOR2_X1 U1924 ( .A(n2242), .B(b[6]), .ZN(n1549) );
  XNOR2_X1 U1925 ( .A(n2140), .B(b[4]), .ZN(n1526) );
  XNOR2_X1 U1926 ( .A(n2245), .B(b[16]), .ZN(n1564) );
  XNOR2_X1 U1927 ( .A(n2266), .B(b[16]), .ZN(n1689) );
  XNOR2_X1 U1928 ( .A(n2256), .B(b[16]), .ZN(n1639) );
  XNOR2_X1 U1929 ( .A(n2250), .B(b[16]), .ZN(n1589) );
  XNOR2_X1 U1930 ( .A(n2242), .B(b[4]), .ZN(n1551) );
  XNOR2_X1 U1931 ( .A(n1989), .B(b[12]), .ZN(n1643) );
  XNOR2_X1 U1932 ( .A(n2245), .B(b[4]), .ZN(n1576) );
  XNOR2_X1 U1933 ( .A(n2238), .B(b[2]), .ZN(n1528) );
  XNOR2_X1 U1934 ( .A(n1996), .B(b[6]), .ZN(n1574) );
  XNOR2_X1 U1935 ( .A(n2271), .B(b[16]), .ZN(n1714) );
  XNOR2_X1 U1936 ( .A(n2250), .B(b[6]), .ZN(n1599) );
  XNOR2_X1 U1937 ( .A(n2262), .B(b[12]), .ZN(n1668) );
  XNOR2_X1 U1938 ( .A(n2241), .B(b[2]), .ZN(n1553) );
  XNOR2_X1 U1939 ( .A(n1977), .B(b[4]), .ZN(n1601) );
  XNOR2_X1 U1940 ( .A(n2276), .B(b[16]), .ZN(n1739) );
  XNOR2_X1 U1941 ( .A(n1998), .B(b[2]), .ZN(n1578) );
  XNOR2_X1 U1942 ( .A(n2268), .B(b[12]), .ZN(n1693) );
  XNOR2_X1 U1943 ( .A(n2254), .B(b[6]), .ZN(n1624) );
  XNOR2_X1 U1944 ( .A(n2270), .B(b[12]), .ZN(n1718) );
  XNOR2_X1 U1945 ( .A(n2271), .B(b[6]), .ZN(n1724) );
  XNOR2_X1 U1946 ( .A(n1990), .B(b[4]), .ZN(n1651) );
  XNOR2_X1 U1947 ( .A(n2275), .B(b[12]), .ZN(n1743) );
  XNOR2_X1 U1948 ( .A(n1967), .B(b[2]), .ZN(n1678) );
  XNOR2_X1 U1949 ( .A(n2266), .B(b[2]), .ZN(n1703) );
  XNOR2_X1 U1950 ( .A(n2253), .B(b[2]), .ZN(n1628) );
  XNOR2_X1 U1951 ( .A(n2263), .B(b[16]), .ZN(n1664) );
  XNOR2_X1 U1952 ( .A(n2268), .B(b[4]), .ZN(n1701) );
  XNOR2_X1 U1953 ( .A(n2262), .B(b[6]), .ZN(n1674) );
  XNOR2_X1 U1954 ( .A(n1967), .B(b[4]), .ZN(n1676) );
  XNOR2_X1 U1955 ( .A(n2257), .B(b[6]), .ZN(n1649) );
  XNOR2_X1 U1956 ( .A(n2268), .B(b[6]), .ZN(n1699) );
  XNOR2_X1 U1957 ( .A(n2257), .B(b[2]), .ZN(n1653) );
  XNOR2_X1 U1958 ( .A(n2275), .B(b[4]), .ZN(n1751) );
  XNOR2_X1 U1959 ( .A(n2271), .B(b[4]), .ZN(n1726) );
  XNOR2_X1 U1960 ( .A(n2276), .B(b[6]), .ZN(n1749) );
  XNOR2_X1 U1961 ( .A(n2254), .B(b[4]), .ZN(n1626) );
  XNOR2_X1 U1962 ( .A(n2249), .B(b[2]), .ZN(n1603) );
  XNOR2_X1 U1963 ( .A(n2271), .B(b[2]), .ZN(n1728) );
  XNOR2_X1 U1964 ( .A(n2275), .B(b[2]), .ZN(n1753) );
  XNOR2_X1 U1965 ( .A(n2280), .B(b[20]), .ZN(n1760) );
  XNOR2_X1 U1966 ( .A(n2278), .B(b[22]), .ZN(n1758) );
  XNOR2_X1 U1967 ( .A(n2263), .B(b[22]), .ZN(n1658) );
  XNOR2_X1 U1968 ( .A(n2241), .B(b[20]), .ZN(n1535) );
  XNOR2_X1 U1969 ( .A(n2265), .B(b[22]), .ZN(n1683) );
  XNOR2_X1 U1970 ( .A(n2239), .B(b[20]), .ZN(n1510) );
  XNOR2_X1 U1971 ( .A(n2241), .B(b[22]), .ZN(n1533) );
  XNOR2_X1 U1972 ( .A(n2247), .B(b[20]), .ZN(n1560) );
  XNOR2_X1 U1973 ( .A(n2247), .B(b[22]), .ZN(n1558) );
  XNOR2_X1 U1974 ( .A(n2256), .B(b[20]), .ZN(n1635) );
  XNOR2_X1 U1975 ( .A(n2253), .B(b[22]), .ZN(n1608) );
  XNOR2_X1 U1976 ( .A(n2271), .B(b[20]), .ZN(n1710) );
  XNOR2_X1 U1977 ( .A(n2271), .B(b[22]), .ZN(n1708) );
  XNOR2_X1 U1978 ( .A(n2253), .B(b[20]), .ZN(n1610) );
  XNOR2_X1 U1979 ( .A(n2266), .B(b[20]), .ZN(n1685) );
  XNOR2_X1 U1980 ( .A(n2239), .B(b[22]), .ZN(n1508) );
  XNOR2_X1 U1981 ( .A(n1990), .B(b[22]), .ZN(n1633) );
  XNOR2_X1 U1982 ( .A(n2274), .B(b[20]), .ZN(n1735) );
  XNOR2_X1 U1983 ( .A(n2263), .B(b[20]), .ZN(n1660) );
  XNOR2_X1 U1984 ( .A(n2280), .B(b[18]), .ZN(n1762) );
  XNOR2_X1 U1985 ( .A(n2241), .B(b[18]), .ZN(n1537) );
  XNOR2_X1 U1986 ( .A(n2140), .B(b[18]), .ZN(n1512) );
  XNOR2_X1 U1987 ( .A(n2247), .B(b[18]), .ZN(n1562) );
  XNOR2_X1 U1988 ( .A(n2242), .B(b[10]), .ZN(n1545) );
  XNOR2_X1 U1989 ( .A(n2242), .B(b[8]), .ZN(n1547) );
  XNOR2_X1 U1990 ( .A(n1998), .B(b[10]), .ZN(n1570) );
  XNOR2_X1 U1991 ( .A(n2239), .B(b[10]), .ZN(n1520) );
  XNOR2_X1 U1992 ( .A(n2140), .B(b[8]), .ZN(n1522) );
  XNOR2_X1 U1993 ( .A(n1990), .B(b[18]), .ZN(n1637) );
  XNOR2_X1 U1994 ( .A(n1997), .B(b[8]), .ZN(n1572) );
  XNOR2_X1 U1995 ( .A(n2270), .B(b[18]), .ZN(n1712) );
  XNOR2_X1 U1996 ( .A(n2275), .B(b[18]), .ZN(n1737) );
  XNOR2_X1 U1997 ( .A(n2256), .B(b[10]), .ZN(n1645) );
  XNOR2_X1 U1998 ( .A(n1989), .B(b[8]), .ZN(n1647) );
  XNOR2_X1 U1999 ( .A(n1967), .B(b[10]), .ZN(n1670) );
  XNOR2_X1 U2000 ( .A(n2267), .B(b[10]), .ZN(n1695) );
  XNOR2_X1 U2001 ( .A(n2267), .B(b[8]), .ZN(n1697) );
  XNOR2_X1 U2002 ( .A(n2262), .B(b[18]), .ZN(n1662) );
  XNOR2_X1 U2003 ( .A(n2267), .B(b[18]), .ZN(n1687) );
  XNOR2_X1 U2004 ( .A(n1967), .B(b[8]), .ZN(n1672) );
  XNOR2_X1 U2005 ( .A(n2274), .B(b[10]), .ZN(n1745) );
  XNOR2_X1 U2006 ( .A(n2276), .B(b[8]), .ZN(n1747) );
  XNOR2_X1 U2007 ( .A(n2272), .B(b[8]), .ZN(n1722) );
  XNOR2_X1 U2008 ( .A(n2272), .B(b[10]), .ZN(n1720) );
  OAI22_X1 U2009 ( .A1(n2220), .A2(n1778), .B1(n1777), .B2(n2006), .ZN(n1479)
         );
  XNOR2_X1 U2010 ( .A(n2276), .B(b[0]), .ZN(n1755) );
  XNOR2_X1 U2011 ( .A(n2254), .B(b[0]), .ZN(n1630) );
  XNOR2_X1 U2012 ( .A(n2268), .B(b[0]), .ZN(n1705) );
  OAI22_X1 U2013 ( .A1(n2220), .A2(n1776), .B1(n1775), .B2(n2005), .ZN(n1477)
         );
  XNOR2_X1 U2014 ( .A(n2271), .B(b[0]), .ZN(n1730) );
  XNOR2_X1 U2015 ( .A(n2245), .B(b[0]), .ZN(n1580) );
  XNOR2_X1 U2016 ( .A(n1990), .B(b[0]), .ZN(n1655) );
  XNOR2_X1 U2017 ( .A(b[23]), .B(n2238), .ZN(n1507) );
  XNOR2_X1 U2018 ( .A(b[3]), .B(n2021), .ZN(n1502) );
  XNOR2_X1 U2019 ( .A(b[3]), .B(n2238), .ZN(n1527) );
  XNOR2_X1 U2020 ( .A(b[3]), .B(n2250), .ZN(n1602) );
  XNOR2_X1 U2021 ( .A(b[3]), .B(n2253), .ZN(n1627) );
  XNOR2_X1 U2022 ( .A(b[7]), .B(n2021), .ZN(n1498) );
  XNOR2_X1 U2023 ( .A(b[7]), .B(n2239), .ZN(n1523) );
  XNOR2_X1 U2024 ( .A(b[5]), .B(n2140), .ZN(n1525) );
  XNOR2_X1 U2025 ( .A(b[9]), .B(n2021), .ZN(n1496) );
  XNOR2_X1 U2026 ( .A(b[9]), .B(n2249), .ZN(n1596) );
  XNOR2_X1 U2027 ( .A(b[5]), .B(n2021), .ZN(n1500) );
  XNOR2_X1 U2028 ( .A(b[9]), .B(n2140), .ZN(n1521) );
  XNOR2_X1 U2029 ( .A(b[1]), .B(n2236), .ZN(n1504) );
  XNOR2_X1 U2030 ( .A(b[7]), .B(n1977), .ZN(n1598) );
  XNOR2_X1 U2031 ( .A(b[1]), .B(n2140), .ZN(n1529) );
  XNOR2_X1 U2032 ( .A(b[5]), .B(n1976), .ZN(n1600) );
  XNOR2_X1 U2033 ( .A(b[1]), .B(n2253), .ZN(n1629) );
  XNOR2_X1 U2034 ( .A(b[13]), .B(n2021), .ZN(n1492) );
  XNOR2_X1 U2035 ( .A(b[15]), .B(n2021), .ZN(n1490) );
  XNOR2_X1 U2036 ( .A(b[17]), .B(n2021), .ZN(n1488) );
  XNOR2_X1 U2037 ( .A(b[19]), .B(n2021), .ZN(n1486) );
  XNOR2_X1 U2038 ( .A(b[11]), .B(n2021), .ZN(n1494) );
  XNOR2_X1 U2039 ( .A(b[21]), .B(n2021), .ZN(n1484) );
  INV_X1 U2040 ( .A(n2093), .ZN(n2132) );
  XNOR2_X1 U2041 ( .A(n2278), .B(b[0]), .ZN(n1780) );
  INV_X1 U2042 ( .A(a[11]), .ZN(n2259) );
  OAI21_X1 U2043 ( .B1(a[0]), .B2(n2138), .A(n2283), .ZN(n1458) );
  INV_X1 U2044 ( .A(n1757), .ZN(n2283) );
  OR2_X1 U2045 ( .A1(n2139), .A2(n2129), .ZN(n277) );
  XNOR2_X1 U2046 ( .A(a[2]), .B(a[3]), .ZN(n2139) );
  XNOR2_X1 U2047 ( .A(n2241), .B(b[0]), .ZN(n1555) );
  XNOR2_X1 U2048 ( .A(n2263), .B(b[0]), .ZN(n1680) );
  INV_X1 U2049 ( .A(a[0]), .ZN(n251) );
  XNOR2_X1 U2050 ( .A(b[23]), .B(n2021), .ZN(n1482) );
  XNOR2_X1 U2051 ( .A(n1998), .B(b[14]), .ZN(n1566) );
  XNOR2_X1 U2052 ( .A(n2243), .B(b[14]), .ZN(n1541) );
  XNOR2_X1 U2053 ( .A(n2262), .B(b[14]), .ZN(n1666) );
  XNOR2_X1 U2054 ( .A(n2275), .B(b[14]), .ZN(n1741) );
  XNOR2_X1 U2055 ( .A(n2272), .B(b[14]), .ZN(n1716) );
  XNOR2_X1 U2056 ( .A(n1977), .B(b[14]), .ZN(n1591) );
  XNOR2_X1 U2057 ( .A(n2238), .B(b[14]), .ZN(n1516) );
  XNOR2_X1 U2058 ( .A(n2278), .B(b[14]), .ZN(n1766) );
  XNOR2_X1 U2059 ( .A(n2253), .B(b[14]), .ZN(n1616) );
  XNOR2_X1 U2060 ( .A(n2257), .B(b[14]), .ZN(n1641) );
  XNOR2_X1 U2061 ( .A(n2268), .B(b[14]), .ZN(n1691) );
  INV_X1 U2062 ( .A(a[7]), .ZN(n2269) );
  INV_X1 U2063 ( .A(a[15]), .ZN(n2251) );
  NAND2_X1 U2064 ( .A1(n839), .A2(n856), .ZN(n514) );
  INV_X1 U2065 ( .A(a[19]), .ZN(n2244) );
  INV_X1 U2066 ( .A(n505), .ZN(n507) );
  OAI21_X1 U2067 ( .B1(n2212), .B2(n2175), .A(n2289), .ZN(n1314) );
  INV_X1 U2068 ( .A(n2092), .ZN(n667) );
  NAND2_X1 U2069 ( .A1(n1159), .A2(n1161), .ZN(n627) );
  NOR2_X1 U2070 ( .A1(n1159), .A2(n1161), .ZN(n626) );
  XNOR2_X1 U2071 ( .A(b[9]), .B(n2276), .ZN(n1746) );
  XNOR2_X1 U2072 ( .A(b[7]), .B(n2274), .ZN(n1748) );
  XNOR2_X1 U2073 ( .A(b[1]), .B(n2274), .ZN(n1754) );
  XNOR2_X1 U2074 ( .A(b[3]), .B(n2275), .ZN(n1752) );
  XNOR2_X1 U2075 ( .A(b[5]), .B(n2275), .ZN(n1750) );
  XNOR2_X1 U2076 ( .A(b[23]), .B(n2275), .ZN(n1732) );
  NOR2_X1 U2077 ( .A1(n856), .A2(n839), .ZN(n2147) );
  NOR2_X1 U2078 ( .A1(n839), .A2(n856), .ZN(n513) );
  NAND2_X1 U2079 ( .A1(n668), .A2(n2090), .ZN(n317) );
  INV_X1 U2080 ( .A(n503), .ZN(n501) );
  NAND2_X1 U2081 ( .A1(n821), .A2(n838), .ZN(n503) );
  INV_X1 U2082 ( .A(a[9]), .ZN(n2264) );
  INV_X1 U2083 ( .A(a[13]), .ZN(n2255) );
  XNOR2_X1 U2084 ( .A(n2021), .B(b[22]), .ZN(n1483) );
  XNOR2_X1 U2085 ( .A(n2021), .B(b[18]), .ZN(n1487) );
  XNOR2_X1 U2086 ( .A(n2021), .B(b[20]), .ZN(n1485) );
  XNOR2_X1 U2087 ( .A(n2021), .B(b[10]), .ZN(n1495) );
  NAND2_X1 U2088 ( .A1(n2021), .A2(n2282), .ZN(n1506) );
  XNOR2_X1 U2089 ( .A(n2021), .B(b[16]), .ZN(n1489) );
  XNOR2_X1 U2090 ( .A(n2021), .B(b[14]), .ZN(n1491) );
  XNOR2_X1 U2091 ( .A(n2021), .B(b[12]), .ZN(n1493) );
  XNOR2_X1 U2092 ( .A(n2021), .B(b[4]), .ZN(n1501) );
  XNOR2_X1 U2093 ( .A(n2021), .B(b[8]), .ZN(n1497) );
  XNOR2_X1 U2094 ( .A(n2021), .B(b[0]), .ZN(n1505) );
  XNOR2_X1 U2095 ( .A(n2021), .B(b[6]), .ZN(n1499) );
  XNOR2_X1 U2096 ( .A(n2021), .B(b[2]), .ZN(n1503) );
  INV_X1 U2097 ( .A(a[23]), .ZN(n2237) );
  OAI21_X1 U2098 ( .B1(n503), .B2(n2092), .A(n496), .ZN(n2148) );
  XNOR2_X1 U2099 ( .A(n515), .B(n318), .ZN(product[28]) );
  NOR2_X1 U2100 ( .A1(n597), .A2(n599), .ZN(n595) );
  XNOR2_X1 U2101 ( .A(b[1]), .B(n2267), .ZN(n1704) );
  XNOR2_X1 U2102 ( .A(b[5]), .B(n2267), .ZN(n1700) );
  XNOR2_X1 U2103 ( .A(b[3]), .B(n2266), .ZN(n1702) );
  XNOR2_X1 U2104 ( .A(b[7]), .B(n2266), .ZN(n1698) );
  XNOR2_X1 U2105 ( .A(b[9]), .B(n2266), .ZN(n1696) );
  XNOR2_X1 U2106 ( .A(b[23]), .B(n2265), .ZN(n1682) );
  NAND2_X1 U2107 ( .A1(n921), .A2(n942), .ZN(n2149) );
  NAND2_X1 U2108 ( .A1(n921), .A2(n923), .ZN(n2150) );
  NAND2_X1 U2109 ( .A1(n942), .A2(n923), .ZN(n2151) );
  NAND3_X1 U2110 ( .A1(n2149), .A2(n2150), .A3(n2151), .ZN(n918) );
  NAND2_X1 U2111 ( .A1(n2252), .A2(n1984), .ZN(n1631) );
  XNOR2_X1 U2112 ( .A(n2252), .B(b[18]), .ZN(n1612) );
  XNOR2_X1 U2113 ( .A(b[5]), .B(n2252), .ZN(n1625) );
  XNOR2_X1 U2114 ( .A(n2252), .B(b[10]), .ZN(n1620) );
  XNOR2_X1 U2115 ( .A(b[7]), .B(n2252), .ZN(n1623) );
  XNOR2_X1 U2116 ( .A(b[23]), .B(n2252), .ZN(n1607) );
  XNOR2_X1 U2117 ( .A(n522), .B(n319), .ZN(product[27]) );
  XNOR2_X1 U2118 ( .A(n497), .B(n316), .ZN(product[30]) );
  XNOR2_X1 U2119 ( .A(n486), .B(n315), .ZN(product[31]) );
  XNOR2_X1 U2120 ( .A(n475), .B(n314), .ZN(product[32]) );
  NAND2_X1 U2121 ( .A1(n899), .A2(n920), .ZN(n2152) );
  NAND2_X1 U2122 ( .A1(n899), .A2(n901), .ZN(n2153) );
  NAND2_X1 U2123 ( .A1(n920), .A2(n901), .ZN(n2154) );
  NAND3_X1 U2124 ( .A1(n2152), .A2(n2153), .A3(n2154), .ZN(n896) );
  OAI21_X1 U2125 ( .B1(n2130), .B2(n2186), .A(n2287), .ZN(n1362) );
  NOR2_X1 U2126 ( .A1(n877), .A2(n896), .ZN(n2155) );
  XNOR2_X1 U2127 ( .A(n1976), .B(b[18]), .ZN(n1587) );
  XNOR2_X1 U2128 ( .A(n2249), .B(b[22]), .ZN(n1583) );
  XNOR2_X1 U2129 ( .A(n2249), .B(b[20]), .ZN(n1585) );
  XNOR2_X1 U2130 ( .A(b[23]), .B(n2250), .ZN(n1582) );
  XNOR2_X1 U2131 ( .A(n1977), .B(b[0]), .ZN(n1605) );
  XNOR2_X1 U2132 ( .A(n1977), .B(b[8]), .ZN(n1597) );
  XNOR2_X1 U2133 ( .A(n2249), .B(b[10]), .ZN(n1595) );
  XNOR2_X1 U2134 ( .A(b[1]), .B(n2250), .ZN(n1604) );
  INV_X1 U2135 ( .A(a[3]), .ZN(n2277) );
  OR2_X1 U2136 ( .A1(n2092), .A2(n502), .ZN(n2157) );
  INV_X1 U2137 ( .A(a[5]), .ZN(n2273) );
  XNOR2_X1 U2138 ( .A(b[3]), .B(n2261), .ZN(n1677) );
  XNOR2_X1 U2139 ( .A(b[9]), .B(n2261), .ZN(n1671) );
  XNOR2_X1 U2140 ( .A(b[1]), .B(n2261), .ZN(n1679) );
  XNOR2_X1 U2141 ( .A(b[5]), .B(n2261), .ZN(n1675) );
  XNOR2_X1 U2142 ( .A(b[7]), .B(n2261), .ZN(n1673) );
  XNOR2_X1 U2143 ( .A(b[23]), .B(n2261), .ZN(n1657) );
  INV_X1 U2144 ( .A(n672), .ZN(n2159) );
  INV_X1 U2145 ( .A(n492), .ZN(n2160) );
  OAI21_X1 U2146 ( .B1(n2137), .B2(n2192), .A(n2285), .ZN(n1410) );
  XNOR2_X1 U2147 ( .A(b[1]), .B(n2245), .ZN(n1579) );
  XNOR2_X1 U2148 ( .A(b[5]), .B(n1997), .ZN(n1575) );
  XNOR2_X1 U2149 ( .A(b[3]), .B(n1997), .ZN(n1577) );
  XNOR2_X1 U2150 ( .A(b[23]), .B(n2247), .ZN(n1557) );
  XNOR2_X1 U2151 ( .A(b[7]), .B(n2245), .ZN(n1573) );
  XNOR2_X1 U2152 ( .A(b[9]), .B(n1996), .ZN(n1571) );
  INV_X2 U2153 ( .A(n2269), .ZN(n2266) );
  XNOR2_X1 U2154 ( .A(b[23]), .B(n2243), .ZN(n1532) );
  XNOR2_X1 U2155 ( .A(b[1]), .B(n2243), .ZN(n1554) );
  XNOR2_X1 U2156 ( .A(b[5]), .B(n2243), .ZN(n1550) );
  XNOR2_X1 U2157 ( .A(b[7]), .B(n2242), .ZN(n1548) );
  XNOR2_X1 U2158 ( .A(b[9]), .B(n2242), .ZN(n1546) );
  XNOR2_X1 U2159 ( .A(b[3]), .B(n2243), .ZN(n1552) );
  XOR2_X1 U2160 ( .A(n863), .B(n882), .Z(n2161) );
  XOR2_X1 U2161 ( .A(n2161), .B(n880), .Z(n859) );
  NAND2_X1 U2162 ( .A1(n863), .A2(n882), .ZN(n2162) );
  NAND2_X1 U2163 ( .A1(n863), .A2(n2031), .ZN(n2163) );
  NAND2_X1 U2164 ( .A1(n882), .A2(n880), .ZN(n2164) );
  NAND3_X1 U2165 ( .A1(n2162), .A2(n2163), .A3(n2164), .ZN(n858) );
  NAND2_X1 U2166 ( .A1(n878), .A2(n861), .ZN(n2165) );
  NAND2_X1 U2167 ( .A1(n878), .A2(n859), .ZN(n2166) );
  NAND2_X1 U2168 ( .A1(n861), .A2(n859), .ZN(n2167) );
  NAND3_X1 U2169 ( .A1(n2165), .A2(n2166), .A3(n2167), .ZN(n856) );
  XNOR2_X1 U2170 ( .A(b[3]), .B(n2256), .ZN(n1652) );
  XNOR2_X1 U2171 ( .A(b[7]), .B(n2258), .ZN(n1648) );
  XNOR2_X1 U2172 ( .A(b[23]), .B(n2258), .ZN(n1632) );
  XNOR2_X1 U2173 ( .A(b[9]), .B(n2257), .ZN(n1646) );
  XNOR2_X1 U2174 ( .A(b[1]), .B(n2258), .ZN(n1654) );
  XNOR2_X1 U2175 ( .A(b[5]), .B(n2258), .ZN(n1650) );
  INV_X1 U2176 ( .A(n2126), .ZN(n2168) );
  XNOR2_X1 U2177 ( .A(b[3]), .B(n2271), .ZN(n1727) );
  XNOR2_X1 U2178 ( .A(b[9]), .B(n2272), .ZN(n1721) );
  XNOR2_X1 U2179 ( .A(b[5]), .B(n2270), .ZN(n1725) );
  XNOR2_X1 U2180 ( .A(b[1]), .B(n2270), .ZN(n1729) );
  XNOR2_X1 U2181 ( .A(b[7]), .B(n2271), .ZN(n1723) );
  XNOR2_X1 U2182 ( .A(b[23]), .B(n2272), .ZN(n1707) );
  INV_X1 U2183 ( .A(a[17]), .ZN(n2248) );
  NOR2_X1 U2184 ( .A1(n896), .A2(n2008), .ZN(n531) );
  NAND2_X1 U2185 ( .A1(n2176), .A2(n2050), .ZN(n320) );
  OR2_X1 U2186 ( .A1(n420), .A2(n347), .ZN(n2170) );
  NAND2_X1 U2187 ( .A1(n426), .A2(n663), .ZN(n420) );
  NAND2_X1 U2188 ( .A1(n356), .A2(n2122), .ZN(n347) );
  XNOR2_X1 U2189 ( .A(n1023), .B(n2171), .ZN(n1021) );
  XNOR2_X1 U2190 ( .A(n1040), .B(n1025), .ZN(n2171) );
  INV_X1 U2191 ( .A(a[21]), .ZN(n2240) );
  INV_X1 U2192 ( .A(n2205), .ZN(n2172) );
  NOR2_X1 U2193 ( .A1(n502), .A2(n495), .ZN(n489) );
  OAI21_X1 U2194 ( .B1(n2218), .B2(n1994), .A(n2284), .ZN(n1434) );
  CLKBUF_X1 U2195 ( .A(n535), .Z(n2174) );
  OAI21_X1 U2196 ( .B1(n2055), .B2(n2230), .A(n2286), .ZN(n1386) );
  NAND2_X1 U2197 ( .A1(n941), .A2(n962), .ZN(n550) );
  NAND2_X1 U2198 ( .A1(n919), .A2(n940), .ZN(n543) );
  INV_X1 U2199 ( .A(n297), .ZN(n2205) );
  OR2_X1 U2200 ( .A1(n2020), .A2(n896), .ZN(n2176) );
  XNOR2_X1 U2201 ( .A(b[13]), .B(n2272), .ZN(n1717) );
  INV_X1 U2202 ( .A(n257), .ZN(n2230) );
  INV_X1 U2203 ( .A(n2264), .ZN(n2260) );
  INV_X1 U2204 ( .A(n2207), .ZN(n2179) );
  OAI22_X1 U2205 ( .A1(n2220), .A2(n1767), .B1(n1766), .B2(n2005), .ZN(n1468)
         );
  OAI22_X1 U2206 ( .A1(n2220), .A2(n1768), .B1(n1767), .B2(n2235), .ZN(n1469)
         );
  OAI22_X1 U2207 ( .A1(n2220), .A2(n1764), .B1(n1763), .B2(n2005), .ZN(n1465)
         );
  OAI22_X1 U2208 ( .A1(n2220), .A2(n1765), .B1(n1764), .B2(n2006), .ZN(n1466)
         );
  OAI22_X1 U2209 ( .A1(n2220), .A2(n1759), .B1(n1758), .B2(n2005), .ZN(n1460)
         );
  OAI22_X1 U2210 ( .A1(n2219), .A2(n1760), .B1(n1759), .B2(n2235), .ZN(n1461)
         );
  OAI22_X1 U2211 ( .A1(n2219), .A2(n1763), .B1(n1762), .B2(n2005), .ZN(n1464)
         );
  OAI22_X1 U2212 ( .A1(n2219), .A2(n1761), .B1(n1760), .B2(n2005), .ZN(n1462)
         );
  OAI22_X1 U2213 ( .A1(n2219), .A2(n1758), .B1(n1757), .B2(n2006), .ZN(n1459)
         );
  XNOR2_X1 U2214 ( .A(b[1]), .B(n2280), .ZN(n1779) );
  OAI22_X1 U2215 ( .A1(n2219), .A2(n1766), .B1(n1765), .B2(n2006), .ZN(n1467)
         );
  OAI22_X1 U2216 ( .A1(n2219), .A2(n1762), .B1(n1761), .B2(n2005), .ZN(n1463)
         );
  XNOR2_X1 U2217 ( .A(b[3]), .B(n2279), .ZN(n1777) );
  XNOR2_X1 U2218 ( .A(b[5]), .B(n2279), .ZN(n1775) );
  XNOR2_X1 U2219 ( .A(b[9]), .B(n2279), .ZN(n1771) );
  XNOR2_X1 U2220 ( .A(b[7]), .B(n2279), .ZN(n1773) );
  XNOR2_X1 U2221 ( .A(b[23]), .B(n2279), .ZN(n1757) );
  OR2_X1 U2222 ( .A1(n2180), .A2(n1622), .ZN(n2181) );
  OR2_X1 U2223 ( .A1(n1621), .A2(n2142), .ZN(n2182) );
  NAND2_X1 U2224 ( .A1(n2181), .A2(n2182), .ZN(n1328) );
  XNOR2_X1 U2225 ( .A(n2254), .B(b[8]), .ZN(n1622) );
  NAND2_X1 U2226 ( .A1(n1023), .A2(n1040), .ZN(n2183) );
  NAND2_X1 U2227 ( .A1(n1023), .A2(n1025), .ZN(n2184) );
  NAND2_X1 U2228 ( .A1(n1040), .A2(n1025), .ZN(n2185) );
  NAND3_X1 U2229 ( .A1(n2183), .A2(n2184), .A3(n2185), .ZN(n1020) );
  NOR2_X1 U2230 ( .A1(n1003), .A2(n1020), .ZN(n569) );
  OAI21_X1 U2231 ( .B1(n2135), .B2(n2158), .A(n2290), .ZN(n1290) );
  INV_X1 U2232 ( .A(n2205), .ZN(n2204) );
  OAI21_X1 U2233 ( .B1(n2136), .B2(n2178), .A(n2288), .ZN(n1338) );
  INV_X1 U2234 ( .A(n295), .ZN(n2207) );
  OAI21_X1 U2235 ( .B1(n2205), .B2(n2127), .A(n2294), .ZN(n1194) );
  OAI22_X1 U2236 ( .A1(n2098), .A2(n1513), .B1(n2038), .B2(n1512), .ZN(n1223)
         );
  OAI22_X1 U2237 ( .A1(n2187), .A2(n1511), .B1(n2038), .B2(n1510), .ZN(n1221)
         );
  OAI22_X1 U2238 ( .A1(n2187), .A2(n1515), .B1(n2038), .B2(n1514), .ZN(n1225)
         );
  OAI22_X1 U2239 ( .A1(n2187), .A2(n1509), .B1(n2038), .B2(n1508), .ZN(n1219)
         );
  OAI22_X1 U2240 ( .A1(n2187), .A2(n1517), .B1(n2038), .B2(n1516), .ZN(n1227)
         );
  OAI21_X1 U2241 ( .B1(n590), .B2(n593), .A(n591), .ZN(n589) );
  NOR2_X1 U2242 ( .A1(n1071), .A2(n1084), .ZN(n590) );
  INV_X1 U2243 ( .A(n2277), .ZN(n2274) );
  INV_X1 U2244 ( .A(n281), .ZN(n2215) );
  OAI21_X1 U2245 ( .B1(n2133), .B2(n2009), .A(n2291), .ZN(n1266) );
  OAI22_X1 U2246 ( .A1(n2014), .A2(n1634), .B1(n2146), .B2(n1633), .ZN(n1339)
         );
  OAI22_X1 U2247 ( .A1(n2015), .A2(n1636), .B1(n2226), .B2(n1635), .ZN(n1341)
         );
  OAI22_X1 U2248 ( .A1(n2213), .A2(n1640), .B1(n2226), .B2(n1639), .ZN(n1345)
         );
  OAI22_X1 U2249 ( .A1(n2015), .A2(n1638), .B1(n2226), .B2(n1637), .ZN(n1343)
         );
  INV_X1 U2250 ( .A(n2207), .ZN(n2206) );
  NOR2_X1 U2251 ( .A1(n919), .A2(n940), .ZN(n2194) );
  NOR2_X1 U2252 ( .A1(n919), .A2(n940), .ZN(n542) );
  OAI21_X1 U2253 ( .B1(n405), .B2(n360), .A(n361), .ZN(n359) );
  XNOR2_X1 U2254 ( .A(b[19]), .B(n1990), .ZN(n1636) );
  XNOR2_X1 U2255 ( .A(b[21]), .B(n1989), .ZN(n1634) );
  INV_X1 U2256 ( .A(n384), .ZN(n657) );
  NOR2_X1 U2257 ( .A1(n389), .A2(n384), .ZN(n382) );
  OAI21_X1 U2258 ( .B1(n390), .B2(n384), .A(n387), .ZN(n383) );
  OAI22_X1 U2259 ( .A1(n2209), .A2(n1536), .B1(n2089), .B2(n1535), .ZN(n1245)
         );
  OAI22_X1 U2260 ( .A1(n2208), .A2(n1534), .B1(n2089), .B2(n1533), .ZN(n1243)
         );
  OAI22_X1 U2261 ( .A1(n2169), .A2(n1542), .B1(n2088), .B2(n1541), .ZN(n1251)
         );
  OAI22_X1 U2262 ( .A1(n2208), .A2(n1540), .B1(n2089), .B2(n1539), .ZN(n1249)
         );
  OAI22_X1 U2263 ( .A1(n2208), .A2(n1538), .B1(n2088), .B2(n1537), .ZN(n1247)
         );
  INV_X1 U2264 ( .A(n2215), .ZN(n2214) );
  NAND2_X1 U2265 ( .A1(n2109), .A2(n461), .ZN(n313) );
  INV_X1 U2266 ( .A(n461), .ZN(n459) );
  AOI21_X1 U2267 ( .B1(n629), .B2(n635), .A(n630), .ZN(n628) );
  OAI21_X1 U2268 ( .B1(n638), .B2(n636), .A(n637), .ZN(n635) );
  OAI21_X1 U2269 ( .B1(n620), .B2(n610), .A(n611), .ZN(n609) );
  NAND2_X1 U2270 ( .A1(n2034), .A2(n2109), .ZN(n456) );
  INV_X1 U2271 ( .A(n400), .ZN(n398) );
  NAND2_X1 U2272 ( .A1(n400), .A2(n2116), .ZN(n389) );
  NOR2_X1 U2273 ( .A1(n590), .A2(n592), .ZN(n588) );
  AOI21_X1 U2274 ( .B1(n565), .B2(n1932), .A(n2053), .ZN(n551) );
  INV_X1 U2275 ( .A(n558), .ZN(n675) );
  INV_X1 U2276 ( .A(n553), .ZN(n555) );
  OAI21_X1 U2277 ( .B1(n558), .B2(n564), .A(n559), .ZN(n553) );
  INV_X1 U2278 ( .A(n542), .ZN(n673) );
  OAI21_X1 U2279 ( .B1(n2126), .B2(n2086), .A(n2292), .ZN(n1242) );
  INV_X1 U2280 ( .A(n277), .ZN(n2218) );
  NAND2_X1 U2281 ( .A1(n1085), .A2(n1098), .ZN(n593) );
  NOR2_X1 U2282 ( .A1(n1085), .A2(n1098), .ZN(n592) );
  OAI21_X1 U2283 ( .B1(n600), .B2(n597), .A(n598), .ZN(n596) );
  INV_X1 U2284 ( .A(n401), .ZN(n399) );
  INV_X1 U2285 ( .A(n421), .ZN(n423) );
  NAND2_X1 U2286 ( .A1(n2008), .A2(n896), .ZN(n532) );
  NAND2_X1 U2287 ( .A1(n1806), .A2(n2030), .ZN(n297) );
  NOR2_X1 U2288 ( .A1(n571), .A2(n569), .ZN(n567) );
  NAND2_X1 U2289 ( .A1(n1003), .A2(n1020), .ZN(n570) );
  INV_X1 U2290 ( .A(n2148), .ZN(n492) );
  NAND2_X1 U2291 ( .A1(n685), .A2(n688), .ZN(n369) );
  NOR2_X1 U2292 ( .A1(n1181), .A2(n1192), .ZN(n644) );
  NAND2_X1 U2293 ( .A1(n1181), .A2(n1192), .ZN(n645) );
  AOI21_X1 U2294 ( .B1(n2097), .B2(n2077), .A(n2094), .ZN(n2196) );
  NAND2_X1 U2295 ( .A1(n983), .A2(n1002), .ZN(n564) );
  INV_X1 U2296 ( .A(n2019), .ZN(n674) );
  NOR2_X1 U2297 ( .A1(n554), .A2(n2019), .ZN(n545) );
  OAI21_X1 U2298 ( .B1(n555), .B2(n2019), .A(n1930), .ZN(n546) );
  NAND2_X1 U2299 ( .A1(n2119), .A2(n2120), .ZN(n599) );
  NAND2_X1 U2300 ( .A1(n963), .A2(n982), .ZN(n559) );
  XNOR2_X1 U2301 ( .A(b[21]), .B(n2243), .ZN(n1534) );
  XNOR2_X1 U2302 ( .A(b[19]), .B(n2241), .ZN(n1536) );
  XNOR2_X1 U2303 ( .A(b[13]), .B(n2241), .ZN(n1542) );
  XNOR2_X1 U2304 ( .A(b[11]), .B(n2242), .ZN(n1544) );
  XNOR2_X1 U2305 ( .A(b[17]), .B(n2241), .ZN(n1538) );
  XNOR2_X1 U2306 ( .A(b[15]), .B(n2241), .ZN(n1540) );
  INV_X1 U2307 ( .A(n420), .ZN(n422) );
  NOR2_X1 U2308 ( .A1(n420), .A2(n347), .ZN(n345) );
  NAND2_X1 U2309 ( .A1(n727), .A2(n736), .ZN(n429) );
  NOR2_X2 U2310 ( .A1(n727), .A2(n736), .ZN(n428) );
  OAI22_X1 U2311 ( .A1(n2210), .A2(n1593), .B1(n1592), .B2(n1965), .ZN(n1300)
         );
  OAI22_X1 U2312 ( .A1(n2210), .A2(n1590), .B1(n1965), .B2(n1589), .ZN(n1297)
         );
  OAI22_X1 U2313 ( .A1(n2004), .A2(n1589), .B1(n1588), .B2(n1965), .ZN(n1296)
         );
  OAI22_X1 U2314 ( .A1(n2003), .A2(n1584), .B1(n2000), .B2(n1583), .ZN(n1291)
         );
  OAI22_X1 U2315 ( .A1(n2003), .A2(n1583), .B1(n1582), .B2(n1974), .ZN(n724)
         );
  OAI22_X1 U2316 ( .A1(n2003), .A2(n1592), .B1(n1964), .B2(n1591), .ZN(n1299)
         );
  OAI22_X1 U2317 ( .A1(n2004), .A2(n1585), .B1(n1584), .B2(n1974), .ZN(n1292)
         );
  OAI22_X1 U2318 ( .A1(n2004), .A2(n1588), .B1(n1965), .B2(n1587), .ZN(n1295)
         );
  OAI22_X1 U2319 ( .A1(n2004), .A2(n1591), .B1(n1590), .B2(n1965), .ZN(n1298)
         );
  OAI22_X1 U2320 ( .A1(n1606), .A2(n1964), .B1(n2211), .B2(n1995), .ZN(n1186)
         );
  OAI22_X1 U2321 ( .A1(n2003), .A2(n1587), .B1(n1586), .B2(n1965), .ZN(n1294)
         );
  OAI22_X1 U2322 ( .A1(n2210), .A2(n1586), .B1(n1965), .B2(n1585), .ZN(n1293)
         );
  AOI21_X1 U2323 ( .B1(n2109), .B2(n2036), .A(n459), .ZN(n457) );
  INV_X1 U2324 ( .A(n508), .ZN(n2197) );
  AOI21_X1 U2325 ( .B1(n511), .B2(n526), .A(n512), .ZN(n506) );
  NAND2_X1 U2326 ( .A1(n761), .A2(n774), .ZN(n461) );
  AOI21_X1 U2327 ( .B1(n2108), .B2(n1956), .A(n2107), .ZN(n572) );
  NAND2_X1 U2328 ( .A1(n2108), .A2(n2111), .ZN(n571) );
  NAND2_X1 U2329 ( .A1(n588), .A2(n2110), .ZN(n582) );
  AOI21_X1 U2330 ( .B1(n589), .B2(n2110), .A(n1959), .ZN(n583) );
  NAND2_X1 U2331 ( .A1(n672), .A2(n2174), .ZN(n321) );
  OAI21_X1 U2332 ( .B1(n2155), .B2(n535), .A(n532), .ZN(n526) );
  NOR2_X1 U2333 ( .A1(n2157), .A2(n480), .ZN(n478) );
  OAI21_X1 U2334 ( .B1(n492), .B2(n480), .A(n481), .ZN(n479) );
  INV_X1 U2335 ( .A(n480), .ZN(n666) );
  NOR2_X1 U2336 ( .A1(n480), .A2(n456), .ZN(n454) );
  NOR2_X2 U2337 ( .A1(n789), .A2(n804), .ZN(n480) );
  NAND2_X1 U2338 ( .A1(n332), .A2(n2124), .ZN(n326) );
  NAND2_X1 U2339 ( .A1(n709), .A2(n716), .ZN(n409) );
  INV_X1 U2340 ( .A(n746), .ZN(n747) );
  AOI21_X1 U2341 ( .B1(n595), .B2(n609), .A(n596), .ZN(n594) );
  NOR2_X1 U2342 ( .A1(n1171), .A2(n1174), .ZN(n633) );
  XNOR2_X1 U2343 ( .A(n504), .B(n317), .ZN(product[29]) );
  INV_X1 U2344 ( .A(n502), .ZN(n668) );
  INV_X1 U2345 ( .A(n2052), .ZN(n523) );
  NAND2_X1 U2346 ( .A1(n2052), .A2(n670), .ZN(n516) );
  INV_X1 U2347 ( .A(n534), .ZN(n672) );
  NAND2_X1 U2348 ( .A1(n525), .A2(n1982), .ZN(n505) );
  NAND2_X1 U2349 ( .A1(n1071), .A2(n1084), .ZN(n591) );
  XNOR2_X1 U2350 ( .A(b[17]), .B(n2260), .ZN(n1663) );
  XNOR2_X1 U2351 ( .A(b[19]), .B(n2260), .ZN(n1661) );
  XNOR2_X1 U2352 ( .A(b[15]), .B(n2260), .ZN(n1665) );
  XNOR2_X1 U2353 ( .A(b[21]), .B(n2260), .ZN(n1659) );
  XNOR2_X1 U2354 ( .A(b[11]), .B(n2260), .ZN(n1669) );
  XNOR2_X1 U2355 ( .A(b[13]), .B(n2260), .ZN(n1667) );
  OAI22_X1 U2356 ( .A1(n1781), .A2(n2235), .B1(n2220), .B2(n2076), .ZN(n1193)
         );
  OAI21_X1 U2357 ( .B1(n456), .B2(n481), .A(n457), .ZN(n455) );
  OAI21_X1 U2358 ( .B1(n503), .B2(n495), .A(n496), .ZN(n490) );
  OAI21_X1 U2359 ( .B1(n594), .B2(n582), .A(n583), .ZN(n581) );
  INV_X1 U2360 ( .A(n1931), .ZN(n524) );
  AOI21_X1 U2361 ( .B1(n1931), .B2(n670), .A(n519), .ZN(n517) );
  INV_X1 U2362 ( .A(n2196), .ZN(n508) );
  NOR2_X1 U2363 ( .A1(n542), .A2(n547), .ZN(n540) );
  OAI21_X1 U2364 ( .B1(n2194), .B2(n550), .A(n543), .ZN(n541) );
  OAI21_X1 U2365 ( .B1(n631), .B2(n634), .A(n632), .ZN(n630) );
  NAND2_X1 U2366 ( .A1(n1171), .A2(n1174), .ZN(n634) );
  NAND2_X1 U2367 ( .A1(n897), .A2(n918), .ZN(n535) );
  XNOR2_X1 U2368 ( .A(b[15]), .B(n1989), .ZN(n1640) );
  XNOR2_X1 U2369 ( .A(b[13]), .B(n2258), .ZN(n1642) );
  XNOR2_X1 U2370 ( .A(b[11]), .B(n2256), .ZN(n1644) );
  XNOR2_X1 U2371 ( .A(b[17]), .B(n2257), .ZN(n1638) );
  NAND2_X1 U2372 ( .A1(n663), .A2(n662), .ZN(n431) );
  NAND2_X1 U2373 ( .A1(n749), .A2(n760), .ZN(n439) );
  NOR2_X1 U2374 ( .A1(n749), .A2(n760), .ZN(n438) );
  INV_X1 U2375 ( .A(n772), .ZN(n773) );
  OAI22_X1 U2376 ( .A1(n2191), .A2(n1733), .B1(n1732), .B2(n2049), .ZN(n2198)
         );
  OAI22_X1 U2377 ( .A1(n2177), .A2(n1620), .B1(n1619), .B2(n2144), .ZN(n1326)
         );
  OAI22_X1 U2378 ( .A1(n2177), .A2(n1626), .B1(n1625), .B2(n1970), .ZN(n1332)
         );
  OAI22_X1 U2379 ( .A1(n2177), .A2(n1623), .B1(n2142), .B2(n1622), .ZN(n1329)
         );
  OAI22_X1 U2380 ( .A1(n2177), .A2(n1625), .B1(n1970), .B2(n1624), .ZN(n1331)
         );
  OAI22_X1 U2381 ( .A1(n2177), .A2(n1621), .B1(n1942), .B2(n1620), .ZN(n1327)
         );
  OAI22_X1 U2382 ( .A1(n1999), .A2(n1629), .B1(n1970), .B2(n1628), .ZN(n1335)
         );
  OAI22_X1 U2383 ( .A1(n2177), .A2(n1627), .B1(n1970), .B2(n1626), .ZN(n1333)
         );
  OAI22_X1 U2384 ( .A1(n287), .A2(n1619), .B1(n1942), .B2(n1618), .ZN(n1325)
         );
  OAI22_X1 U2385 ( .A1(n1999), .A2(n1624), .B1(n1623), .B2(n2142), .ZN(n1330)
         );
  AOI21_X1 U2386 ( .B1(n333), .B2(n2124), .A(n2125), .ZN(n327) );
  OAI21_X1 U2387 ( .B1(n337), .B2(n334), .A(n335), .ZN(n333) );
  OAI22_X1 U2388 ( .A1(n1972), .A2(n1483), .B1(n1482), .B2(n1986), .ZN(n676)
         );
  OAI22_X1 U2389 ( .A1(n1973), .A2(n1484), .B1(n1986), .B2(n1483), .ZN(n1195)
         );
  NAND2_X1 U2390 ( .A1(n717), .A2(n726), .ZN(n418) );
  OAI22_X1 U2391 ( .A1(n1972), .A2(n1485), .B1(n1484), .B2(n1986), .ZN(n1196)
         );
  OAI22_X1 U2392 ( .A1(n1972), .A2(n1491), .B1(n1490), .B2(n1986), .ZN(n1202)
         );
  OAI22_X1 U2393 ( .A1(n1973), .A2(n1488), .B1(n1986), .B2(n1487), .ZN(n1199)
         );
  OAI22_X1 U2394 ( .A1(n1972), .A2(n1487), .B1(n1486), .B2(n1986), .ZN(n1198)
         );
  OAI22_X1 U2395 ( .A1(n1973), .A2(n1486), .B1(n1986), .B2(n1485), .ZN(n1197)
         );
  OAI22_X1 U2396 ( .A1(n1973), .A2(n1490), .B1(n1986), .B2(n1489), .ZN(n1201)
         );
  OAI22_X1 U2397 ( .A1(n1972), .A2(n1489), .B1(n1488), .B2(n1986), .ZN(n1200)
         );
  OAI22_X1 U2398 ( .A1(n1506), .A2(n2221), .B1(n2204), .B2(n2237), .ZN(n1182)
         );
  OAI22_X1 U2399 ( .A1(n1492), .A2(n1973), .B1(n1986), .B2(n1491), .ZN(n1203)
         );
  OAI22_X1 U2400 ( .A1(n1973), .A2(n1493), .B1(n1492), .B2(n1986), .ZN(n1204)
         );
  OAI22_X1 U2401 ( .A1(n2193), .A2(n1695), .B1(n1694), .B2(n2228), .ZN(n1398)
         );
  OAI22_X1 U2402 ( .A1(n2193), .A2(n1704), .B1(n2002), .B2(n1703), .ZN(n1407)
         );
  OAI22_X1 U2403 ( .A1(n2193), .A2(n1701), .B1(n1700), .B2(n2228), .ZN(n1404)
         );
  OAI22_X1 U2404 ( .A1(n2193), .A2(n1702), .B1(n2228), .B2(n1701), .ZN(n1405)
         );
  OAI22_X1 U2405 ( .A1(n2193), .A2(n1698), .B1(n2228), .B2(n1697), .ZN(n1401)
         );
  OAI22_X1 U2406 ( .A1(n2193), .A2(n1705), .B1(n1704), .B2(n2228), .ZN(n1408)
         );
  OAI22_X1 U2407 ( .A1(n2193), .A2(n1694), .B1(n2228), .B2(n1693), .ZN(n1397)
         );
  OAI22_X1 U2408 ( .A1(n2193), .A2(n1696), .B1(n2002), .B2(n1695), .ZN(n1399)
         );
  OAI22_X1 U2409 ( .A1(n2193), .A2(n1700), .B1(n2228), .B2(n1699), .ZN(n1403)
         );
  OAI22_X1 U2410 ( .A1(n2096), .A2(n1699), .B1(n1698), .B2(n2228), .ZN(n1402)
         );
  OAI22_X1 U2411 ( .A1(n2193), .A2(n1703), .B1(n1702), .B2(n2228), .ZN(n1406)
         );
  OAI22_X1 U2412 ( .A1(n2096), .A2(n1697), .B1(n1696), .B2(n2228), .ZN(n1400)
         );
  NAND2_X1 U2413 ( .A1(n1814), .A2(n257), .ZN(n281) );
  INV_X1 U2414 ( .A(n513), .ZN(n669) );
  NOR2_X1 U2415 ( .A1(n513), .A2(n520), .ZN(n511) );
  OAI21_X1 U2416 ( .B1(n2147), .B2(n521), .A(n514), .ZN(n512) );
  XNOR2_X1 U2417 ( .A(n2035), .B(n1237), .ZN(n939) );
  OR2_X1 U2418 ( .A1(n1215), .A2(n1237), .ZN(n938) );
  NAND2_X1 U2419 ( .A1(n1165), .A2(n1170), .ZN(n632) );
  XNOR2_X1 U2420 ( .A(b[21]), .B(n1997), .ZN(n1559) );
  XNOR2_X1 U2421 ( .A(b[15]), .B(n2247), .ZN(n1565) );
  XNOR2_X1 U2422 ( .A(b[11]), .B(n1998), .ZN(n1569) );
  XNOR2_X1 U2423 ( .A(b[17]), .B(n2247), .ZN(n1563) );
  XNOR2_X1 U2424 ( .A(b[13]), .B(n2247), .ZN(n1567) );
  XNOR2_X1 U2425 ( .A(b[19]), .B(n2245), .ZN(n1561) );
  XNOR2_X1 U2426 ( .A(b[17]), .B(n1976), .ZN(n1588) );
  XNOR2_X1 U2427 ( .A(b[13]), .B(n1976), .ZN(n1592) );
  XNOR2_X1 U2428 ( .A(b[15]), .B(n2249), .ZN(n1590) );
  XNOR2_X1 U2429 ( .A(b[19]), .B(n2249), .ZN(n1586) );
  XNOR2_X1 U2430 ( .A(b[21]), .B(n1977), .ZN(n1584) );
  XNOR2_X1 U2431 ( .A(b[11]), .B(n1976), .ZN(n1594) );
  AOI21_X1 U2432 ( .B1(n540), .B2(n553), .A(n541), .ZN(n539) );
  NAND2_X1 U2433 ( .A1(n2033), .A2(n552), .ZN(n538) );
  AOI21_X1 U2434 ( .B1(n508), .B2(n465), .A(n466), .ZN(n464) );
  AOI21_X1 U2435 ( .B1(n508), .B2(n668), .A(n501), .ZN(n499) );
  AOI21_X1 U2436 ( .B1(n508), .B2(n478), .A(n479), .ZN(n477) );
  AOI21_X1 U2437 ( .B1(n508), .B2(n2156), .A(n2160), .ZN(n488) );
  NAND2_X1 U2438 ( .A1(n1372), .A2(n1284), .ZN(n2199) );
  NAND2_X1 U2439 ( .A1(n1284), .A2(n1438), .ZN(n2200) );
  NAND2_X1 U2440 ( .A1(n1372), .A2(n1438), .ZN(n2201) );
  NAND3_X1 U2441 ( .A1(n2199), .A2(n2200), .A3(n2201), .ZN(n996) );
  AOI21_X1 U2442 ( .B1(n2054), .B2(n2188), .A(n451), .ZN(n2203) );
  AOI21_X1 U2443 ( .B1(n2054), .B2(n2188), .A(n451), .ZN(n2202) );
  AOI21_X1 U2444 ( .B1(n537), .B2(n2188), .A(n451), .ZN(n301) );
  NAND2_X1 U2445 ( .A1(n1953), .A2(n378), .ZN(n305) );
  NAND2_X1 U2446 ( .A1(n382), .A2(n1953), .ZN(n371) );
  AOI21_X1 U2447 ( .B1(n383), .B2(n1953), .A(n376), .ZN(n372) );
  NAND2_X1 U2448 ( .A1(n345), .A2(n2123), .ZN(n336) );
  NAND2_X1 U2449 ( .A1(n1953), .A2(n2121), .ZN(n364) );
  OAI21_X1 U2450 ( .B1(n421), .B2(n402), .A(n405), .ZN(n401) );
  OAI21_X1 U2451 ( .B1(n428), .B2(n436), .A(n429), .ZN(n427) );
  XNOR2_X1 U2452 ( .A(n437), .B(n311), .ZN(product[35]) );
  NAND2_X1 U2453 ( .A1(n805), .A2(n820), .ZN(n496) );
  XNOR2_X1 U2454 ( .A(b[17]), .B(n2278), .ZN(n1763) );
  XNOR2_X1 U2455 ( .A(b[13]), .B(n2280), .ZN(n1767) );
  XNOR2_X1 U2456 ( .A(b[21]), .B(n2280), .ZN(n1759) );
  XNOR2_X1 U2457 ( .A(b[15]), .B(n2279), .ZN(n1765) );
  XNOR2_X1 U2458 ( .A(b[11]), .B(n2278), .ZN(n1769) );
  XNOR2_X1 U2459 ( .A(b[19]), .B(n2279), .ZN(n1761) );
  XNOR2_X1 U2460 ( .A(n430), .B(n310), .ZN(product[36]) );
  OAI22_X1 U2461 ( .A1(n2014), .A2(n1637), .B1(n1636), .B2(n2146), .ZN(n1342)
         );
  OAI22_X1 U2462 ( .A1(n2015), .A2(n1635), .B1(n1634), .B2(n2146), .ZN(n1340)
         );
  OAI22_X1 U2463 ( .A1(n2014), .A2(n1652), .B1(n2226), .B2(n1651), .ZN(n1357)
         );
  OAI22_X1 U2464 ( .A1(n2015), .A2(n1649), .B1(n1648), .B2(n2226), .ZN(n1354)
         );
  OAI22_X1 U2465 ( .A1(n2015), .A2(n1653), .B1(n1652), .B2(n2146), .ZN(n1358)
         );
  OAI22_X1 U2466 ( .A1(n2015), .A2(n1648), .B1(n2226), .B2(n1647), .ZN(n1353)
         );
  OAI22_X1 U2467 ( .A1(n2213), .A2(n1639), .B1(n1638), .B2(n2146), .ZN(n1344)
         );
  OAI22_X1 U2468 ( .A1(n2015), .A2(n1647), .B1(n1646), .B2(n2226), .ZN(n1352)
         );
  OAI22_X1 U2469 ( .A1(n2014), .A2(n1654), .B1(n2226), .B2(n1653), .ZN(n1359)
         );
  OAI22_X1 U2470 ( .A1(n2015), .A2(n1650), .B1(n2226), .B2(n1649), .ZN(n1355)
         );
  OAI22_X1 U2471 ( .A1(n2015), .A2(n1645), .B1(n1644), .B2(n2226), .ZN(n1350)
         );
  OAI22_X1 U2472 ( .A1(n2213), .A2(n1655), .B1(n1654), .B2(n2146), .ZN(n1360)
         );
  OAI22_X1 U2473 ( .A1(n2014), .A2(n1641), .B1(n1640), .B2(n2146), .ZN(n1346)
         );
  OAI22_X1 U2474 ( .A1(n2014), .A2(n1644), .B1(n2146), .B2(n1643), .ZN(n1349)
         );
  OAI22_X1 U2475 ( .A1(n1656), .A2(n2146), .B1(n2014), .B2(n2259), .ZN(n1188)
         );
  OAI22_X1 U2476 ( .A1(n2015), .A2(n1633), .B1(n1632), .B2(n2146), .ZN(n772)
         );
  OAI22_X1 U2477 ( .A1(n2015), .A2(n1643), .B1(n1642), .B2(n2146), .ZN(n1348)
         );
  OAI22_X1 U2478 ( .A1(n2213), .A2(n1651), .B1(n1650), .B2(n2226), .ZN(n1356)
         );
  OAI22_X1 U2479 ( .A1(n2014), .A2(n1646), .B1(n2146), .B2(n1645), .ZN(n1351)
         );
  OAI22_X1 U2480 ( .A1(n1756), .A2(n2233), .B1(n2191), .B2(n2011), .ZN(n1192)
         );
  OAI22_X1 U2481 ( .A1(n2190), .A2(n1738), .B1(n2233), .B2(n1737), .ZN(n1439)
         );
  OAI22_X1 U2482 ( .A1(n2195), .A2(n1741), .B1(n1740), .B2(n2049), .ZN(n1442)
         );
  OAI22_X1 U2483 ( .A1(n2191), .A2(n1740), .B1(n2233), .B2(n1739), .ZN(n1441)
         );
  OAI22_X1 U2484 ( .A1(n2195), .A2(n1735), .B1(n1734), .B2(n2233), .ZN(n1436)
         );
  OAI22_X1 U2485 ( .A1(n2195), .A2(n1739), .B1(n1738), .B2(n2049), .ZN(n1440)
         );
  OAI22_X1 U2486 ( .A1(n2195), .A2(n1742), .B1(n2233), .B2(n1741), .ZN(n1443)
         );
  OAI22_X1 U2487 ( .A1(n2195), .A2(n1734), .B1(n2049), .B2(n1733), .ZN(n1435)
         );
  OAI22_X1 U2488 ( .A1(n2190), .A2(n1736), .B1(n2049), .B2(n1735), .ZN(n1437)
         );
  OAI22_X1 U2489 ( .A1(n2195), .A2(n1737), .B1(n1736), .B2(n2048), .ZN(n1438)
         );
  OAI22_X1 U2490 ( .A1(n2195), .A2(n1743), .B1(n1742), .B2(n2048), .ZN(n1444)
         );
  XNOR2_X1 U2491 ( .A(n419), .B(n309), .ZN(product[37]) );
  OAI22_X1 U2492 ( .A1(n2098), .A2(n1508), .B1(n1507), .B2(n2001), .ZN(n682)
         );
  OAI22_X1 U2493 ( .A1(n2187), .A2(n1518), .B1(n1517), .B2(n2001), .ZN(n1228)
         );
  OAI22_X1 U2494 ( .A1(n2187), .A2(n1522), .B1(n1521), .B2(n2038), .ZN(n1232)
         );
  OAI22_X1 U2495 ( .A1(n2187), .A2(n1510), .B1(n1509), .B2(n2001), .ZN(n1220)
         );
  OAI22_X1 U2496 ( .A1(n2187), .A2(n1521), .B1(n2038), .B2(n1520), .ZN(n1231)
         );
  OAI22_X1 U2497 ( .A1(n2187), .A2(n1519), .B1(n2038), .B2(n1518), .ZN(n1229)
         );
  OAI22_X1 U2498 ( .A1(n2187), .A2(n1514), .B1(n1513), .B2(n2001), .ZN(n1224)
         );
  OAI22_X1 U2499 ( .A1(n2187), .A2(n1520), .B1(n1519), .B2(n2038), .ZN(n1230)
         );
  OAI22_X1 U2500 ( .A1(n2187), .A2(n1512), .B1(n1511), .B2(n2001), .ZN(n1222)
         );
  OAI22_X1 U2501 ( .A1(n2187), .A2(n1525), .B1(n2038), .B2(n1524), .ZN(n1235)
         );
  OAI22_X1 U2502 ( .A1(n2187), .A2(n1523), .B1(n2038), .B2(n1522), .ZN(n1233)
         );
  OAI22_X1 U2503 ( .A1(n2206), .A2(n1526), .B1(n1525), .B2(n2038), .ZN(n1236)
         );
  OAI22_X1 U2504 ( .A1(n1531), .A2(n2001), .B1(n2187), .B2(n1968), .ZN(n1183)
         );
  OAI22_X1 U2505 ( .A1(n1524), .A2(n2179), .B1(n1523), .B2(n2038), .ZN(n1234)
         );
  OAI22_X1 U2506 ( .A1(n2206), .A2(n1528), .B1(n1527), .B2(n2038), .ZN(n1238)
         );
  OAI22_X1 U2507 ( .A1(n2187), .A2(n1516), .B1(n1515), .B2(n2001), .ZN(n1226)
         );
  OAI22_X1 U2508 ( .A1(n2179), .A2(n1529), .B1(n2038), .B2(n1528), .ZN(n1239)
         );
  OAI22_X1 U2509 ( .A1(n2179), .A2(n1527), .B1(n2038), .B2(n1526), .ZN(n1237)
         );
  OAI22_X1 U2510 ( .A1(n2206), .A2(n1530), .B1(n1529), .B2(n2038), .ZN(n1240)
         );
  NAND2_X1 U2511 ( .A1(n1807), .A2(n2095), .ZN(n295) );
  NAND2_X1 U2512 ( .A1(n465), .A2(n507), .ZN(n463) );
  NAND2_X1 U2513 ( .A1(n507), .A2(n668), .ZN(n498) );
  NAND2_X1 U2514 ( .A1(n507), .A2(n2156), .ZN(n487) );
  NAND2_X1 U2515 ( .A1(n478), .A2(n507), .ZN(n476) );
  OAI22_X1 U2516 ( .A1(n1987), .A2(n1571), .B1(n2223), .B2(n1570), .ZN(n1279)
         );
  OAI22_X1 U2517 ( .A1(n1929), .A2(n1580), .B1(n1579), .B2(n2222), .ZN(n1288)
         );
  OAI22_X1 U2518 ( .A1(n1929), .A2(n1570), .B1(n1569), .B2(n2223), .ZN(n1278)
         );
  OAI22_X1 U2519 ( .A1(n2040), .A2(n1573), .B1(n2222), .B2(n1572), .ZN(n1281)
         );
  OAI22_X1 U2520 ( .A1(n1987), .A2(n1579), .B1(n2222), .B2(n1578), .ZN(n1287)
         );
  OAI22_X1 U2521 ( .A1(n1929), .A2(n1575), .B1(n2222), .B2(n1574), .ZN(n1283)
         );
  OAI22_X1 U2522 ( .A1(n2040), .A2(n1569), .B1(n2222), .B2(n1568), .ZN(n1277)
         );
  OAI22_X1 U2523 ( .A1(n2040), .A2(n1572), .B1(n1571), .B2(n2223), .ZN(n1280)
         );
  OAI22_X1 U2524 ( .A1(n2040), .A2(n1578), .B1(n1577), .B2(n2222), .ZN(n1286)
         );
  OAI22_X1 U2525 ( .A1(n2040), .A2(n1574), .B1(n1573), .B2(n2223), .ZN(n1282)
         );
  OAI22_X1 U2526 ( .A1(n2040), .A2(n1577), .B1(n2222), .B2(n1576), .ZN(n1285)
         );
  OAI22_X1 U2527 ( .A1(n1929), .A2(n1576), .B1(n1575), .B2(n2222), .ZN(n1284)
         );
  XNOR2_X1 U2528 ( .A(n410), .B(n308), .ZN(product[38]) );
  OAI22_X1 U2529 ( .A1(n2190), .A2(n1753), .B1(n1752), .B2(n2233), .ZN(n1454)
         );
  OAI22_X1 U2530 ( .A1(n2191), .A2(n1747), .B1(n1746), .B2(n2233), .ZN(n1448)
         );
  OAI22_X1 U2531 ( .A1(n2190), .A2(n1750), .B1(n2049), .B2(n1749), .ZN(n1451)
         );
  OAI22_X1 U2532 ( .A1(n2191), .A2(n1749), .B1(n1748), .B2(n2049), .ZN(n1450)
         );
  OAI22_X1 U2533 ( .A1(n2191), .A2(n1745), .B1(n1744), .B2(n2233), .ZN(n1446)
         );
  OAI22_X1 U2534 ( .A1(n2190), .A2(n1748), .B1(n2049), .B2(n1747), .ZN(n1449)
         );
  OAI22_X1 U2535 ( .A1(n2195), .A2(n1744), .B1(n2233), .B2(n1743), .ZN(n1445)
         );
  OAI22_X1 U2536 ( .A1(n2195), .A2(n1746), .B1(n2049), .B2(n1745), .ZN(n1447)
         );
  OAI22_X1 U2537 ( .A1(n2191), .A2(n1754), .B1(n2049), .B2(n1753), .ZN(n1455)
         );
  OAI22_X1 U2538 ( .A1(n2190), .A2(n1752), .B1(n2049), .B2(n1751), .ZN(n1453)
         );
  OAI22_X1 U2539 ( .A1(n2195), .A2(n1751), .B1(n1750), .B2(n2233), .ZN(n1452)
         );
  OAI22_X1 U2540 ( .A1(n2195), .A2(n1755), .B1(n1754), .B2(n2233), .ZN(n1456)
         );
  XNOR2_X1 U2541 ( .A(n397), .B(n307), .ZN(product[39]) );
  OAI22_X1 U2542 ( .A1(n2063), .A2(n1661), .B1(n2037), .B2(n1660), .ZN(n1365)
         );
  OAI22_X1 U2543 ( .A1(n2063), .A2(n1660), .B1(n1659), .B2(n1981), .ZN(n1364)
         );
  OAI22_X1 U2544 ( .A1(n2063), .A2(n1663), .B1(n2227), .B2(n1662), .ZN(n1367)
         );
  OAI22_X1 U2545 ( .A1(n1681), .A2(n1981), .B1(n2062), .B2(n2264), .ZN(n1189)
         );
  OAI22_X1 U2546 ( .A1(n2062), .A2(n1664), .B1(n1663), .B2(n1981), .ZN(n1368)
         );
  OAI22_X1 U2547 ( .A1(n2062), .A2(n1665), .B1(n2227), .B2(n1664), .ZN(n1369)
         );
  OAI22_X1 U2548 ( .A1(n2062), .A2(n1658), .B1(n1657), .B2(n1981), .ZN(n802)
         );
  OAI22_X1 U2549 ( .A1(n2063), .A2(n1667), .B1(n2227), .B2(n1666), .ZN(n1371)
         );
  OAI22_X1 U2550 ( .A1(n2070), .A2(n1662), .B1(n1661), .B2(n1981), .ZN(n1366)
         );
  OAI22_X1 U2551 ( .A1(n2063), .A2(n1666), .B1(n1665), .B2(n1981), .ZN(n1370)
         );
  XNOR2_X1 U2552 ( .A(b[17]), .B(n2267), .ZN(n1688) );
  OAI22_X1 U2553 ( .A1(n2070), .A2(n1659), .B1(n2227), .B2(n1658), .ZN(n1363)
         );
  XNOR2_X1 U2554 ( .A(b[19]), .B(n2268), .ZN(n1686) );
  XNOR2_X1 U2555 ( .A(b[11]), .B(n2266), .ZN(n1694) );
  XNOR2_X1 U2556 ( .A(b[21]), .B(n2266), .ZN(n1684) );
  XNOR2_X1 U2557 ( .A(b[15]), .B(n2268), .ZN(n1690) );
  XNOR2_X1 U2558 ( .A(b[13]), .B(n2266), .ZN(n1692) );
  XNOR2_X1 U2559 ( .A(n388), .B(n306), .ZN(product[40]) );
  OAI22_X1 U2560 ( .A1(n2062), .A2(n1671), .B1(n2227), .B2(n1670), .ZN(n1375)
         );
  OAI22_X1 U2561 ( .A1(n2063), .A2(n1672), .B1(n1671), .B2(n2227), .ZN(n1376)
         );
  OAI22_X1 U2562 ( .A1(n2062), .A2(n1679), .B1(n2227), .B2(n1678), .ZN(n1383)
         );
  OAI22_X1 U2563 ( .A1(n2062), .A2(n1677), .B1(n2227), .B2(n1676), .ZN(n1381)
         );
  OAI22_X1 U2564 ( .A1(n2062), .A2(n1675), .B1(n2227), .B2(n1674), .ZN(n1379)
         );
  OAI22_X1 U2565 ( .A1(n2070), .A2(n1669), .B1(n2227), .B2(n1668), .ZN(n1373)
         );
  OAI22_X1 U2566 ( .A1(n2063), .A2(n1676), .B1(n1675), .B2(n2227), .ZN(n1380)
         );
  OAI22_X1 U2567 ( .A1(n2063), .A2(n1670), .B1(n1669), .B2(n2227), .ZN(n1374)
         );
  OAI22_X1 U2568 ( .A1(n2062), .A2(n1680), .B1(n1679), .B2(n1981), .ZN(n1384)
         );
  OAI22_X1 U2569 ( .A1(n2062), .A2(n1678), .B1(n1677), .B2(n1981), .ZN(n1382)
         );
  OAI22_X1 U2570 ( .A1(n2062), .A2(n1674), .B1(n1673), .B2(n2227), .ZN(n1378)
         );
  OAI22_X1 U2571 ( .A1(n2063), .A2(n1673), .B1(n2227), .B2(n1672), .ZN(n1377)
         );
  OAI22_X1 U2572 ( .A1(n1731), .A2(n2141), .B1(n2217), .B2(n2273), .ZN(n1191)
         );
  OAI22_X1 U2573 ( .A1(n2216), .A2(n1718), .B1(n1717), .B2(n2141), .ZN(n1420)
         );
  OAI22_X1 U2574 ( .A1(n2069), .A2(n1711), .B1(n2231), .B2(n1710), .ZN(n1413)
         );
  OAI22_X1 U2575 ( .A1(n2217), .A2(n1717), .B1(n2231), .B2(n1716), .ZN(n1419)
         );
  OAI22_X1 U2576 ( .A1(n2069), .A2(n1713), .B1(n2231), .B2(n1712), .ZN(n1415)
         );
  OAI22_X1 U2577 ( .A1(n2217), .A2(n1709), .B1(n2231), .B2(n1708), .ZN(n1411)
         );
  OAI22_X1 U2578 ( .A1(n2069), .A2(n1710), .B1(n1709), .B2(n2141), .ZN(n1412)
         );
  OAI22_X1 U2579 ( .A1(n2216), .A2(n1715), .B1(n2231), .B2(n1714), .ZN(n1417)
         );
  OAI22_X1 U2580 ( .A1(n2216), .A2(n1716), .B1(n1715), .B2(n2141), .ZN(n1418)
         );
  OAI22_X1 U2581 ( .A1(n2216), .A2(n1708), .B1(n1707), .B2(n2141), .ZN(n874)
         );
  OAI22_X1 U2582 ( .A1(n2216), .A2(n1714), .B1(n1713), .B2(n2141), .ZN(n1416)
         );
  OAI22_X1 U2583 ( .A1(n2217), .A2(n1712), .B1(n1711), .B2(n2141), .ZN(n1414)
         );
  XNOR2_X1 U2584 ( .A(b[11]), .B(n2274), .ZN(n1744) );
  XNOR2_X1 U2585 ( .A(b[21]), .B(n2275), .ZN(n1734) );
  XNOR2_X1 U2586 ( .A(b[15]), .B(n2276), .ZN(n1740) );
  XNOR2_X1 U2587 ( .A(b[19]), .B(n2274), .ZN(n1736) );
  XNOR2_X1 U2588 ( .A(b[17]), .B(n2274), .ZN(n1738) );
  XNOR2_X1 U2589 ( .A(b[13]), .B(n2276), .ZN(n1742) );
  XNOR2_X1 U2590 ( .A(n379), .B(n305), .ZN(product[41]) );
  INV_X1 U2591 ( .A(n916), .ZN(n917) );
  OAI21_X1 U2592 ( .B1(n421), .B2(n347), .A(n348), .ZN(n346) );
  OAI22_X1 U2593 ( .A1(n2177), .A2(n1613), .B1(n1942), .B2(n1612), .ZN(n1319)
         );
  OAI22_X1 U2594 ( .A1(n1999), .A2(n1612), .B1(n1611), .B2(n2143), .ZN(n1318)
         );
  OAI22_X1 U2595 ( .A1(n1999), .A2(n1617), .B1(n1970), .B2(n1616), .ZN(n1323)
         );
  OAI22_X1 U2596 ( .A1(n1999), .A2(n1630), .B1(n1629), .B2(n2144), .ZN(n1336)
         );
  OAI22_X1 U2597 ( .A1(n1631), .A2(n2143), .B1(n1999), .B2(n1988), .ZN(n1187)
         );
  OAI22_X1 U2598 ( .A1(n1999), .A2(n1611), .B1(n1942), .B2(n1610), .ZN(n1317)
         );
  OAI22_X1 U2599 ( .A1(n2177), .A2(n1610), .B1(n1609), .B2(n2144), .ZN(n1316)
         );
  OAI22_X1 U2600 ( .A1(n1999), .A2(n1615), .B1(n1970), .B2(n1614), .ZN(n1321)
         );
  OAI22_X1 U2601 ( .A1(n1999), .A2(n1609), .B1(n1942), .B2(n1608), .ZN(n1315)
         );
  OAI22_X1 U2602 ( .A1(n1999), .A2(n1618), .B1(n1617), .B2(n2144), .ZN(n1324)
         );
  OAI22_X1 U2603 ( .A1(n2180), .A2(n1616), .B1(n1615), .B2(n2143), .ZN(n1322)
         );
  OAI22_X1 U2604 ( .A1(n2177), .A2(n1608), .B1(n1607), .B2(n2143), .ZN(n746)
         );
  OAI22_X1 U2605 ( .A1(n2177), .A2(n1628), .B1(n1627), .B2(n2143), .ZN(n1334)
         );
  NAND2_X1 U2606 ( .A1(n2142), .A2(n1811), .ZN(n287) );
  XNOR2_X1 U2607 ( .A(n370), .B(n304), .ZN(product[42]) );
  OAI22_X1 U2608 ( .A1(n2169), .A2(n1535), .B1(n1534), .B2(n2088), .ZN(n1244)
         );
  OAI22_X1 U2609 ( .A1(n2209), .A2(n1537), .B1(n1536), .B2(n2087), .ZN(n1246)
         );
  OAI22_X1 U2610 ( .A1(n2209), .A2(n1543), .B1(n1542), .B2(n2089), .ZN(n1252)
         );
  OAI22_X1 U2611 ( .A1(n1556), .A2(n2088), .B1(n2208), .B2(n1945), .ZN(n1184)
         );
  OAI22_X1 U2612 ( .A1(n2169), .A2(n1533), .B1(n1532), .B2(n2088), .ZN(n692)
         );
  OAI22_X1 U2613 ( .A1(n2208), .A2(n1541), .B1(n1540), .B2(n2089), .ZN(n1250)
         );
  OAI22_X1 U2614 ( .A1(n2209), .A2(n1539), .B1(n1538), .B2(n2089), .ZN(n1248)
         );
  NAND2_X1 U2615 ( .A1(n2034), .A2(n474), .ZN(n314) );
  AOI21_X1 U2616 ( .B1(n2034), .B2(n483), .A(n2036), .ZN(n468) );
  NAND2_X1 U2617 ( .A1(n666), .A2(n2034), .ZN(n467) );
  OAI22_X1 U2618 ( .A1(n1973), .A2(n1497), .B1(n1496), .B2(n1986), .ZN(n1208)
         );
  OAI22_X1 U2619 ( .A1(n1973), .A2(n1496), .B1(n1986), .B2(n1495), .ZN(n1207)
         );
  OAI22_X1 U2620 ( .A1(n1502), .A2(n1971), .B1(n1986), .B2(n1501), .ZN(n1213)
         );
  OAI22_X1 U2621 ( .A1(n1972), .A2(n1495), .B1(n1494), .B2(n1986), .ZN(n1206)
         );
  OAI22_X1 U2622 ( .A1(n1971), .A2(n1501), .B1(n1500), .B2(n2221), .ZN(n1212)
         );
  OAI22_X1 U2623 ( .A1(n2204), .A2(n1505), .B1(n1504), .B2(n2221), .ZN(n1216)
         );
  OAI22_X1 U2624 ( .A1(n1972), .A2(n1494), .B1(n1986), .B2(n1493), .ZN(n1205)
         );
  OAI22_X1 U2625 ( .A1(n2172), .A2(n1503), .B1(n1502), .B2(n2221), .ZN(n1214)
         );
  OAI22_X1 U2626 ( .A1(n1972), .A2(n1500), .B1(n1986), .B2(n1499), .ZN(n1211)
         );
  OAI22_X1 U2627 ( .A1(n2172), .A2(n1504), .B1(n2221), .B2(n1503), .ZN(n1215)
         );
  OAI22_X1 U2628 ( .A1(n2172), .A2(n1498), .B1(n2221), .B2(n1497), .ZN(n1209)
         );
  OAI22_X1 U2629 ( .A1(n2204), .A2(n1499), .B1(n1498), .B2(n2221), .ZN(n1210)
         );
  XNOR2_X1 U2630 ( .A(b[21]), .B(n2140), .ZN(n1509) );
  XNOR2_X1 U2631 ( .A(b[17]), .B(n2140), .ZN(n1513) );
  XNOR2_X1 U2632 ( .A(b[11]), .B(n2239), .ZN(n1519) );
  XNOR2_X1 U2633 ( .A(b[19]), .B(n2239), .ZN(n1511) );
  XNOR2_X1 U2634 ( .A(b[13]), .B(n2140), .ZN(n1517) );
  XNOR2_X1 U2635 ( .A(b[15]), .B(n2239), .ZN(n1515) );
  OAI22_X1 U2636 ( .A1(n2070), .A2(n1668), .B1(n1667), .B2(n1981), .ZN(n1372)
         );
  XNOR2_X1 U2637 ( .A(a[6]), .B(a[5]), .ZN(n257) );
  XNOR2_X1 U2638 ( .A(b[17]), .B(n2270), .ZN(n1713) );
  XNOR2_X1 U2639 ( .A(b[19]), .B(n2272), .ZN(n1711) );
  XNOR2_X1 U2640 ( .A(b[15]), .B(n2271), .ZN(n1715) );
  XNOR2_X1 U2641 ( .A(b[11]), .B(n2270), .ZN(n1719) );
  XNOR2_X1 U2642 ( .A(b[21]), .B(n2270), .ZN(n1709) );
  XNOR2_X1 U2643 ( .A(n353), .B(n303), .ZN(product[43]) );
  OAI22_X1 U2644 ( .A1(n2209), .A2(n1544), .B1(n2089), .B2(n1543), .ZN(n1253)
         );
  OAI22_X1 U2645 ( .A1(n2169), .A2(n1552), .B1(n2088), .B2(n1551), .ZN(n1261)
         );
  OAI22_X1 U2646 ( .A1(n2208), .A2(n1549), .B1(n1548), .B2(n2087), .ZN(n1258)
         );
  OAI22_X1 U2647 ( .A1(n2168), .A2(n1548), .B1(n2089), .B2(n1547), .ZN(n1257)
         );
  OAI22_X1 U2648 ( .A1(n2209), .A2(n1555), .B1(n1554), .B2(n2088), .ZN(n1264)
         );
  OAI22_X1 U2649 ( .A1(n2168), .A2(n1547), .B1(n1546), .B2(n2089), .ZN(n1256)
         );
  OAI22_X1 U2650 ( .A1(n2169), .A2(n1546), .B1(n2087), .B2(n1545), .ZN(n1255)
         );
  OAI22_X1 U2651 ( .A1(n2169), .A2(n1550), .B1(n2087), .B2(n1549), .ZN(n1259)
         );
  OAI22_X1 U2652 ( .A1(n2169), .A2(n1545), .B1(n1544), .B2(n2087), .ZN(n1254)
         );
  OAI22_X1 U2653 ( .A1(n2168), .A2(n1554), .B1(n2088), .B2(n1553), .ZN(n1263)
         );
  OAI22_X1 U2654 ( .A1(n2209), .A2(n1551), .B1(n1550), .B2(n2087), .ZN(n1260)
         );
  OAI22_X1 U2655 ( .A1(n2168), .A2(n1553), .B1(n1552), .B2(n2088), .ZN(n1262)
         );
  INV_X1 U2656 ( .A(n346), .ZN(n344) );
  AOI21_X1 U2657 ( .B1(n346), .B2(n2123), .A(n339), .ZN(n337) );
  NAND2_X1 U2658 ( .A1(n694), .A2(n689), .ZN(n378) );
  OAI22_X1 U2659 ( .A1(n2210), .A2(n1602), .B1(n1965), .B2(n1601), .ZN(n1309)
         );
  OAI22_X1 U2660 ( .A1(n2003), .A2(n1600), .B1(n1965), .B2(n1599), .ZN(n1307)
         );
  OAI22_X1 U2661 ( .A1(n2210), .A2(n1601), .B1(n1600), .B2(n1965), .ZN(n1308)
         );
  OAI22_X1 U2662 ( .A1(n2211), .A2(n1594), .B1(n1964), .B2(n1593), .ZN(n1301)
         );
  OAI22_X1 U2663 ( .A1(n2211), .A2(n1596), .B1(n1964), .B2(n1595), .ZN(n1303)
         );
  OAI22_X1 U2664 ( .A1(n2004), .A2(n1598), .B1(n1965), .B2(n1597), .ZN(n1305)
         );
  OAI22_X1 U2665 ( .A1(n2004), .A2(n1595), .B1(n1594), .B2(n1964), .ZN(n1302)
         );
  OAI22_X1 U2666 ( .A1(n2210), .A2(n1597), .B1(n1596), .B2(n1965), .ZN(n1304)
         );
  OAI22_X1 U2667 ( .A1(n2003), .A2(n1603), .B1(n1602), .B2(n1965), .ZN(n1310)
         );
  OAI22_X1 U2668 ( .A1(n2003), .A2(n1604), .B1(n1965), .B2(n1603), .ZN(n1311)
         );
  OAI22_X1 U2669 ( .A1(n2210), .A2(n1599), .B1(n1598), .B2(n1965), .ZN(n1306)
         );
  OAI22_X1 U2670 ( .A1(n2211), .A2(n1605), .B1(n1604), .B2(n1964), .ZN(n1312)
         );
  XNOR2_X1 U2671 ( .A(b[19]), .B(n2254), .ZN(n1611) );
  XNOR2_X1 U2672 ( .A(b[11]), .B(n2253), .ZN(n1619) );
  XNOR2_X1 U2673 ( .A(b[17]), .B(n2254), .ZN(n1613) );
  XNOR2_X1 U2674 ( .A(b[13]), .B(n2253), .ZN(n1617) );
  XNOR2_X1 U2675 ( .A(b[21]), .B(n2253), .ZN(n1609) );
  XNOR2_X1 U2676 ( .A(b[15]), .B(n2253), .ZN(n1615) );
  NAND2_X1 U2677 ( .A1(n489), .A2(n454), .ZN(n452) );
  AOI21_X1 U2678 ( .B1(n490), .B2(n454), .A(n455), .ZN(n453) );
  OAI22_X1 U2679 ( .A1(n2195), .A2(n1733), .B1(n1732), .B2(n2233), .ZN(n916)
         );
  OAI21_X1 U2680 ( .B1(n506), .B2(n452), .A(n453), .ZN(n451) );
  XNOR2_X1 U2681 ( .A(n462), .B(n313), .ZN(product[33]) );
  XOR2_X1 U2682 ( .A(n1992), .B(n321), .Z(product[25]) );
  OAI21_X1 U2683 ( .B1(n1993), .B2(n516), .A(n517), .ZN(n515) );
  OAI21_X1 U2684 ( .B1(n1991), .B2(n523), .A(n524), .ZN(n522) );
  OAI21_X1 U2685 ( .B1(n1993), .B2(n463), .A(n464), .ZN(n462) );
  OAI21_X1 U2686 ( .B1(n1991), .B2(n2159), .A(n2174), .ZN(n533) );
  OAI21_X1 U2687 ( .B1(n1991), .B2(n476), .A(n477), .ZN(n475) );
  OAI21_X1 U2688 ( .B1(n1992), .B2(n487), .A(n488), .ZN(n486) );
  OAI21_X1 U2689 ( .B1(n1992), .B2(n498), .A(n499), .ZN(n497) );
  OAI21_X1 U2690 ( .B1(n1993), .B2(n505), .A(n2197), .ZN(n504) );
  OAI22_X1 U2691 ( .A1(n2069), .A2(n1727), .B1(n2141), .B2(n1726), .ZN(n1429)
         );
  OAI22_X1 U2692 ( .A1(n2217), .A2(n1720), .B1(n1719), .B2(n2231), .ZN(n1422)
         );
  OAI22_X1 U2693 ( .A1(n2216), .A2(n1721), .B1(n2231), .B2(n1720), .ZN(n1423)
         );
  OAI22_X1 U2694 ( .A1(n2217), .A2(n1726), .B1(n1725), .B2(n2231), .ZN(n1428)
         );
  OAI22_X1 U2695 ( .A1(n2217), .A2(n1730), .B1(n1729), .B2(n2141), .ZN(n1432)
         );
  OAI22_X1 U2696 ( .A1(n2069), .A2(n1725), .B1(n2231), .B2(n1724), .ZN(n1427)
         );
  OAI22_X1 U2697 ( .A1(n2217), .A2(n1723), .B1(n2231), .B2(n1722), .ZN(n1425)
         );
  OAI22_X1 U2698 ( .A1(n2069), .A2(n1728), .B1(n1727), .B2(n2141), .ZN(n1430)
         );
  OAI22_X1 U2699 ( .A1(n2217), .A2(n1729), .B1(n2231), .B2(n1728), .ZN(n1431)
         );
  OAI22_X1 U2700 ( .A1(n2216), .A2(n1722), .B1(n1721), .B2(n2231), .ZN(n1424)
         );
  OAI22_X1 U2701 ( .A1(n2217), .A2(n1719), .B1(n2231), .B2(n1718), .ZN(n1421)
         );
  OAI22_X1 U2702 ( .A1(n2217), .A2(n1724), .B1(n1723), .B2(n2231), .ZN(n1426)
         );
  INV_X1 U2703 ( .A(n325), .ZN(product[47]) );
  AOI21_X1 U2704 ( .B1(n423), .B2(n356), .A(n359), .ZN(n355) );
  NAND2_X1 U2705 ( .A1(n422), .A2(n356), .ZN(n354) );
  OAI22_X1 U2706 ( .A1(n1929), .A2(n1563), .B1(n2223), .B2(n1562), .ZN(n1271)
         );
  OAI22_X1 U2707 ( .A1(n1987), .A2(n1566), .B1(n1565), .B2(n2223), .ZN(n1274)
         );
  OAI22_X1 U2708 ( .A1(n1929), .A2(n1561), .B1(n2222), .B2(n1560), .ZN(n1269)
         );
  OAI22_X1 U2709 ( .A1(n1929), .A2(n1567), .B1(n2222), .B2(n1566), .ZN(n1275)
         );
  OAI22_X1 U2710 ( .A1(n1929), .A2(n1564), .B1(n1563), .B2(n2223), .ZN(n1272)
         );
  OAI22_X1 U2711 ( .A1(n1929), .A2(n1560), .B1(n1559), .B2(n2222), .ZN(n1268)
         );
  OAI22_X1 U2712 ( .A1(n1929), .A2(n1559), .B1(n2222), .B2(n1558), .ZN(n1267)
         );
  OAI22_X1 U2713 ( .A1(n1581), .A2(n2223), .B1(n1929), .B2(n2248), .ZN(n1185)
         );
  OAI22_X1 U2714 ( .A1(n1987), .A2(n1565), .B1(n2222), .B2(n1564), .ZN(n1273)
         );
  INV_X1 U2715 ( .A(n706), .ZN(n707) );
  OAI22_X1 U2716 ( .A1(n1987), .A2(n1562), .B1(n1561), .B2(n2223), .ZN(n1270)
         );
  OAI22_X1 U2717 ( .A1(n2040), .A2(n1568), .B1(n1567), .B2(n2222), .ZN(n1276)
         );
  OAI22_X1 U2718 ( .A1(n1929), .A2(n1558), .B1(n1557), .B2(n2223), .ZN(n706)
         );
  XNOR2_X1 U2719 ( .A(n342), .B(n302), .ZN(product[44]) );
  OAI21_X1 U2720 ( .B1(n2007), .B2(n326), .A(n327), .ZN(n325) );
  OAI21_X1 U2721 ( .B1(n2203), .B2(n411), .A(n412), .ZN(n410) );
  OAI21_X1 U2722 ( .B1(n301), .B2(n431), .A(n432), .ZN(n430) );
  OAI21_X1 U2723 ( .B1(n2203), .B2(n354), .A(n355), .ZN(n353) );
  OAI21_X1 U2724 ( .B1(n301), .B2(n420), .A(n421), .ZN(n419) );
  OAI21_X1 U2725 ( .B1(n2202), .B2(n398), .A(n399), .ZN(n397) );
  OAI21_X1 U2726 ( .B1(n301), .B2(n438), .A(n439), .ZN(n437) );
  OAI21_X1 U2727 ( .B1(n301), .B2(n2170), .A(n344), .ZN(n342) );
  OAI21_X1 U2728 ( .B1(n2203), .B2(n389), .A(n390), .ZN(n388) );
  OAI21_X1 U2729 ( .B1(n2203), .B2(n371), .A(n372), .ZN(n370) );
  OAI21_X1 U2730 ( .B1(n2202), .B2(n380), .A(n381), .ZN(n379) );
  OAI22_X1 U2731 ( .A1(n2193), .A2(n1691), .B1(n1690), .B2(n2002), .ZN(n1394)
         );
  OAI22_X1 U2732 ( .A1(n2193), .A2(n1686), .B1(n2228), .B2(n1685), .ZN(n1389)
         );
  OAI22_X1 U2733 ( .A1(n2193), .A2(n1689), .B1(n1688), .B2(n2002), .ZN(n1392)
         );
  OAI22_X1 U2734 ( .A1(n2193), .A2(n1690), .B1(n2002), .B2(n1689), .ZN(n1393)
         );
  OAI22_X1 U2735 ( .A1(n2193), .A2(n1687), .B1(n1686), .B2(n2002), .ZN(n1390)
         );
  OAI22_X1 U2736 ( .A1(n2193), .A2(n1692), .B1(n2002), .B2(n1691), .ZN(n1395)
         );
  OAI22_X1 U2737 ( .A1(n2193), .A2(n1685), .B1(n1684), .B2(n2002), .ZN(n1388)
         );
  OAI22_X1 U2738 ( .A1(n2193), .A2(n1688), .B1(n2228), .B2(n1687), .ZN(n1391)
         );
  INV_X1 U2739 ( .A(n836), .ZN(n837) );
  OAI22_X1 U2740 ( .A1(n2193), .A2(n1684), .B1(n2228), .B2(n1683), .ZN(n1387)
         );
  OAI22_X1 U2741 ( .A1(n2214), .A2(n1693), .B1(n1692), .B2(n2228), .ZN(n1396)
         );
  OAI22_X1 U2742 ( .A1(n1706), .A2(n2002), .B1(n2096), .B2(n2269), .ZN(n1190)
         );
  INV_X2 U2743 ( .A(n2135), .ZN(n2210) );
  INV_X2 U2744 ( .A(n2273), .ZN(n2271) );
  INV_X1 U2745 ( .A(n2177), .ZN(n2212) );
  INV_X1 U2746 ( .A(n2128), .ZN(n2223) );
  INV_X1 U2747 ( .A(n2129), .ZN(n2233) );
  INV_X1 U2748 ( .A(n1968), .ZN(n2239) );
  INV_X1 U2749 ( .A(n2248), .ZN(n2245) );
  INV_X1 U2750 ( .A(n2248), .ZN(n2247) );
  INV_X1 U2751 ( .A(n2255), .ZN(n2252) );
  INV_X1 U2752 ( .A(n2259), .ZN(n2258) );
  INV_X1 U2753 ( .A(n2264), .ZN(n2263) );
  INV_X1 U2754 ( .A(n2269), .ZN(n2268) );
  INV_X1 U2755 ( .A(n2273), .ZN(n2270) );
  INV_X1 U2756 ( .A(n2273), .ZN(n2272) );
  INV_X1 U2757 ( .A(n2277), .ZN(n2276) );
  INV_X1 U2758 ( .A(n1936), .ZN(n2280) );
endmodule


module iir_filter_DW_mult_tc_0 ( a, b, product );
  input [23:0] a;
  input [23:0] b;
  output [47:0] product;
  wire   n251, n285, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n323, n325, n326, n327, n332, n333, n334, n335, n336, n337, n339,
         n341, n342, n343, n344, n345, n346, n347, n348, n350, n352, n353,
         n354, n355, n356, n359, n360, n361, n362, n363, n364, n365, n367,
         n369, n370, n371, n372, n376, n378, n379, n380, n381, n382, n383,
         n384, n387, n388, n389, n390, n394, n396, n397, n398, n399, n400,
         n401, n402, n405, n407, n409, n410, n411, n412, n416, n418, n419,
         n420, n421, n422, n423, n426, n427, n428, n429, n430, n431, n432,
         n434, n435, n436, n437, n438, n439, n445, n450, n451, n452, n453,
         n454, n455, n456, n457, n459, n461, n462, n463, n464, n465, n466,
         n467, n468, n472, n474, n475, n476, n477, n478, n479, n480, n481,
         n483, n486, n487, n488, n489, n490, n492, n495, n496, n497, n498,
         n499, n501, n502, n503, n504, n505, n506, n508, n511, n512, n513,
         n514, n515, n516, n517, n519, n520, n521, n522, n523, n524, n525,
         n526, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n550, n551, n552, n553,
         n554, n555, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n581, n582, n583, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n609, n610, n611, n620, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n643, n644, n645, n646,
         n657, n661, n662, n666, n667, n668, n671, n674, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1806, n1808, n1809, n1810, n1812, n1813,
         n1817, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324;

  FA_X1 U546 ( .A(n1195), .B(n682), .CI(n1218), .CO(n678), .S(n679) );
  FA_X1 U547 ( .A(n683), .B(n1196), .CI(n686), .CO(n680), .S(n681) );
  FA_X1 U549 ( .A(n690), .B(n1242), .CI(n687), .CO(n684), .S(n685) );
  FA_X1 U550 ( .A(n1219), .B(n692), .CI(n1197), .CO(n686), .S(n687) );
  FA_X1 U551 ( .A(n691), .B(n698), .CI(n696), .CO(n688), .S(n689) );
  FA_X1 U552 ( .A(n1198), .B(n1220), .CI(n693), .CO(n690), .S(n691) );
  FA_X1 U554 ( .A(n702), .B(n699), .CI(n697), .CO(n694), .S(n695) );
  FA_X1 U555 ( .A(n1266), .B(n1243), .CI(n704), .CO(n696), .S(n697) );
  FA_X1 U556 ( .A(n1221), .B(n1199), .CI(n706), .CO(n698), .S(n699) );
  FA_X1 U557 ( .A(n710), .B(n712), .CI(n703), .CO(n700), .S(n701) );
  FA_X1 U558 ( .A(n714), .B(n1244), .CI(n705), .CO(n702), .S(n703) );
  FA_X1 U559 ( .A(n1222), .B(n1200), .CI(n707), .CO(n704), .S(n705) );
  FA_X1 U561 ( .A(n718), .B(n713), .CI(n711), .CO(n708), .S(n709) );
  FA_X1 U562 ( .A(n715), .B(n722), .CI(n720), .CO(n710), .S(n711) );
  FA_X1 U563 ( .A(n1245), .B(n1223), .CI(n1290), .CO(n712), .S(n713) );
  FA_X1 U564 ( .A(n1267), .B(n1201), .CI(n724), .CO(n714), .S(n715) );
  FA_X1 U565 ( .A(n728), .B(n721), .CI(n719), .CO(n716), .S(n717) );
  FA_X1 U566 ( .A(n723), .B(n732), .CI(n730), .CO(n718), .S(n719) );
  FA_X1 U567 ( .A(n1202), .B(n1246), .CI(n734), .CO(n720), .S(n721) );
  FA_X1 U568 ( .A(n1268), .B(n1224), .CI(n725), .CO(n722), .S(n723) );
  FA_X1 U570 ( .A(n738), .B(n731), .CI(n729), .CO(n726), .S(n727) );
  FA_X1 U571 ( .A(n735), .B(n733), .CI(n740), .CO(n728), .S(n729) );
  FA_X1 U572 ( .A(n744), .B(n1314), .CI(n742), .CO(n730), .S(n731) );
  FA_X1 U573 ( .A(n1225), .B(n1291), .CI(n1269), .CO(n732), .S(n733) );
  FA_X1 U574 ( .A(n746), .B(n1203), .CI(n1247), .CO(n734), .S(n735) );
  FA_X1 U575 ( .A(n750), .B(n741), .CI(n739), .CO(n736), .S(n737) );
  FA_X1 U576 ( .A(n754), .B(n745), .CI(n752), .CO(n738), .S(n739) );
  FA_X1 U577 ( .A(n756), .B(n758), .CI(n743), .CO(n740), .S(n741) );
  FA_X1 U578 ( .A(n1226), .B(n1204), .CI(n1270), .CO(n742), .S(n743) );
  FA_X1 U579 ( .A(n1292), .B(n1248), .CI(n747), .CO(n744), .S(n745) );
  FA_X1 U581 ( .A(n762), .B(n753), .CI(n751), .CO(n748), .S(n749) );
  FA_X1 U582 ( .A(n755), .B(n766), .CI(n764), .CO(n750), .S(n751) );
  FA_X1 U583 ( .A(n757), .B(n768), .CI(n759), .CO(n752), .S(n753) );
  FA_X1 U584 ( .A(n1338), .B(n1271), .CI(n770), .CO(n754), .S(n755) );
  FA_X1 U585 ( .A(n1249), .B(n1293), .CI(n1315), .CO(n756), .S(n757) );
  FA_X1 U586 ( .A(n772), .B(n1205), .CI(n1227), .CO(n758), .S(n759) );
  FA_X1 U587 ( .A(n776), .B(n765), .CI(n763), .CO(n760), .S(n761) );
  FA_X1 U588 ( .A(n767), .B(n780), .CI(n778), .CO(n762), .S(n763) );
  FA_X1 U589 ( .A(n771), .B(n769), .CI(n782), .CO(n764), .S(n765) );
  FA_X1 U590 ( .A(n786), .B(n1228), .CI(n784), .CO(n766), .S(n767) );
  FA_X1 U591 ( .A(n1294), .B(n1206), .CI(n1272), .CO(n768), .S(n769) );
  FA_X1 U592 ( .A(n1316), .B(n1250), .CI(n773), .CO(n770), .S(n771) );
  FA_X1 U594 ( .A(n790), .B(n779), .CI(n777), .CO(n774), .S(n775) );
  FA_X1 U595 ( .A(n781), .B(n794), .CI(n792), .CO(n776), .S(n777) );
  FA_X1 U596 ( .A(n796), .B(n787), .CI(n783), .CO(n778), .S(n779) );
  FA_X1 U597 ( .A(n798), .B(n800), .CI(n785), .CO(n780), .S(n781) );
  FA_X1 U598 ( .A(n1339), .B(n1229), .CI(n1362), .CO(n782), .S(n783) );
  FA_X1 U599 ( .A(n1273), .B(n1317), .CI(n1295), .CO(n784), .S(n785) );
  FA_X1 U600 ( .A(n1251), .B(n1207), .CI(n2012), .CO(n786), .S(n787) );
  FA_X1 U601 ( .A(n806), .B(n793), .CI(n791), .CO(n788), .S(n789) );
  FA_X1 U602 ( .A(n795), .B(n810), .CI(n808), .CO(n790), .S(n791) );
  FA_X1 U603 ( .A(n797), .B(n801), .CI(n812), .CO(n792), .S(n793) );
  FA_X1 U604 ( .A(n814), .B(n816), .CI(n799), .CO(n794), .S(n795) );
  FA_X1 U606 ( .A(n1208), .B(n1318), .CI(n1230), .CO(n798), .S(n799) );
  FA_X1 U607 ( .A(n1340), .B(n1252), .CI(n803), .CO(n800), .S(n801) );
  FA_X1 U609 ( .A(n822), .B(n809), .CI(n807), .CO(n804), .S(n805) );
  FA_X1 U610 ( .A(n811), .B(n826), .CI(n824), .CO(n806), .S(n807) );
  FA_X1 U611 ( .A(n828), .B(n819), .CI(n813), .CO(n808), .S(n809) );
  FA_X1 U612 ( .A(n815), .B(n832), .CI(n817), .CO(n810), .S(n811) );
  FA_X1 U613 ( .A(n834), .B(n1386), .CI(n830), .CO(n812), .S(n813) );
  FA_X1 U614 ( .A(n1319), .B(n1253), .CI(n1341), .CO(n814), .S(n815) );
  FA_X1 U615 ( .A(n1231), .B(n1297), .CI(n1275), .CO(n816), .S(n817) );
  FA_X1 U618 ( .A(n827), .B(n844), .CI(n842), .CO(n822), .S(n823) );
  FA_X1 U619 ( .A(n846), .B(n848), .CI(n829), .CO(n824), .S(n825) );
  FA_X1 U620 ( .A(n835), .B(n831), .CI(n833), .CO(n826), .S(n827) );
  FA_X1 U621 ( .A(n850), .B(n854), .CI(n852), .CO(n828), .S(n829) );
  FA_X1 U622 ( .A(n1254), .B(n1320), .CI(n1298), .CO(n830), .S(n831) );
  FA_X1 U623 ( .A(n1232), .B(n1364), .CI(n1342), .CO(n832), .S(n833) );
  FA_X1 U624 ( .A(n1276), .B(n1210), .CI(n837), .CO(n834), .S(n835) );
  FA_X1 U626 ( .A(n858), .B(n843), .CI(n841), .CO(n838), .S(n839) );
  FA_X1 U627 ( .A(n845), .B(n847), .CI(n860), .CO(n840), .S(n841) );
  FA_X1 U628 ( .A(n864), .B(n849), .CI(n862), .CO(n842), .S(n843) );
  FA_X1 U629 ( .A(n855), .B(n853), .CI(n866), .CO(n844), .S(n845) );
  FA_X1 U630 ( .A(n868), .B(n870), .CI(n851), .CO(n846), .S(n847) );
  FA_X1 U631 ( .A(n1410), .B(n1365), .CI(n872), .CO(n848), .S(n849) );
  FA_X1 U632 ( .A(n1343), .B(n1277), .CI(n1299), .CO(n850), .S(n851) );
  FA_X1 U633 ( .A(n1255), .B(n1321), .CI(n1983), .CO(n852), .S(n853) );
  FA_X1 U634 ( .A(n1387), .B(n1211), .CI(n1233), .CO(n854), .S(n855) );
  FA_X1 U637 ( .A(n867), .B(n884), .CI(n865), .CO(n860), .S(n861) );
  FA_X1 U638 ( .A(n873), .B(n888), .CI(n886), .CO(n862), .S(n863) );
  FA_X1 U639 ( .A(n869), .B(n890), .CI(n871), .CO(n864), .S(n865) );
  FA_X1 U640 ( .A(n894), .B(n1300), .CI(n892), .CO(n866), .S(n867) );
  FA_X1 U641 ( .A(n1234), .B(n1322), .CI(n1256), .CO(n868), .S(n869) );
  FA_X1 U642 ( .A(n1344), .B(n1212), .CI(n1366), .CO(n870), .S(n871) );
  FA_X1 U643 ( .A(n1388), .B(n1278), .CI(n875), .CO(n872), .S(n873) );
  FA_X1 U645 ( .A(n898), .B(n881), .CI(n879), .CO(n876), .S(n877) );
  FA_X1 U646 ( .A(n883), .B(n885), .CI(n900), .CO(n878), .S(n879) );
  FA_X1 U649 ( .A(n895), .B(n908), .CI(n891), .CO(n884), .S(n885) );
  FA_X1 U650 ( .A(n914), .B(n910), .CI(n912), .CO(n886), .S(n887) );
  FA_X1 U651 ( .A(n1367), .B(n1389), .CI(n1434), .CO(n888), .S(n889) );
  FA_X1 U652 ( .A(n1257), .B(n1301), .CI(n1345), .CO(n890), .S(n891) );
  FA_X1 U653 ( .A(n2042), .B(n1323), .CI(n1279), .CO(n892), .S(n893) );
  FA_X1 U654 ( .A(n1411), .B(n1213), .CI(n1235), .CO(n894), .S(n895) );
  FA_X1 U655 ( .A(n920), .B(n901), .CI(n899), .CO(n896), .S(n897) );
  FA_X1 U656 ( .A(n903), .B(n924), .CI(n922), .CO(n898), .S(n899) );
  FA_X1 U658 ( .A(n909), .B(n930), .CI(n928), .CO(n902), .S(n903) );
  FA_X1 U659 ( .A(n915), .B(n911), .CI(n913), .CO(n904), .S(n905) );
  FA_X1 U660 ( .A(n932), .B(n936), .CI(n934), .CO(n906), .S(n907) );
  FA_X1 U661 ( .A(n1368), .B(n1390), .CI(n938), .CO(n908), .S(n909) );
  FA_X1 U662 ( .A(n1346), .B(n1280), .CI(n1324), .CO(n910), .S(n911) );
  FA_X1 U663 ( .A(n1412), .B(n1236), .CI(n1258), .CO(n912), .S(n913) );
  FA_X1 U664 ( .A(n917), .B(n1214), .CI(n1302), .CO(n914), .S(n915) );
  FA_X1 U666 ( .A(n942), .B(n923), .CI(n921), .CO(n918), .S(n919) );
  FA_X1 U667 ( .A(n925), .B(n927), .CI(n944), .CO(n920), .S(n921) );
  FA_X1 U668 ( .A(n929), .B(n948), .CI(n946), .CO(n922), .S(n923) );
  FA_X1 U669 ( .A(n950), .B(n935), .CI(n931), .CO(n924), .S(n925) );
  FA_X1 U671 ( .A(n954), .B(n958), .CI(n956), .CO(n928), .S(n929) );
  FA_X1 U672 ( .A(n1458), .B(n960), .CI(n939), .CO(n930), .S(n931) );
  FA_X1 U674 ( .A(n1281), .B(n1369), .CI(n1391), .CO(n934), .S(n935) );
  FA_X1 U675 ( .A(n1259), .B(n1347), .CI(n1303), .CO(n936), .S(n937) );
  FA_X1 U680 ( .A(n951), .B(n970), .CI(n968), .CO(n944), .S(n945) );
  FA_X1 U682 ( .A(n955), .B(n974), .CI(n957), .CO(n948), .S(n949) );
  FA_X1 U683 ( .A(n976), .B(n980), .CI(n978), .CO(n950), .S(n951) );
  FA_X1 U685 ( .A(n1282), .B(n1304), .CI(n1414), .CO(n954), .S(n955) );
  FA_X1 U686 ( .A(n1370), .B(n1459), .CI(n1436), .CO(n956), .S(n957) );
  FA_X1 U687 ( .A(n1260), .B(n1348), .CI(n1182), .CO(n958), .S(n959) );
  HA_X1 U688 ( .A(n1238), .B(n1216), .CO(n960), .S(n961) );
  FA_X1 U689 ( .A(n984), .B(n967), .CI(n965), .CO(n962), .S(n963) );
  FA_X1 U690 ( .A(n969), .B(n971), .CI(n986), .CO(n964), .S(n965) );
  FA_X1 U691 ( .A(n973), .B(n990), .CI(n988), .CO(n966), .S(n967) );
  FA_X1 U693 ( .A(n977), .B(n998), .CI(n979), .CO(n970), .S(n971) );
  FA_X1 U696 ( .A(n1327), .B(n1437), .CI(n1305), .CO(n976), .S(n977) );
  FA_X1 U697 ( .A(n1460), .B(n1371), .CI(n1283), .CO(n978), .S(n979) );
  FA_X1 U698 ( .A(n1349), .B(n1239), .CI(n1261), .CO(n980), .S(n981) );
  FA_X1 U699 ( .A(n1004), .B(n987), .CI(n985), .CO(n982), .S(n983) );
  FA_X1 U700 ( .A(n989), .B(n991), .CI(n1006), .CO(n984), .S(n985) );
  FA_X1 U701 ( .A(n993), .B(n1010), .CI(n1008), .CO(n986), .S(n987) );
  FA_X1 U702 ( .A(n999), .B(n997), .CI(n1012), .CO(n988), .S(n989) );
  FA_X1 U703 ( .A(n1014), .B(n1016), .CI(n995), .CO(n990), .S(n991) );
  FA_X1 U704 ( .A(n1001), .B(n1394), .CI(n1018), .CO(n992), .S(n993) );
  FA_X1 U705 ( .A(n1306), .B(n1416), .CI(n1328), .CO(n994), .S(n995) );
  FA_X1 U707 ( .A(n1461), .B(n1350), .CI(n1183), .CO(n998), .S(n999) );
  FA_X1 U709 ( .A(n1022), .B(n1007), .CI(n1005), .CO(n1002), .S(n1003) );
  FA_X1 U710 ( .A(n1009), .B(n1011), .CI(n1024), .CO(n1004), .S(n1005) );
  FA_X1 U711 ( .A(n1013), .B(n1028), .CI(n1026), .CO(n1006), .S(n1007) );
  FA_X1 U712 ( .A(n1019), .B(n1015), .CI(n1017), .CO(n1008), .S(n1009) );
  FA_X1 U713 ( .A(n1241), .B(n1034), .CI(n1030), .CO(n1010), .S(n1011) );
  FA_X1 U714 ( .A(n1036), .B(n1439), .CI(n1032), .CO(n1012), .S(n1013) );
  FA_X1 U715 ( .A(n1395), .B(n1462), .CI(n1417), .CO(n1014), .S(n1015) );
  FA_X1 U716 ( .A(n1307), .B(n1329), .CI(n1373), .CO(n1016), .S(n1017) );
  FA_X1 U717 ( .A(n1351), .B(n1285), .CI(n1263), .CO(n1018), .S(n1019) );
  FA_X1 U718 ( .A(n1023), .B(n1025), .CI(n1040), .CO(n1020), .S(n1021) );
  FA_X1 U720 ( .A(n1046), .B(n1035), .CI(n1029), .CO(n1024), .S(n1025) );
  FA_X1 U721 ( .A(n1033), .B(n1048), .CI(n1031), .CO(n1026), .S(n1027) );
  FA_X1 U722 ( .A(n1052), .B(n1037), .CI(n1050), .CO(n1028), .S(n1029) );
  FA_X1 U723 ( .A(n1352), .B(n1440), .CI(n1418), .CO(n1030), .S(n1031) );
  FA_X1 U724 ( .A(n1463), .B(n1396), .CI(n1330), .CO(n1032), .S(n1033) );
  FA_X1 U725 ( .A(n1184), .B(n1308), .CI(n1374), .CO(n1034), .S(n1035) );
  HA_X1 U726 ( .A(n1264), .B(n1286), .CO(n1036), .S(n1037) );
  FA_X1 U728 ( .A(n1058), .B(n1047), .CI(n1045), .CO(n1040), .S(n1041) );
  FA_X1 U730 ( .A(n1049), .B(n1265), .CI(n1051), .CO(n1044), .S(n1045) );
  FA_X1 U731 ( .A(n1064), .B(n1068), .CI(n1066), .CO(n1046), .S(n1047) );
  FA_X1 U732 ( .A(n1397), .B(n1441), .CI(n1419), .CO(n1048), .S(n1049) );
  FA_X1 U733 ( .A(n1331), .B(n1353), .CI(n1375), .CO(n1050), .S(n1051) );
  FA_X1 U735 ( .A(n1072), .B(n1059), .CI(n1057), .CO(n1054), .S(n1055) );
  FA_X1 U736 ( .A(n1074), .B(n1063), .CI(n1061), .CO(n1056), .S(n1057) );
  FA_X1 U737 ( .A(n1067), .B(n1065), .CI(n1076), .CO(n1058), .S(n1059) );
  FA_X1 U738 ( .A(n1080), .B(n1082), .CI(n1078), .CO(n1060), .S(n1061) );
  FA_X1 U739 ( .A(n1398), .B(n1420), .CI(n1069), .CO(n1062), .S(n1063) );
  FA_X1 U740 ( .A(n1442), .B(n1354), .CI(n1332), .CO(n1064), .S(n1065) );
  FA_X1 U741 ( .A(n1465), .B(n1376), .CI(n1185), .CO(n1066), .S(n1067) );
  HA_X1 U742 ( .A(n1288), .B(n1310), .CO(n1068), .S(n1069) );
  FA_X1 U743 ( .A(n1086), .B(n1075), .CI(n1073), .CO(n1070), .S(n1071) );
  FA_X1 U744 ( .A(n1088), .B(n1090), .CI(n1077), .CO(n1072), .S(n1073) );
  FA_X1 U745 ( .A(n1083), .B(n1081), .CI(n1079), .CO(n1074), .S(n1075) );
  FA_X1 U746 ( .A(n1092), .B(n1094), .CI(n1289), .CO(n1076), .S(n1077) );
  FA_X1 U747 ( .A(n1399), .B(n1421), .CI(n1096), .CO(n1078), .S(n1079) );
  FA_X1 U748 ( .A(n1377), .B(n1443), .CI(n1355), .CO(n1080), .S(n1081) );
  FA_X1 U749 ( .A(n1311), .B(n1466), .CI(n1333), .CO(n1082), .S(n1083) );
  FA_X1 U750 ( .A(n1100), .B(n1089), .CI(n1087), .CO(n1084), .S(n1085) );
  FA_X1 U751 ( .A(n1102), .B(n1104), .CI(n1091), .CO(n1086), .S(n1087) );
  FA_X1 U752 ( .A(n1093), .B(n1106), .CI(n1095), .CO(n1088), .S(n1089) );
  FA_X1 U753 ( .A(n1097), .B(n1422), .CI(n1108), .CO(n1090), .S(n1091) );
  FA_X1 U754 ( .A(n1356), .B(n1378), .CI(n1444), .CO(n1092), .S(n1093) );
  FA_X1 U755 ( .A(n1186), .B(n1400), .CI(n1467), .CO(n1094), .S(n1095) );
  HA_X1 U756 ( .A(n1334), .B(n1312), .CO(n1096), .S(n1097) );
  FA_X1 U757 ( .A(n1103), .B(n1112), .CI(n1101), .CO(n1098), .S(n1099) );
  FA_X1 U758 ( .A(n1114), .B(n1109), .CI(n1105), .CO(n1100), .S(n1101) );
  FA_X1 U759 ( .A(n1313), .B(n1116), .CI(n1107), .CO(n1102), .S(n1103) );
  FA_X1 U760 ( .A(n1120), .B(n1423), .CI(n1118), .CO(n1104), .S(n1105) );
  FA_X1 U761 ( .A(n1379), .B(n1445), .CI(n1401), .CO(n1106), .S(n1107) );
  FA_X1 U762 ( .A(n1335), .B(n1468), .CI(n1357), .CO(n1108), .S(n1109) );
  FA_X1 U763 ( .A(n1124), .B(n1115), .CI(n1113), .CO(n1110), .S(n1111) );
  FA_X1 U764 ( .A(n1119), .B(n1117), .CI(n1126), .CO(n1112), .S(n1113) );
  FA_X1 U765 ( .A(n1130), .B(n1121), .CI(n1128), .CO(n1114), .S(n1115) );
  FA_X1 U766 ( .A(n1380), .B(n1446), .CI(n1424), .CO(n1116), .S(n1117) );
  FA_X1 U767 ( .A(n1469), .B(n1402), .CI(n1187), .CO(n1118), .S(n1119) );
  HA_X1 U768 ( .A(n1336), .B(n1358), .CO(n1120), .S(n1121) );
  FA_X1 U769 ( .A(n1127), .B(n1134), .CI(n1125), .CO(n1122), .S(n1123) );
  FA_X1 U770 ( .A(n1131), .B(n1129), .CI(n1136), .CO(n1124), .S(n1125) );
  FA_X1 U771 ( .A(n1138), .B(n1140), .CI(n1337), .CO(n1126), .S(n1127) );
  FA_X1 U772 ( .A(n1403), .B(n1447), .CI(n1425), .CO(n1128), .S(n1129) );
  FA_X1 U773 ( .A(n1359), .B(n1470), .CI(n1381), .CO(n1130), .S(n1131) );
  FA_X1 U774 ( .A(n1144), .B(n1137), .CI(n1135), .CO(n1132), .S(n1133) );
  FA_X1 U775 ( .A(n1146), .B(n1148), .CI(n1139), .CO(n1134), .S(n1135) );
  FA_X1 U776 ( .A(n1404), .B(n1448), .CI(n1141), .CO(n1136), .S(n1137) );
  FA_X1 U777 ( .A(n1471), .B(n1188), .CI(n1426), .CO(n1138), .S(n1139) );
  HA_X1 U778 ( .A(n1360), .B(n1382), .CO(n1140), .S(n1141) );
  FA_X1 U779 ( .A(n1152), .B(n1147), .CI(n1145), .CO(n1142), .S(n1143) );
  FA_X1 U780 ( .A(n1361), .B(n1154), .CI(n1149), .CO(n1144), .S(n1145) );
  FA_X1 U781 ( .A(n1427), .B(n1449), .CI(n1156), .CO(n1146), .S(n1147) );
  FA_X1 U782 ( .A(n1383), .B(n1472), .CI(n1405), .CO(n1148), .S(n1149) );
  FA_X1 U783 ( .A(n1160), .B(n1155), .CI(n1153), .CO(n1150), .S(n1151) );
  FA_X1 U784 ( .A(n1157), .B(n1473), .CI(n1162), .CO(n1152), .S(n1153) );
  FA_X1 U785 ( .A(n1450), .B(n1428), .CI(n1189), .CO(n1154), .S(n1155) );
  HA_X1 U786 ( .A(n1384), .B(n1406), .CO(n1156), .S(n1157) );
  FA_X1 U787 ( .A(n1163), .B(n1385), .CI(n1164), .CO(n1158), .S(n1159) );
  FA_X1 U788 ( .A(n1168), .B(n1429), .CI(n1166), .CO(n1160), .S(n1161) );
  FA_X1 U789 ( .A(n1451), .B(n1474), .CI(n1407), .CO(n1162), .S(n1163) );
  FA_X1 U790 ( .A(n1172), .B(n1169), .CI(n1167), .CO(n1164), .S(n1165) );
  FA_X1 U791 ( .A(n1452), .B(n1475), .CI(n1190), .CO(n1166), .S(n1167) );
  HA_X1 U792 ( .A(n1408), .B(n1430), .CO(n1168), .S(n1169) );
  FA_X1 U793 ( .A(n1409), .B(n1176), .CI(n1173), .CO(n1170), .S(n1171) );
  FA_X1 U794 ( .A(n1476), .B(n1453), .CI(n1431), .CO(n1172), .S(n1173) );
  FA_X1 U795 ( .A(n1191), .B(n1454), .CI(n1177), .CO(n1174), .S(n1175) );
  HA_X1 U796 ( .A(n1432), .B(n1477), .CO(n1176), .S(n1177) );
  FA_X1 U797 ( .A(n1455), .B(n1478), .CI(n1180), .CO(n1178), .S(n1179) );
  HA_X1 U798 ( .A(n1456), .B(n1479), .CO(n1180), .S(n1181) );
  CLKBUF_X1 U1448 ( .A(n919), .Z(n1929) );
  XOR2_X1 U1449 ( .A(n1262), .B(n1240), .Z(n1001) );
  INV_X1 U1450 ( .A(n1930), .ZN(n1000) );
  NAND2_X1 U1451 ( .A1(n1240), .A2(n1262), .ZN(n1930) );
  INV_X1 U1452 ( .A(n2300), .ZN(n1931) );
  INV_X2 U1453 ( .A(n2131), .ZN(n2226) );
  OR2_X1 U1454 ( .A1(n1021), .A2(n1038), .ZN(n1932) );
  BUF_X2 U1455 ( .A(n251), .Z(n2257) );
  AND2_X2 U1456 ( .A1(n1817), .A2(n2257), .ZN(n2133) );
  INV_X1 U1457 ( .A(n2143), .ZN(n1933) );
  BUF_X1 U1458 ( .A(n2085), .Z(n2149) );
  INV_X1 U1459 ( .A(a[15]), .ZN(n1934) );
  XNOR2_X1 U1460 ( .A(n544), .B(n1935), .ZN(product[24]) );
  AND2_X1 U1461 ( .A1(n2195), .A2(n2005), .ZN(n1935) );
  INV_X1 U1462 ( .A(a[9]), .ZN(n1936) );
  XNOR2_X1 U1463 ( .A(n1937), .B(n818), .ZN(n797) );
  XNOR2_X1 U1464 ( .A(n1274), .B(n1296), .ZN(n1937) );
  INV_X1 U1465 ( .A(n2273), .ZN(n2269) );
  INV_X2 U1466 ( .A(n2264), .ZN(n1977) );
  XNOR2_X1 U1467 ( .A(a[0]), .B(n2311), .ZN(n1817) );
  INV_X1 U1468 ( .A(a[23]), .ZN(n1938) );
  INV_X2 U1469 ( .A(n1938), .ZN(n1939) );
  INV_X2 U1470 ( .A(n2018), .ZN(n2243) );
  INV_X2 U1471 ( .A(n2131), .ZN(n2160) );
  BUF_X1 U1472 ( .A(a[16]), .Z(n2024) );
  CLKBUF_X1 U1473 ( .A(n2051), .Z(n2151) );
  CLKBUF_X3 U1474 ( .A(n2051), .Z(n2152) );
  CLKBUF_X3 U1475 ( .A(n2051), .Z(n2153) );
  INV_X1 U1476 ( .A(n2134), .ZN(n2229) );
  XNOR2_X1 U1477 ( .A(n1940), .B(n975), .ZN(n969) );
  XNOR2_X1 U1478 ( .A(n981), .B(n992), .ZN(n1940) );
  INV_X2 U1479 ( .A(n2295), .ZN(n2292) );
  XOR2_X1 U1480 ( .A(n1393), .B(n1415), .Z(n1941) );
  XOR2_X1 U1481 ( .A(n1941), .B(n1000), .Z(n975) );
  NAND2_X1 U1482 ( .A1(n1393), .A2(n1415), .ZN(n1942) );
  NAND2_X1 U1483 ( .A1(n1393), .A2(n1000), .ZN(n1943) );
  NAND2_X1 U1484 ( .A1(n1415), .A2(n1000), .ZN(n1944) );
  NAND3_X1 U1485 ( .A1(n1942), .A2(n1943), .A3(n1944), .ZN(n974) );
  NAND2_X1 U1486 ( .A1(n981), .A2(n992), .ZN(n1945) );
  NAND2_X1 U1487 ( .A1(n981), .A2(n975), .ZN(n1946) );
  NAND2_X1 U1488 ( .A1(n992), .A2(n975), .ZN(n1947) );
  NAND3_X1 U1489 ( .A1(n1945), .A2(n1946), .A3(n1947), .ZN(n968) );
  BUF_X2 U1490 ( .A(n2085), .Z(n2147) );
  NOR2_X1 U1491 ( .A1(n1003), .A2(n1020), .ZN(n1948) );
  CLKBUF_X2 U1492 ( .A(a[19]), .Z(n1981) );
  BUF_X1 U1493 ( .A(n2132), .Z(n1992) );
  BUF_X1 U1494 ( .A(a[18]), .Z(n1949) );
  XOR2_X1 U1495 ( .A(n840), .B(n825), .Z(n1950) );
  XOR2_X1 U1496 ( .A(n823), .B(n1950), .Z(n821) );
  NAND2_X1 U1497 ( .A1(n823), .A2(n840), .ZN(n1951) );
  NAND2_X1 U1498 ( .A1(n823), .A2(n825), .ZN(n1952) );
  NAND2_X1 U1499 ( .A1(n840), .A2(n825), .ZN(n1953) );
  NAND3_X1 U1500 ( .A1(n1951), .A2(n1952), .A3(n1953), .ZN(n820) );
  BUF_X1 U1501 ( .A(n2108), .Z(n2107) );
  BUF_X1 U1502 ( .A(n553), .Z(n2055) );
  CLKBUF_X3 U1503 ( .A(a[11]), .Z(n1954) );
  INV_X1 U1504 ( .A(n2134), .ZN(n1956) );
  INV_X1 U1505 ( .A(n2134), .ZN(n1955) );
  INV_X1 U1506 ( .A(n2069), .ZN(n2191) );
  BUF_X1 U1507 ( .A(n2085), .Z(n2148) );
  BUF_X1 U1508 ( .A(n285), .Z(n2208) );
  AND2_X1 U1509 ( .A1(n1193), .A2(n1481), .ZN(n1957) );
  OR2_X1 U1510 ( .A1(n1457), .A2(n1480), .ZN(n1958) );
  OR2_X1 U1511 ( .A1(n1179), .A2(n1433), .ZN(n1959) );
  AND2_X1 U1512 ( .A1(n1123), .A2(n1132), .ZN(n1960) );
  AND2_X1 U1513 ( .A1(n1143), .A2(n1150), .ZN(n1961) );
  AND2_X1 U1514 ( .A1(n1151), .A2(n1158), .ZN(n1962) );
  BUF_X2 U1515 ( .A(a[13]), .Z(n2043) );
  XNOR2_X1 U1516 ( .A(a[22]), .B(a[21]), .ZN(n1963) );
  XNOR2_X1 U1517 ( .A(a[10]), .B(a[9]), .ZN(n1964) );
  AND2_X1 U1518 ( .A1(n1457), .A2(n1480), .ZN(n1965) );
  AND2_X1 U1519 ( .A1(n1179), .A2(n1433), .ZN(n1966) );
  AND2_X1 U1520 ( .A1(n1111), .A2(n1122), .ZN(n1967) );
  AND2_X1 U1521 ( .A1(n1133), .A2(n1142), .ZN(n1968) );
  AND2_X1 U1522 ( .A1(n1055), .A2(n1070), .ZN(n1969) );
  AND2_X1 U1523 ( .A1(n1021), .A2(n1038), .ZN(n1970) );
  OR2_X1 U1524 ( .A1(n1151), .A2(n1158), .ZN(n1971) );
  XNOR2_X1 U1525 ( .A(n560), .B(n1972), .ZN(product[22]) );
  AND2_X1 U1526 ( .A1(n2054), .A2(n559), .ZN(n1972) );
  XNOR2_X1 U1527 ( .A(n2108), .B(n1973), .ZN(product[34]) );
  AND2_X1 U1528 ( .A1(n2167), .A2(n439), .ZN(n1973) );
  BUF_X1 U1529 ( .A(n536), .Z(n1974) );
  BUF_X1 U1530 ( .A(n536), .Z(n1976) );
  BUF_X1 U1531 ( .A(n536), .Z(n1975) );
  INV_X2 U1532 ( .A(n2307), .ZN(n2025) );
  INV_X2 U1533 ( .A(n2307), .ZN(n2304) );
  INV_X1 U1534 ( .A(n2181), .ZN(n1978) );
  INV_X2 U1535 ( .A(n2140), .ZN(n2232) );
  INV_X1 U1536 ( .A(n554), .ZN(n1979) );
  NAND2_X2 U1537 ( .A1(n1806), .A2(n1963), .ZN(n1980) );
  XNOR2_X1 U1538 ( .A(a[6]), .B(a[7]), .ZN(n2136) );
  NAND2_X2 U1539 ( .A1(n1806), .A2(n1963), .ZN(n2130) );
  CLKBUF_X1 U1540 ( .A(n2290), .Z(n1982) );
  OAI22_X1 U1541 ( .A1(n2149), .A2(n1708), .B1(n1707), .B2(n2253), .ZN(n1983)
         );
  XNOR2_X1 U1542 ( .A(a[16]), .B(a[15]), .ZN(n1984) );
  BUF_X1 U1543 ( .A(n2159), .Z(n1985) );
  XNOR2_X1 U1544 ( .A(a[6]), .B(n2302), .ZN(n1987) );
  XNOR2_X1 U1545 ( .A(a[6]), .B(n2302), .ZN(n1986) );
  XNOR2_X1 U1546 ( .A(a[6]), .B(n2301), .ZN(n2168) );
  INV_X2 U1547 ( .A(n2133), .ZN(n1988) );
  INV_X1 U1548 ( .A(n2133), .ZN(n2237) );
  XNOR2_X1 U1549 ( .A(a[12]), .B(n2281), .ZN(n2111) );
  INV_X1 U1550 ( .A(n2246), .ZN(n1989) );
  INV_X1 U1551 ( .A(n2270), .ZN(n1990) );
  INV_X2 U1552 ( .A(n2196), .ZN(n2247) );
  INV_X1 U1553 ( .A(n2032), .ZN(n2196) );
  NOR2_X1 U1554 ( .A1(n513), .A2(n520), .ZN(n1991) );
  INV_X2 U1555 ( .A(n2302), .ZN(n2297) );
  INV_X1 U1556 ( .A(n2301), .ZN(n2298) );
  XOR2_X1 U1557 ( .A(a[20]), .B(a[19]), .Z(n2132) );
  CLKBUF_X3 U1558 ( .A(n285), .Z(n1993) );
  OAI22_X1 U1559 ( .A1(n2152), .A2(n1737), .B1(n1736), .B2(n2256), .ZN(n1994)
         );
  CLKBUF_X1 U1560 ( .A(n2259), .Z(n1995) );
  BUF_X2 U1561 ( .A(n2259), .Z(n1997) );
  CLKBUF_X2 U1562 ( .A(n2259), .Z(n1996) );
  BUF_X4 U1563 ( .A(b[0]), .Z(n1998) );
  CLKBUF_X1 U1564 ( .A(n2043), .Z(n1999) );
  INV_X1 U1565 ( .A(n2265), .ZN(n2000) );
  INV_X1 U1566 ( .A(n423), .ZN(n2001) );
  INV_X1 U1567 ( .A(n1936), .ZN(n2002) );
  INV_X1 U1568 ( .A(n2285), .ZN(n2004) );
  INV_X1 U1569 ( .A(n2285), .ZN(n2003) );
  BUF_X1 U1570 ( .A(n543), .Z(n2005) );
  CLKBUF_X3 U1571 ( .A(n2224), .Z(n2014) );
  BUF_X2 U1572 ( .A(n2224), .Z(n2015) );
  INV_X1 U1573 ( .A(n2143), .ZN(n2006) );
  INV_X1 U1574 ( .A(n2085), .ZN(n2143) );
  INV_X1 U1575 ( .A(n1992), .ZN(n2007) );
  AND2_X1 U1576 ( .A1(n1813), .A2(n2101), .ZN(n2008) );
  AND2_X1 U1577 ( .A1(n1813), .A2(n2101), .ZN(n2009) );
  XOR2_X1 U1578 ( .A(a[22]), .B(a[21]), .Z(n2010) );
  NOR2_X1 U1579 ( .A1(n513), .A2(n520), .ZN(n511) );
  INV_X1 U1580 ( .A(n2141), .ZN(n2011) );
  INV_X1 U1581 ( .A(n2051), .ZN(n2141) );
  BUF_X1 U1582 ( .A(n802), .Z(n2012) );
  CLKBUF_X1 U1583 ( .A(n2224), .Z(n2013) );
  INV_X1 U1584 ( .A(n2138), .ZN(n2224) );
  OAI22_X1 U1585 ( .A1(n2130), .A2(n1504), .B1(n2238), .B2(n1503), .ZN(n2016)
         );
  XNOR2_X1 U1586 ( .A(a[2]), .B(n2310), .ZN(n2017) );
  XNOR2_X1 U1587 ( .A(a[2]), .B(n2310), .ZN(n2146) );
  XNOR2_X1 U1588 ( .A(a[8]), .B(a[7]), .ZN(n2101) );
  CLKBUF_X1 U1589 ( .A(n2197), .Z(n2018) );
  OAI21_X1 U1590 ( .B1(n531), .B2(n535), .A(n532), .ZN(n2019) );
  NOR2_X1 U1591 ( .A1(n2021), .A2(n534), .ZN(n2020) );
  NOR2_X1 U1592 ( .A1(n877), .A2(n896), .ZN(n2021) );
  NOR2_X1 U1593 ( .A1(n2021), .A2(n534), .ZN(n525) );
  NOR2_X1 U1594 ( .A1(n877), .A2(n896), .ZN(n531) );
  CLKBUF_X1 U1595 ( .A(n568), .Z(n2022) );
  XNOR2_X1 U1596 ( .A(a[20]), .B(a[21]), .ZN(n2139) );
  XOR2_X1 U1597 ( .A(a[4]), .B(a[3]), .Z(n2137) );
  XNOR2_X1 U1598 ( .A(n906), .B(n2023), .ZN(n883) );
  XNOR2_X1 U1599 ( .A(n893), .B(n889), .ZN(n2023) );
  XOR2_X1 U1600 ( .A(n1949), .B(a[19]), .Z(n1808) );
  XOR2_X1 U1601 ( .A(a[16]), .B(a[15]), .Z(n2192) );
  NAND3_X1 U1602 ( .A1(n2062), .A2(n2063), .A3(n2064), .ZN(n2026) );
  INV_X1 U1603 ( .A(n2192), .ZN(n2245) );
  XOR2_X1 U1604 ( .A(n904), .B(n887), .Z(n2027) );
  XOR2_X1 U1605 ( .A(n902), .B(n2027), .Z(n881) );
  NAND2_X1 U1606 ( .A1(n902), .A2(n904), .ZN(n2028) );
  NAND2_X1 U1607 ( .A1(n902), .A2(n887), .ZN(n2029) );
  NAND2_X1 U1608 ( .A1(n904), .A2(n887), .ZN(n2030) );
  NAND3_X1 U1609 ( .A1(n2028), .A2(n2029), .A3(n2030), .ZN(n880) );
  INV_X1 U1610 ( .A(n2101), .ZN(n2181) );
  INV_X1 U1611 ( .A(n2186), .ZN(n2031) );
  XNOR2_X1 U1612 ( .A(a[14]), .B(a[13]), .ZN(n2032) );
  INV_X1 U1613 ( .A(n1988), .ZN(n2033) );
  INV_X2 U1614 ( .A(n2133), .ZN(n2236) );
  INV_X1 U1615 ( .A(n2014), .ZN(n2034) );
  XOR2_X1 U1616 ( .A(a[18]), .B(a[17]), .Z(n2197) );
  INV_X1 U1617 ( .A(n2290), .ZN(n2287) );
  INV_X1 U1618 ( .A(n2264), .ZN(n2262) );
  INV_X1 U1619 ( .A(n501), .ZN(n2035) );
  INV_X1 U1620 ( .A(n2109), .ZN(n2037) );
  INV_X1 U1621 ( .A(n2109), .ZN(n2036) );
  INV_X1 U1622 ( .A(n2109), .ZN(n2249) );
  XNOR2_X1 U1623 ( .A(n2038), .B(n953), .ZN(n947) );
  XNOR2_X1 U1624 ( .A(n972), .B(n959), .ZN(n2038) );
  XNOR2_X1 U1625 ( .A(n2039), .B(n966), .ZN(n943) );
  XNOR2_X1 U1626 ( .A(n947), .B(n949), .ZN(n2039) );
  NAND3_X1 U1627 ( .A1(n2211), .A2(n2212), .A3(n2213), .ZN(n2040) );
  INV_X1 U1628 ( .A(a[21]), .ZN(n2264) );
  CLKBUF_X1 U1629 ( .A(n2100), .Z(n2041) );
  INV_X1 U1630 ( .A(n917), .ZN(n2042) );
  INV_X2 U1631 ( .A(n2146), .ZN(n2256) );
  XOR2_X1 U1632 ( .A(n1363), .B(n1209), .Z(n2044) );
  XOR2_X1 U1633 ( .A(n2044), .B(n2221), .Z(n819) );
  NAND2_X1 U1634 ( .A1(n1363), .A2(n1209), .ZN(n2045) );
  NAND2_X1 U1635 ( .A1(n1363), .A2(n2221), .ZN(n2046) );
  NAND2_X1 U1636 ( .A1(n1209), .A2(n2221), .ZN(n2047) );
  NAND3_X1 U1637 ( .A1(n2045), .A2(n2046), .A3(n2047), .ZN(n818) );
  NAND2_X1 U1638 ( .A1(n1274), .A2(n1296), .ZN(n2048) );
  NAND2_X1 U1639 ( .A1(n1274), .A2(n818), .ZN(n2049) );
  NAND2_X1 U1640 ( .A1(n1296), .A2(n818), .ZN(n2050) );
  NAND3_X1 U1641 ( .A1(n2048), .A2(n2049), .A3(n2050), .ZN(n796) );
  OR2_X2 U1642 ( .A1(n2142), .A2(n2017), .ZN(n2051) );
  NOR2_X1 U1643 ( .A1(n839), .A2(n856), .ZN(n2052) );
  NOR2_X1 U1644 ( .A1(n2139), .A2(n2132), .ZN(n2138) );
  INV_X1 U1645 ( .A(n1964), .ZN(n2109) );
  INV_X1 U1646 ( .A(n2135), .ZN(n2053) );
  INV_X1 U1647 ( .A(n1936), .ZN(n2288) );
  XNOR2_X1 U1648 ( .A(a[10]), .B(n2284), .ZN(n1812) );
  INV_X1 U1649 ( .A(n2285), .ZN(n2283) );
  OR2_X1 U1650 ( .A1(n963), .A2(n982), .ZN(n2054) );
  INV_X2 U1651 ( .A(n2140), .ZN(n2057) );
  INV_X1 U1652 ( .A(n2140), .ZN(n2056) );
  INV_X1 U1653 ( .A(n2009), .ZN(n2234) );
  CLKBUF_X1 U1654 ( .A(n581), .Z(n2058) );
  NOR2_X1 U1655 ( .A1(n820), .A2(n805), .ZN(n2059) );
  NOR2_X1 U1656 ( .A1(n805), .A2(n820), .ZN(n495) );
  OR2_X2 U1657 ( .A1(n2136), .A2(n2168), .ZN(n2100) );
  OR2_X2 U1658 ( .A1(n2136), .A2(n1987), .ZN(n2074) );
  CLKBUF_X1 U1659 ( .A(n535), .Z(n2060) );
  XOR2_X1 U1660 ( .A(n1438), .B(n1284), .Z(n2061) );
  XOR2_X1 U1661 ( .A(n1372), .B(n2061), .Z(n997) );
  NAND2_X1 U1662 ( .A1(n1372), .A2(n1994), .ZN(n2062) );
  NAND2_X1 U1663 ( .A1(n1372), .A2(n1284), .ZN(n2063) );
  NAND2_X1 U1664 ( .A1(n1994), .A2(n1284), .ZN(n2064) );
  NAND3_X1 U1665 ( .A1(n2062), .A2(n2063), .A3(n2064), .ZN(n996) );
  XOR2_X1 U1666 ( .A(n863), .B(n882), .Z(n2065) );
  XOR2_X1 U1667 ( .A(n880), .B(n2065), .Z(n859) );
  NAND2_X1 U1668 ( .A1(n880), .A2(n863), .ZN(n2066) );
  NAND2_X1 U1669 ( .A1(n880), .A2(n882), .ZN(n2067) );
  NAND2_X1 U1670 ( .A1(n863), .A2(n882), .ZN(n2068) );
  NAND3_X1 U1671 ( .A1(n2066), .A2(n2067), .A3(n2068), .ZN(n858) );
  XNOR2_X1 U1672 ( .A(a[14]), .B(n2278), .ZN(n1810) );
  INV_X1 U1673 ( .A(n1934), .ZN(n2275) );
  XNOR2_X1 U1674 ( .A(a[11]), .B(a[12]), .ZN(n2069) );
  INV_X2 U1675 ( .A(n2191), .ZN(n2248) );
  XNOR2_X1 U1676 ( .A(n2024), .B(n2272), .ZN(n1809) );
  XNOR2_X1 U1677 ( .A(n2070), .B(n1042), .ZN(n1023) );
  XNOR2_X1 U1678 ( .A(n1027), .B(n1044), .ZN(n2070) );
  BUF_X1 U1679 ( .A(n2228), .Z(n2154) );
  OAI21_X1 U1680 ( .B1(n503), .B2(n2059), .A(n496), .ZN(n2071) );
  NOR2_X1 U1681 ( .A1(n547), .A2(n542), .ZN(n2072) );
  CLKBUF_X1 U1682 ( .A(n839), .Z(n2073) );
  BUF_X2 U1683 ( .A(n2228), .Z(n2156) );
  AND2_X2 U1684 ( .A1(n2111), .A2(n2069), .ZN(n2140) );
  INV_X1 U1685 ( .A(n2074), .ZN(n2135) );
  BUF_X2 U1686 ( .A(n2228), .Z(n2155) );
  XOR2_X1 U1687 ( .A(n933), .B(n937), .Z(n2075) );
  XOR2_X1 U1688 ( .A(n2075), .B(n952), .Z(n927) );
  NAND2_X1 U1689 ( .A1(n933), .A2(n937), .ZN(n2076) );
  NAND2_X1 U1690 ( .A1(n933), .A2(n952), .ZN(n2077) );
  NAND2_X1 U1691 ( .A1(n937), .A2(n952), .ZN(n2078) );
  NAND3_X1 U1692 ( .A1(n2076), .A2(n2077), .A3(n2078), .ZN(n926) );
  XOR2_X1 U1693 ( .A(n907), .B(n905), .Z(n2079) );
  XOR2_X1 U1694 ( .A(n2079), .B(n926), .Z(n901) );
  NAND2_X1 U1695 ( .A1(n907), .A2(n905), .ZN(n2080) );
  NAND2_X1 U1696 ( .A1(n907), .A2(n926), .ZN(n2081) );
  NAND2_X1 U1697 ( .A1(n905), .A2(n926), .ZN(n2082) );
  NAND3_X1 U1698 ( .A1(n2080), .A2(n2081), .A3(n2082), .ZN(n900) );
  XOR2_X1 U1699 ( .A(n1238), .B(n1216), .Z(n2083) );
  OAI21_X1 U1700 ( .B1(n531), .B2(n535), .A(n532), .ZN(n526) );
  CLKBUF_X1 U1701 ( .A(n490), .Z(n2084) );
  OR2_X2 U1702 ( .A1(n2137), .A2(n2144), .ZN(n2085) );
  XOR2_X1 U1703 ( .A(n1062), .B(n1053), .Z(n2086) );
  XOR2_X1 U1704 ( .A(n2086), .B(n1060), .Z(n1043) );
  NAND2_X1 U1705 ( .A1(n1062), .A2(n1053), .ZN(n2087) );
  NAND2_X1 U1706 ( .A1(n1062), .A2(n1060), .ZN(n2088) );
  NAND2_X1 U1707 ( .A1(n1053), .A2(n1060), .ZN(n2089) );
  NAND3_X1 U1708 ( .A1(n2087), .A2(n2088), .A3(n2089), .ZN(n1042) );
  NAND2_X1 U1709 ( .A1(n1027), .A2(n1044), .ZN(n2090) );
  NAND2_X1 U1710 ( .A1(n1027), .A2(n1042), .ZN(n2091) );
  NAND2_X1 U1711 ( .A1(n1044), .A2(n1042), .ZN(n2092) );
  NAND3_X1 U1712 ( .A1(n2090), .A2(n2091), .A3(n2092), .ZN(n1022) );
  XOR2_X1 U1713 ( .A(n964), .B(n945), .Z(n2093) );
  XOR2_X1 U1714 ( .A(n2093), .B(n943), .Z(n941) );
  NAND2_X1 U1715 ( .A1(n947), .A2(n949), .ZN(n2094) );
  NAND2_X1 U1716 ( .A1(n966), .A2(n947), .ZN(n2095) );
  NAND2_X1 U1717 ( .A1(n949), .A2(n966), .ZN(n2096) );
  NAND3_X1 U1718 ( .A1(n2094), .A2(n2095), .A3(n2096), .ZN(n942) );
  NAND2_X1 U1719 ( .A1(n964), .A2(n945), .ZN(n2097) );
  NAND2_X1 U1720 ( .A1(n964), .A2(n943), .ZN(n2098) );
  NAND2_X1 U1721 ( .A1(n945), .A2(n943), .ZN(n2099) );
  NAND3_X1 U1722 ( .A1(n2097), .A2(n2098), .A3(n2099), .ZN(n940) );
  AND2_X2 U1723 ( .A1(n1810), .A2(n2032), .ZN(n2134) );
  XNOR2_X1 U1724 ( .A(a[22]), .B(n2261), .ZN(n1806) );
  INV_X2 U1725 ( .A(n2181), .ZN(n2250) );
  XOR2_X1 U1726 ( .A(n1309), .B(n1464), .Z(n2102) );
  XOR2_X1 U1727 ( .A(n2102), .B(n1287), .Z(n1053) );
  NAND2_X1 U1728 ( .A1(n1287), .A2(n1309), .ZN(n2103) );
  NAND2_X1 U1729 ( .A1(n1287), .A2(n1464), .ZN(n2104) );
  NAND2_X1 U1730 ( .A1(n1309), .A2(n1464), .ZN(n2105) );
  NAND3_X1 U1731 ( .A1(n2103), .A2(n2104), .A3(n2105), .ZN(n1052) );
  AOI21_X1 U1732 ( .B1(n2058), .B2(n567), .A(n2022), .ZN(n2106) );
  INV_X2 U1733 ( .A(n2145), .ZN(n2227) );
  AND2_X2 U1734 ( .A1(n1809), .A2(n1984), .ZN(n2145) );
  AND2_X1 U1735 ( .A1(n2219), .A2(n2220), .ZN(n2108) );
  AND2_X1 U1736 ( .A1(n2219), .A2(n2220), .ZN(n2215) );
  NOR2_X1 U1737 ( .A1(n695), .A2(n700), .ZN(n384) );
  OR2_X1 U1738 ( .A1(n717), .A2(n726), .ZN(n2118) );
  OR2_X1 U1739 ( .A1(n709), .A2(n716), .ZN(n2119) );
  OR2_X1 U1740 ( .A1(n1143), .A2(n1150), .ZN(n2110) );
  INV_X2 U1741 ( .A(n2267), .ZN(n2265) );
  NOR2_X1 U1742 ( .A1(n2186), .A2(n467), .ZN(n465) );
  INV_X1 U1743 ( .A(n435), .ZN(n662) );
  OAI21_X1 U1744 ( .B1(n492), .B2(n467), .A(n468), .ZN(n466) );
  INV_X1 U1745 ( .A(n481), .ZN(n483) );
  NAND2_X1 U1746 ( .A1(n666), .A2(n481), .ZN(n315) );
  NAND2_X1 U1747 ( .A1(n667), .A2(n496), .ZN(n316) );
  NAND2_X1 U1748 ( .A1(n671), .A2(n532), .ZN(n320) );
  NAND2_X1 U1749 ( .A1(n662), .A2(n436), .ZN(n311) );
  INV_X1 U1750 ( .A(n2167), .ZN(n438) );
  AOI21_X1 U1751 ( .B1(n565), .B2(n561), .A(n562), .ZN(n560) );
  INV_X1 U1752 ( .A(n439), .ZN(n445) );
  XOR2_X1 U1753 ( .A(n551), .B(n323), .Z(product[23]) );
  AOI21_X1 U1754 ( .B1(n662), .B2(n445), .A(n434), .ZN(n432) );
  INV_X1 U1755 ( .A(n436), .ZN(n434) );
  NOR2_X1 U1756 ( .A1(n402), .A2(n360), .ZN(n356) );
  INV_X1 U1757 ( .A(n563), .ZN(n561) );
  INV_X1 U1758 ( .A(n564), .ZN(n562) );
  NAND2_X1 U1759 ( .A1(n2167), .A2(n662), .ZN(n431) );
  INV_X1 U1760 ( .A(n382), .ZN(n380) );
  AOI21_X1 U1761 ( .B1(n426), .B2(n445), .A(n427), .ZN(n421) );
  NOR2_X1 U1762 ( .A1(n737), .A2(n748), .ZN(n435) );
  AOI21_X1 U1763 ( .B1(n2119), .B2(n416), .A(n407), .ZN(n405) );
  INV_X1 U1764 ( .A(n409), .ZN(n407) );
  NOR2_X1 U1765 ( .A1(n384), .A2(n364), .ZN(n362) );
  OAI21_X1 U1766 ( .B1(n590), .B2(n593), .A(n591), .ZN(n589) );
  AND2_X1 U1767 ( .A1(n1039), .A2(n1054), .ZN(n2112) );
  NAND2_X1 U1768 ( .A1(n657), .A2(n387), .ZN(n306) );
  INV_X1 U1769 ( .A(n384), .ZN(n657) );
  NOR2_X1 U1770 ( .A1(n963), .A2(n982), .ZN(n558) );
  NAND2_X1 U1771 ( .A1(n789), .A2(n804), .ZN(n481) );
  NOR2_X1 U1772 ( .A1(n1071), .A2(n1084), .ZN(n590) );
  NOR2_X1 U1773 ( .A1(n435), .A2(n428), .ZN(n426) );
  NAND2_X1 U1774 ( .A1(n737), .A2(n748), .ZN(n436) );
  NAND2_X1 U1775 ( .A1(n2185), .A2(n514), .ZN(n318) );
  NAND2_X1 U1776 ( .A1(n2119), .A2(n409), .ZN(n308) );
  NAND2_X1 U1777 ( .A1(n422), .A2(n2118), .ZN(n411) );
  NAND2_X1 U1778 ( .A1(n2120), .A2(n396), .ZN(n307) );
  NAND2_X1 U1779 ( .A1(n661), .A2(n429), .ZN(n310) );
  AOI21_X1 U1780 ( .B1(n565), .B2(n545), .A(n546), .ZN(n544) );
  OR2_X1 U1781 ( .A1(n761), .A2(n774), .ZN(n2113) );
  AOI21_X1 U1782 ( .B1(n423), .B2(n2118), .A(n416), .ZN(n412) );
  NOR2_X1 U1783 ( .A1(n389), .A2(n384), .ZN(n382) );
  INV_X1 U1784 ( .A(n396), .ZN(n394) );
  NAND2_X1 U1785 ( .A1(n362), .A2(n2120), .ZN(n360) );
  NAND2_X1 U1786 ( .A1(n821), .A2(n838), .ZN(n503) );
  INV_X1 U1787 ( .A(n378), .ZN(n376) );
  NAND2_X1 U1788 ( .A1(n2118), .A2(n2119), .ZN(n402) );
  OR2_X1 U1789 ( .A1(n1039), .A2(n1054), .ZN(n2114) );
  OR2_X1 U1790 ( .A1(n1055), .A2(n1070), .ZN(n2115) );
  XNOR2_X1 U1791 ( .A(n859), .B(n2116), .ZN(n857) );
  XNOR2_X1 U1792 ( .A(n878), .B(n861), .ZN(n2116) );
  XNOR2_X1 U1793 ( .A(n1041), .B(n2117), .ZN(n1039) );
  XNOR2_X1 U1794 ( .A(n1056), .B(n1043), .ZN(n2117) );
  INV_X1 U1795 ( .A(n352), .ZN(n350) );
  OAI21_X1 U1796 ( .B1(n628), .B2(n626), .A(n627), .ZN(n625) );
  OR2_X2 U1797 ( .A1(n701), .A2(n708), .ZN(n2120) );
  OAI21_X1 U1798 ( .B1(n405), .B2(n360), .A(n361), .ZN(n359) );
  AOI21_X1 U1799 ( .B1(n362), .B2(n394), .A(n363), .ZN(n361) );
  OAI21_X1 U1800 ( .B1(n364), .B2(n387), .A(n365), .ZN(n363) );
  AOI21_X1 U1801 ( .B1(n376), .B2(n2125), .A(n367), .ZN(n365) );
  AOI21_X1 U1802 ( .B1(n2122), .B2(n1960), .A(n1967), .ZN(n600) );
  OR2_X1 U1803 ( .A1(n1133), .A2(n1142), .ZN(n2121) );
  AOI21_X1 U1804 ( .B1(n629), .B2(n635), .A(n630), .ZN(n628) );
  OAI21_X1 U1805 ( .B1(n638), .B2(n636), .A(n637), .ZN(n635) );
  NOR2_X1 U1806 ( .A1(n633), .A2(n631), .ZN(n629) );
  OAI21_X1 U1807 ( .B1(n631), .B2(n634), .A(n632), .ZN(n630) );
  NAND2_X1 U1808 ( .A1(n2125), .A2(n369), .ZN(n304) );
  NAND2_X1 U1809 ( .A1(n2127), .A2(n341), .ZN(n302) );
  NAND2_X1 U1810 ( .A1(n2126), .A2(n352), .ZN(n303) );
  NAND2_X1 U1811 ( .A1(n695), .A2(n700), .ZN(n387) );
  AOI21_X1 U1812 ( .B1(n2121), .B2(n1961), .A(n1968), .ZN(n611) );
  OR2_X1 U1813 ( .A1(n1111), .A2(n1122), .ZN(n2122) );
  INV_X1 U1814 ( .A(n369), .ZN(n367) );
  OR2_X1 U1815 ( .A1(n694), .A2(n689), .ZN(n2123) );
  NAND2_X1 U1816 ( .A1(n2110), .A2(n2121), .ZN(n610) );
  NAND2_X1 U1817 ( .A1(n1085), .A2(n1098), .ZN(n593) );
  OR2_X1 U1818 ( .A1(n1123), .A2(n1132), .ZN(n2124) );
  INV_X1 U1819 ( .A(n2311), .ZN(n2308) );
  NOR2_X1 U1820 ( .A1(n1165), .A2(n1170), .ZN(n631) );
  NAND2_X1 U1821 ( .A1(n678), .A2(n677), .ZN(n335) );
  INV_X1 U1822 ( .A(n341), .ZN(n339) );
  AOI21_X1 U1823 ( .B1(n643), .B2(n1959), .A(n1966), .ZN(n638) );
  OAI21_X1 U1824 ( .B1(n646), .B2(n644), .A(n645), .ZN(n643) );
  AOI21_X1 U1825 ( .B1(n1958), .B2(n1957), .A(n1965), .ZN(n646) );
  OR2_X1 U1826 ( .A1(n685), .A2(n688), .ZN(n2125) );
  BUF_X2 U1827 ( .A(n2032), .Z(n2150) );
  NOR2_X1 U1828 ( .A1(n1175), .A2(n1178), .ZN(n636) );
  OR2_X1 U1829 ( .A1(n681), .A2(n684), .ZN(n2126) );
  NOR2_X1 U1830 ( .A1(n1159), .A2(n1161), .ZN(n626) );
  OR2_X1 U1831 ( .A1(n679), .A2(n680), .ZN(n2127) );
  NAND2_X1 U1832 ( .A1(n681), .A2(n684), .ZN(n352) );
  NAND2_X1 U1833 ( .A1(n679), .A2(n680), .ZN(n341) );
  NAND2_X1 U1834 ( .A1(n1175), .A2(n1178), .ZN(n637) );
  NAND2_X1 U1835 ( .A1(n1159), .A2(n1161), .ZN(n627) );
  INV_X1 U1836 ( .A(n676), .ZN(n677) );
  OR2_X1 U1837 ( .A1(n1194), .A2(n676), .ZN(n2128) );
  NOR2_X1 U1838 ( .A1(n678), .A2(n677), .ZN(n334) );
  AND2_X1 U1839 ( .A1(n1194), .A2(n676), .ZN(n2129) );
  INV_X1 U1840 ( .A(n2278), .ZN(n2276) );
  INV_X1 U1841 ( .A(n2302), .ZN(n2299) );
  INV_X1 U1842 ( .A(n2261), .ZN(n2259) );
  INV_X1 U1843 ( .A(n2010), .ZN(n2238) );
  INV_X1 U1844 ( .A(n1507), .ZN(n2323) );
  INV_X1 U1845 ( .A(n682), .ZN(n683) );
  INV_X1 U1846 ( .A(n2017), .ZN(n2255) );
  INV_X1 U1847 ( .A(n2132), .ZN(n2241) );
  INV_X1 U1848 ( .A(n1986), .ZN(n2252) );
  INV_X1 U1849 ( .A(n1992), .ZN(n2240) );
  INV_X1 U1850 ( .A(n2010), .ZN(n2239) );
  INV_X1 U1851 ( .A(n2197), .ZN(n2242) );
  OAI21_X1 U1852 ( .B1(n2141), .B2(n2017), .A(n2314), .ZN(n1434) );
  NAND2_X1 U1853 ( .A1(n1181), .A2(n1192), .ZN(n645) );
  NOR2_X1 U1854 ( .A1(n1181), .A2(n1192), .ZN(n644) );
  INV_X1 U1855 ( .A(n692), .ZN(n693) );
  OAI22_X1 U1856 ( .A1(n1955), .A2(n1586), .B1(n2247), .B2(n1585), .ZN(n1293)
         );
  INV_X1 U1857 ( .A(n1532), .ZN(n2322) );
  OAI22_X1 U1858 ( .A1(n2230), .A2(n1584), .B1(n2247), .B2(n1583), .ZN(n1291)
         );
  OAI22_X1 U1859 ( .A1(n1955), .A2(n1592), .B1(n2150), .B2(n1591), .ZN(n1299)
         );
  OAI22_X1 U1860 ( .A1(n1955), .A2(n1588), .B1(n2247), .B2(n1587), .ZN(n1295)
         );
  OAI22_X1 U1861 ( .A1(n2230), .A2(n1590), .B1(n2247), .B2(n1589), .ZN(n1297)
         );
  INV_X1 U1862 ( .A(n1707), .ZN(n2315) );
  INV_X1 U1863 ( .A(n1682), .ZN(n2316) );
  INV_X1 U1864 ( .A(n1557), .ZN(n2321) );
  INV_X1 U1865 ( .A(n1607), .ZN(n2319) );
  OAI22_X1 U1866 ( .A1(n2226), .A2(n1538), .B1(n2244), .B2(n1537), .ZN(n1247)
         );
  INV_X1 U1867 ( .A(n724), .ZN(n725) );
  CLKBUF_X1 U1868 ( .A(n251), .Z(n2258) );
  INV_X1 U1869 ( .A(n1732), .ZN(n2314) );
  INV_X1 U1870 ( .A(n1582), .ZN(n2320) );
  INV_X1 U1871 ( .A(n1632), .ZN(n2318) );
  INV_X1 U1872 ( .A(n1657), .ZN(n2317) );
  INV_X1 U1873 ( .A(n1482), .ZN(n2324) );
  XNOR2_X1 U1874 ( .A(n2294), .B(b[22]), .ZN(n1683) );
  XNOR2_X1 U1875 ( .A(n2275), .B(b[16]), .ZN(n1589) );
  XNOR2_X1 U1876 ( .A(n2265), .B(b[18]), .ZN(n1537) );
  XNOR2_X1 U1877 ( .A(n2277), .B(b[14]), .ZN(n1591) );
  XNOR2_X1 U1878 ( .A(n2276), .B(b[22]), .ZN(n1583) );
  XNOR2_X1 U1879 ( .A(n2274), .B(b[18]), .ZN(n1587) );
  XNOR2_X1 U1880 ( .A(n2277), .B(b[20]), .ZN(n1585) );
  XNOR2_X1 U1881 ( .A(n2309), .B(b[22]), .ZN(n1758) );
  XNOR2_X1 U1882 ( .A(n2308), .B(b[18]), .ZN(n1762) );
  XNOR2_X1 U1883 ( .A(n2309), .B(b[16]), .ZN(n1764) );
  XNOR2_X1 U1884 ( .A(n2308), .B(b[10]), .ZN(n1770) );
  XNOR2_X1 U1885 ( .A(n2308), .B(b[14]), .ZN(n1766) );
  XNOR2_X1 U1886 ( .A(n2308), .B(b[6]), .ZN(n1774) );
  XNOR2_X1 U1887 ( .A(n2308), .B(b[8]), .ZN(n1772) );
  XNOR2_X1 U1888 ( .A(n2308), .B(b[4]), .ZN(n1776) );
  XNOR2_X1 U1889 ( .A(n2263), .B(b[18]), .ZN(n1512) );
  XNOR2_X1 U1890 ( .A(n2002), .B(b[16]), .ZN(n1664) );
  XNOR2_X1 U1891 ( .A(n2293), .B(b[18]), .ZN(n1687) );
  XNOR2_X1 U1892 ( .A(n2262), .B(b[4]), .ZN(n1526) );
  XNOR2_X1 U1893 ( .A(n2280), .B(b[14]), .ZN(n1616) );
  XNOR2_X1 U1894 ( .A(n2289), .B(b[18]), .ZN(n1662) );
  XNOR2_X1 U1895 ( .A(n2270), .B(b[8]), .ZN(n1572) );
  XNOR2_X1 U1896 ( .A(n2270), .B(b[10]), .ZN(n1570) );
  XNOR2_X1 U1897 ( .A(n2271), .B(b[22]), .ZN(n1558) );
  XNOR2_X1 U1898 ( .A(n1977), .B(b[16]), .ZN(n1514) );
  XNOR2_X1 U1899 ( .A(n2265), .B(b[4]), .ZN(n1551) );
  XNOR2_X1 U1900 ( .A(n2270), .B(b[14]), .ZN(n1566) );
  XNOR2_X1 U1901 ( .A(n2043), .B(b[16]), .ZN(n1614) );
  XNOR2_X1 U1902 ( .A(n2265), .B(b[10]), .ZN(n1545) );
  XNOR2_X1 U1903 ( .A(n2274), .B(b[10]), .ZN(n1595) );
  XNOR2_X1 U1904 ( .A(n2004), .B(b[18]), .ZN(n1637) );
  XNOR2_X1 U1905 ( .A(n2263), .B(b[8]), .ZN(n1522) );
  XNOR2_X1 U1906 ( .A(n2280), .B(b[10]), .ZN(n1620) );
  XNOR2_X1 U1907 ( .A(n2265), .B(b[8]), .ZN(n1547) );
  XNOR2_X1 U1908 ( .A(n2283), .B(b[16]), .ZN(n1639) );
  XNOR2_X1 U1909 ( .A(n2266), .B(b[22]), .ZN(n1533) );
  XNOR2_X1 U1910 ( .A(n2270), .B(b[6]), .ZN(n1574) );
  XNOR2_X1 U1911 ( .A(n2287), .B(b[14]), .ZN(n1666) );
  XNOR2_X1 U1912 ( .A(n2276), .B(b[8]), .ZN(n1597) );
  XNOR2_X1 U1913 ( .A(n2294), .B(b[16]), .ZN(n1689) );
  XNOR2_X1 U1914 ( .A(n2280), .B(b[18]), .ZN(n1612) );
  XNOR2_X1 U1915 ( .A(n2263), .B(b[10]), .ZN(n1520) );
  XNOR2_X1 U1916 ( .A(n2282), .B(b[14]), .ZN(n1641) );
  XNOR2_X1 U1917 ( .A(n2265), .B(b[6]), .ZN(n1549) );
  XNOR2_X1 U1918 ( .A(n2299), .B(b[18]), .ZN(n1712) );
  XNOR2_X1 U1919 ( .A(n2288), .B(b[22]), .ZN(n1658) );
  XNOR2_X1 U1920 ( .A(n2305), .B(b[22]), .ZN(n1733) );
  XNOR2_X1 U1921 ( .A(n2265), .B(b[14]), .ZN(n1541) );
  XNOR2_X1 U1922 ( .A(n2263), .B(b[6]), .ZN(n1524) );
  XNOR2_X1 U1923 ( .A(n2003), .B(b[22]), .ZN(n1633) );
  XNOR2_X1 U1924 ( .A(n2025), .B(b[18]), .ZN(n1737) );
  XNOR2_X1 U1925 ( .A(n2293), .B(b[14]), .ZN(n1691) );
  XNOR2_X1 U1926 ( .A(n2270), .B(b[4]), .ZN(n1576) );
  XNOR2_X1 U1927 ( .A(n2271), .B(b[16]), .ZN(n1564) );
  XNOR2_X1 U1928 ( .A(n2300), .B(b[16]), .ZN(n1714) );
  XNOR2_X1 U1929 ( .A(n2275), .B(b[6]), .ZN(n1599) );
  XNOR2_X1 U1930 ( .A(n2280), .B(b[8]), .ZN(n1622) );
  XNOR2_X1 U1931 ( .A(n2270), .B(b[18]), .ZN(n1562) );
  XNOR2_X1 U1932 ( .A(n2300), .B(b[22]), .ZN(n1708) );
  XNOR2_X1 U1933 ( .A(n2266), .B(b[16]), .ZN(n1539) );
  XNOR2_X1 U1934 ( .A(n2263), .B(b[14]), .ZN(n1516) );
  XNOR2_X1 U1935 ( .A(n2282), .B(b[10]), .ZN(n1645) );
  XNOR2_X1 U1936 ( .A(n2043), .B(b[22]), .ZN(n1608) );
  XNOR2_X1 U1937 ( .A(n2283), .B(b[4]), .ZN(n1651) );
  XNOR2_X1 U1938 ( .A(n2004), .B(b[6]), .ZN(n1649) );
  XNOR2_X1 U1939 ( .A(n2003), .B(b[8]), .ZN(n1647) );
  XNOR2_X1 U1940 ( .A(n2276), .B(b[4]), .ZN(n1601) );
  XNOR2_X1 U1941 ( .A(n2287), .B(b[10]), .ZN(n1670) );
  XNOR2_X1 U1942 ( .A(n2025), .B(b[14]), .ZN(n1741) );
  XNOR2_X1 U1943 ( .A(n2002), .B(b[8]), .ZN(n1672) );
  XNOR2_X1 U1944 ( .A(n2299), .B(b[6]), .ZN(n1724) );
  XNOR2_X1 U1945 ( .A(n2280), .B(b[6]), .ZN(n1624) );
  XNOR2_X1 U1946 ( .A(n2293), .B(b[8]), .ZN(n1697) );
  XNOR2_X1 U1947 ( .A(n2002), .B(b[6]), .ZN(n1674) );
  XNOR2_X1 U1948 ( .A(n2280), .B(b[4]), .ZN(n1626) );
  XNOR2_X1 U1949 ( .A(n2293), .B(b[10]), .ZN(n1695) );
  XNOR2_X1 U1950 ( .A(n2025), .B(b[16]), .ZN(n1739) );
  XNOR2_X1 U1951 ( .A(n2025), .B(b[4]), .ZN(n1751) );
  XNOR2_X1 U1952 ( .A(n2293), .B(b[4]), .ZN(n1701) );
  XNOR2_X1 U1953 ( .A(n2299), .B(b[14]), .ZN(n1716) );
  XNOR2_X1 U1954 ( .A(n2299), .B(b[4]), .ZN(n1726) );
  XNOR2_X1 U1955 ( .A(n2304), .B(b[10]), .ZN(n1745) );
  XNOR2_X1 U1956 ( .A(n2304), .B(b[6]), .ZN(n1749) );
  XNOR2_X1 U1957 ( .A(n2287), .B(b[4]), .ZN(n1676) );
  XNOR2_X1 U1958 ( .A(n2299), .B(b[8]), .ZN(n1722) );
  XNOR2_X1 U1959 ( .A(n2293), .B(b[6]), .ZN(n1699) );
  XNOR2_X1 U1960 ( .A(n2304), .B(b[8]), .ZN(n1747) );
  XNOR2_X1 U1961 ( .A(n1977), .B(b[22]), .ZN(n1508) );
  XNOR2_X1 U1962 ( .A(n2299), .B(b[10]), .ZN(n1720) );
  XNOR2_X1 U1963 ( .A(b[23]), .B(n2003), .ZN(n1632) );
  XNOR2_X1 U1964 ( .A(n2309), .B(b[20]), .ZN(n1760) );
  XNOR2_X1 U1965 ( .A(n2308), .B(b[2]), .ZN(n1778) );
  XNOR2_X1 U1966 ( .A(n2308), .B(b[12]), .ZN(n1768) );
  XNOR2_X1 U1967 ( .A(n2266), .B(b[20]), .ZN(n1535) );
  XNOR2_X1 U1968 ( .A(n2274), .B(b[12]), .ZN(n1593) );
  XNOR2_X1 U1969 ( .A(n2294), .B(b[20]), .ZN(n1685) );
  XNOR2_X1 U1970 ( .A(n2282), .B(b[12]), .ZN(n1643) );
  XNOR2_X1 U1971 ( .A(n2271), .B(b[20]), .ZN(n1560) );
  XNOR2_X1 U1972 ( .A(n2265), .B(b[12]), .ZN(n1543) );
  XNOR2_X1 U1973 ( .A(n2003), .B(b[20]), .ZN(n1635) );
  XNOR2_X1 U1974 ( .A(n2270), .B(b[12]), .ZN(n1568) );
  XNOR2_X1 U1975 ( .A(n2305), .B(b[20]), .ZN(n1735) );
  XNOR2_X1 U1976 ( .A(n2280), .B(b[12]), .ZN(n1618) );
  XNOR2_X1 U1977 ( .A(n2263), .B(b[20]), .ZN(n1510) );
  XNOR2_X1 U1978 ( .A(n1977), .B(b[12]), .ZN(n1518) );
  XNOR2_X1 U1979 ( .A(n2288), .B(b[20]), .ZN(n1660) );
  XNOR2_X1 U1980 ( .A(n2043), .B(b[20]), .ZN(n1610) );
  XNOR2_X1 U1981 ( .A(n2265), .B(b[2]), .ZN(n1553) );
  XNOR2_X1 U1982 ( .A(n2280), .B(b[2]), .ZN(n1628) );
  XNOR2_X1 U1983 ( .A(n2293), .B(b[12]), .ZN(n1693) );
  XNOR2_X1 U1984 ( .A(n2283), .B(b[2]), .ZN(n1653) );
  XNOR2_X1 U1985 ( .A(n2276), .B(b[2]), .ZN(n1603) );
  XNOR2_X1 U1986 ( .A(n2299), .B(b[12]), .ZN(n1718) );
  XNOR2_X1 U1987 ( .A(n2270), .B(b[2]), .ZN(n1578) );
  XNOR2_X1 U1988 ( .A(n2293), .B(b[2]), .ZN(n1703) );
  XNOR2_X1 U1989 ( .A(n2304), .B(b[12]), .ZN(n1743) );
  XNOR2_X1 U1990 ( .A(n2288), .B(b[2]), .ZN(n1678) );
  XNOR2_X1 U1991 ( .A(n2299), .B(b[2]), .ZN(n1728) );
  XNOR2_X1 U1992 ( .A(n2304), .B(b[2]), .ZN(n1753) );
  XNOR2_X1 U1993 ( .A(b[5]), .B(n2004), .ZN(n1650) );
  XNOR2_X1 U1994 ( .A(b[3]), .B(n2004), .ZN(n1652) );
  AND2_X2 U1995 ( .A1(n1808), .A2(n2242), .ZN(n2131) );
  XNOR2_X1 U1996 ( .A(b[23]), .B(n2305), .ZN(n1732) );
  XNOR2_X1 U1997 ( .A(b[23]), .B(n2269), .ZN(n1557) );
  XNOR2_X1 U1998 ( .A(b[23]), .B(n1999), .ZN(n1607) );
  XNOR2_X1 U1999 ( .A(b[23]), .B(n2288), .ZN(n1657) );
  XNOR2_X1 U2000 ( .A(b[23]), .B(n1981), .ZN(n1532) );
  XNOR2_X1 U2001 ( .A(b[9]), .B(n2269), .ZN(n1571) );
  XNOR2_X1 U2002 ( .A(b[1]), .B(n1995), .ZN(n1504) );
  XNOR2_X1 U2003 ( .A(b[7]), .B(n1981), .ZN(n1548) );
  XNOR2_X1 U2004 ( .A(b[9]), .B(n1981), .ZN(n1546) );
  XNOR2_X1 U2005 ( .A(b[7]), .B(n2269), .ZN(n1573) );
  XNOR2_X1 U2006 ( .A(b[3]), .B(n1997), .ZN(n1502) );
  XNOR2_X1 U2007 ( .A(b[5]), .B(n1996), .ZN(n1500) );
  XNOR2_X1 U2008 ( .A(b[7]), .B(n1995), .ZN(n1498) );
  XNOR2_X1 U2009 ( .A(b[5]), .B(n2269), .ZN(n1575) );
  XNOR2_X1 U2010 ( .A(b[5]), .B(n1981), .ZN(n1550) );
  XNOR2_X1 U2011 ( .A(b[9]), .B(n2043), .ZN(n1621) );
  XNOR2_X1 U2012 ( .A(b[9]), .B(n1996), .ZN(n1496) );
  XNOR2_X1 U2013 ( .A(b[3]), .B(n1981), .ZN(n1552) );
  XNOR2_X1 U2014 ( .A(b[1]), .B(n1981), .ZN(n1554) );
  XNOR2_X1 U2015 ( .A(b[7]), .B(n2043), .ZN(n1623) );
  XNOR2_X1 U2016 ( .A(b[9]), .B(n1954), .ZN(n1646) );
  XNOR2_X1 U2017 ( .A(b[3]), .B(n2269), .ZN(n1577) );
  XNOR2_X1 U2018 ( .A(b[3]), .B(n2043), .ZN(n1627) );
  XNOR2_X1 U2019 ( .A(b[7]), .B(n2288), .ZN(n1673) );
  XNOR2_X1 U2020 ( .A(b[1]), .B(n2002), .ZN(n1679) );
  XNOR2_X1 U2021 ( .A(b[5]), .B(n2289), .ZN(n1675) );
  XNOR2_X1 U2022 ( .A(b[5]), .B(n2304), .ZN(n1750) );
  XNOR2_X1 U2023 ( .A(b[3]), .B(n2289), .ZN(n1677) );
  XNOR2_X1 U2024 ( .A(b[7]), .B(n2025), .ZN(n1748) );
  XNOR2_X1 U2025 ( .A(b[1]), .B(n2269), .ZN(n1579) );
  XNOR2_X1 U2026 ( .A(b[9]), .B(n2288), .ZN(n1671) );
  XNOR2_X1 U2027 ( .A(b[1]), .B(n2304), .ZN(n1754) );
  XNOR2_X1 U2028 ( .A(b[1]), .B(n1999), .ZN(n1629) );
  XNOR2_X1 U2029 ( .A(b[3]), .B(n2025), .ZN(n1752) );
  XNOR2_X1 U2030 ( .A(b[7]), .B(n1954), .ZN(n1648) );
  XNOR2_X1 U2031 ( .A(b[5]), .B(n2043), .ZN(n1625) );
  XNOR2_X1 U2032 ( .A(b[9]), .B(n2025), .ZN(n1746) );
  XNOR2_X1 U2033 ( .A(b[1]), .B(n1954), .ZN(n1654) );
  XNOR2_X1 U2034 ( .A(b[15]), .B(n1997), .ZN(n1490) );
  XNOR2_X1 U2035 ( .A(b[17]), .B(n1996), .ZN(n1488) );
  XNOR2_X1 U2036 ( .A(b[13]), .B(n1997), .ZN(n1492) );
  XNOR2_X1 U2037 ( .A(b[11]), .B(n1997), .ZN(n1494) );
  XNOR2_X1 U2038 ( .A(b[19]), .B(n1996), .ZN(n1486) );
  XNOR2_X1 U2039 ( .A(b[21]), .B(n1997), .ZN(n1484) );
  XNOR2_X1 U2040 ( .A(a[2]), .B(n2303), .ZN(n2142) );
  XNOR2_X1 U2041 ( .A(a[4]), .B(n2298), .ZN(n2144) );
  INV_X1 U2042 ( .A(a[23]), .ZN(n2261) );
  XOR2_X1 U2043 ( .A(a[8]), .B(n2286), .Z(n1813) );
  OAI21_X1 U2044 ( .B1(a[0]), .B2(n2033), .A(n2313), .ZN(n1458) );
  INV_X1 U2045 ( .A(n1757), .ZN(n2313) );
  INV_X1 U2046 ( .A(a[0]), .ZN(n251) );
  XNOR2_X1 U2047 ( .A(b[23]), .B(n1996), .ZN(n1482) );
  INV_X1 U2048 ( .A(n2020), .ZN(n523) );
  NAND2_X1 U2049 ( .A1(n2020), .A2(n2180), .ZN(n516) );
  OAI21_X1 U2050 ( .B1(n2131), .B2(n2018), .A(n2322), .ZN(n1242) );
  INV_X1 U2051 ( .A(n2285), .ZN(n2282) );
  INV_X1 U2052 ( .A(n2145), .ZN(n2228) );
  BUF_X2 U2053 ( .A(n2069), .Z(n2157) );
  NOR2_X1 U2054 ( .A1(n919), .A2(n940), .ZN(n2158) );
  INV_X1 U2055 ( .A(n2131), .ZN(n2159) );
  OAI21_X1 U2056 ( .B1(n2140), .B2(n2191), .A(n2319), .ZN(n1314) );
  INV_X1 U2057 ( .A(n2137), .ZN(n2254) );
  NAND2_X1 U2058 ( .A1(n906), .A2(n893), .ZN(n2161) );
  NAND2_X1 U2059 ( .A1(n906), .A2(n889), .ZN(n2162) );
  NAND2_X1 U2060 ( .A1(n893), .A2(n889), .ZN(n2163) );
  NAND3_X1 U2061 ( .A1(n2161), .A2(n2162), .A3(n2163), .ZN(n882) );
  NAND2_X1 U2062 ( .A1(n1041), .A2(n1056), .ZN(n2164) );
  NAND2_X1 U2063 ( .A1(n1041), .A2(n1043), .ZN(n2165) );
  NAND2_X1 U2064 ( .A1(n1056), .A2(n1043), .ZN(n2166) );
  NAND3_X1 U2065 ( .A1(n2164), .A2(n2165), .A3(n2166), .ZN(n1038) );
  NOR2_X1 U2066 ( .A1(n1978), .A2(n2312), .ZN(n1385) );
  NOR2_X1 U2067 ( .A1(n2253), .A2(n2312), .ZN(n1433) );
  NOR2_X1 U2068 ( .A1(n2251), .A2(n2312), .ZN(n1409) );
  NOR2_X1 U2069 ( .A1(n2243), .A2(n2312), .ZN(n1265) );
  NOR2_X1 U2070 ( .A1(n2150), .A2(n2312), .ZN(n1313) );
  NOR2_X1 U2071 ( .A1(n2241), .A2(n2312), .ZN(n1241) );
  NOR2_X1 U2072 ( .A1(n2036), .A2(n2312), .ZN(n1361) );
  NOR2_X1 U2073 ( .A1(n2248), .A2(n2312), .ZN(n1337) );
  NOR2_X1 U2074 ( .A1(n2246), .A2(n2312), .ZN(n1289) );
  NAND2_X1 U2075 ( .A1(n2299), .A2(n2312), .ZN(n1731) );
  NAND2_X1 U2076 ( .A1(n2025), .A2(n2312), .ZN(n1756) );
  NOR2_X1 U2077 ( .A1(n2255), .A2(n2312), .ZN(n1457) );
  NAND2_X1 U2078 ( .A1(n2308), .A2(n2312), .ZN(n1781) );
  NAND2_X1 U2079 ( .A1(n2280), .A2(n2312), .ZN(n1631) );
  NAND2_X1 U2080 ( .A1(n2270), .A2(n2312), .ZN(n1581) );
  NAND2_X1 U2081 ( .A1(n2287), .A2(n2312), .ZN(n1681) );
  NAND2_X1 U2082 ( .A1(n2263), .A2(n2312), .ZN(n1531) );
  XNOR2_X1 U2083 ( .A(n2043), .B(n1998), .ZN(n1630) );
  NAND2_X1 U2084 ( .A1(n2293), .A2(n2312), .ZN(n1706) );
  XNOR2_X1 U2085 ( .A(n2309), .B(n1998), .ZN(n1780) );
  NAND2_X1 U2086 ( .A1(n2265), .A2(n2312), .ZN(n1556) );
  XNOR2_X1 U2087 ( .A(n2300), .B(n1998), .ZN(n1730) );
  XNOR2_X1 U2088 ( .A(n2294), .B(n1998), .ZN(n1705) );
  XNOR2_X1 U2089 ( .A(n2283), .B(n1998), .ZN(n1655) );
  NAND2_X1 U2090 ( .A1(n2003), .A2(n2312), .ZN(n1656) );
  NAND2_X1 U2091 ( .A1(n2276), .A2(n2312), .ZN(n1606) );
  XNOR2_X1 U2092 ( .A(n2271), .B(n1998), .ZN(n1580) );
  XNOR2_X1 U2093 ( .A(n2289), .B(n1998), .ZN(n1680) );
  XNOR2_X1 U2094 ( .A(n2025), .B(n1998), .ZN(n1755) );
  XNOR2_X1 U2095 ( .A(n2266), .B(n1998), .ZN(n1555) );
  XNOR2_X1 U2096 ( .A(n2275), .B(n1998), .ZN(n1605) );
  XNOR2_X1 U2097 ( .A(n2262), .B(n1998), .ZN(n1530) );
  INV_X1 U2098 ( .A(n383), .ZN(n381) );
  OR2_X2 U2099 ( .A1(n749), .A2(n760), .ZN(n2167) );
  NAND2_X1 U2100 ( .A1(n674), .A2(n550), .ZN(n323) );
  OR2_X1 U2101 ( .A1(n1021), .A2(n1038), .ZN(n2169) );
  AND2_X1 U2102 ( .A1(n1806), .A2(n1963), .ZN(n2170) );
  NAND2_X1 U2103 ( .A1(n859), .A2(n878), .ZN(n2171) );
  NAND2_X1 U2104 ( .A1(n859), .A2(n861), .ZN(n2172) );
  NAND2_X1 U2105 ( .A1(n878), .A2(n861), .ZN(n2173) );
  NAND3_X1 U2106 ( .A1(n2171), .A2(n2172), .A3(n2173), .ZN(n856) );
  XNOR2_X1 U2107 ( .A(n2174), .B(n1413), .ZN(n933) );
  XNOR2_X1 U2108 ( .A(n1435), .B(n1325), .ZN(n2174) );
  XNOR2_X1 U2109 ( .A(b[23]), .B(n1977), .ZN(n1507) );
  XNOR2_X1 U2110 ( .A(b[9]), .B(n1977), .ZN(n1521) );
  XNOR2_X1 U2111 ( .A(b[5]), .B(n1977), .ZN(n1525) );
  XNOR2_X1 U2112 ( .A(b[7]), .B(n1977), .ZN(n1523) );
  XNOR2_X1 U2113 ( .A(b[1]), .B(n2262), .ZN(n1529) );
  OAI21_X1 U2114 ( .B1(n2134), .B2(n2196), .A(n2320), .ZN(n1290) );
  XNOR2_X1 U2115 ( .A(b[1]), .B(n2297), .ZN(n1729) );
  XNOR2_X1 U2116 ( .A(b[9]), .B(n2297), .ZN(n1721) );
  XNOR2_X1 U2117 ( .A(b[3]), .B(n2297), .ZN(n1727) );
  XNOR2_X1 U2118 ( .A(b[5]), .B(n2297), .ZN(n1725) );
  XNOR2_X1 U2119 ( .A(b[7]), .B(n2297), .ZN(n1723) );
  XNOR2_X1 U2120 ( .A(b[23]), .B(n2297), .ZN(n1707) );
  XNOR2_X1 U2121 ( .A(n2260), .B(b[22]), .ZN(n1483) );
  XNOR2_X1 U2122 ( .A(n2260), .B(b[18]), .ZN(n1487) );
  XNOR2_X1 U2123 ( .A(n1939), .B(b[20]), .ZN(n1485) );
  XNOR2_X1 U2124 ( .A(n1939), .B(b[10]), .ZN(n1495) );
  XNOR2_X1 U2125 ( .A(n1939), .B(b[16]), .ZN(n1489) );
  XNOR2_X1 U2126 ( .A(n2260), .B(b[12]), .ZN(n1493) );
  XNOR2_X1 U2127 ( .A(n2260), .B(b[6]), .ZN(n1499) );
  XNOR2_X1 U2128 ( .A(n1939), .B(b[4]), .ZN(n1501) );
  XNOR2_X1 U2129 ( .A(n2260), .B(b[14]), .ZN(n1491) );
  XNOR2_X1 U2130 ( .A(n1939), .B(n1998), .ZN(n1505) );
  XNOR2_X1 U2131 ( .A(n2260), .B(b[8]), .ZN(n1497) );
  XNOR2_X1 U2132 ( .A(n2260), .B(b[2]), .ZN(n1503) );
  INV_X2 U2133 ( .A(n1938), .ZN(n2260) );
  XNOR2_X1 U2134 ( .A(b[23]), .B(n2277), .ZN(n1582) );
  XNOR2_X1 U2135 ( .A(b[3]), .B(n2274), .ZN(n1602) );
  XNOR2_X1 U2136 ( .A(b[5]), .B(n2274), .ZN(n1600) );
  XNOR2_X1 U2137 ( .A(b[9]), .B(n2276), .ZN(n1596) );
  XNOR2_X1 U2138 ( .A(b[7]), .B(n2275), .ZN(n1598) );
  XNOR2_X1 U2139 ( .A(b[1]), .B(n2276), .ZN(n1604) );
  NAND2_X1 U2140 ( .A1(n1413), .A2(n1435), .ZN(n2175) );
  NAND2_X1 U2141 ( .A1(n1413), .A2(n1325), .ZN(n2176) );
  NAND2_X1 U2142 ( .A1(n1435), .A2(n1325), .ZN(n2177) );
  NAND3_X1 U2143 ( .A1(n2175), .A2(n2176), .A3(n2177), .ZN(n932) );
  OR2_X1 U2144 ( .A1(n2149), .A2(n1711), .ZN(n2178) );
  OR2_X1 U2145 ( .A1(n2254), .A2(n1710), .ZN(n2179) );
  NAND2_X1 U2146 ( .A1(n2178), .A2(n2179), .ZN(n1413) );
  XNOR2_X1 U2147 ( .A(n2300), .B(b[20]), .ZN(n1710) );
  NAND2_X1 U2148 ( .A1(n941), .A2(n962), .ZN(n550) );
  OAI21_X1 U2149 ( .B1(n2135), .B2(n1986), .A(n2316), .ZN(n1386) );
  OR2_X1 U2150 ( .A1(n857), .A2(n876), .ZN(n2180) );
  INV_X1 U2151 ( .A(n2290), .ZN(n2286) );
  AOI21_X1 U2152 ( .B1(n625), .B2(n1971), .A(n1962), .ZN(n620) );
  OAI22_X1 U2153 ( .A1(n1988), .A2(n1772), .B1(n1771), .B2(n2258), .ZN(n1473)
         );
  OAI22_X1 U2154 ( .A1(n2236), .A2(n1777), .B1(n1776), .B2(n2257), .ZN(n1478)
         );
  OAI22_X1 U2155 ( .A1(n1988), .A2(n1769), .B1(n1768), .B2(n2257), .ZN(n1470)
         );
  OAI22_X1 U2156 ( .A1(n1988), .A2(n1780), .B1(n1779), .B2(n2258), .ZN(n1481)
         );
  OAI22_X1 U2157 ( .A1(n1988), .A2(n1773), .B1(n1772), .B2(n2258), .ZN(n1474)
         );
  OAI22_X1 U2158 ( .A1(n1988), .A2(n1776), .B1(n1775), .B2(n2258), .ZN(n1477)
         );
  OAI22_X1 U2159 ( .A1(n2236), .A2(n1779), .B1(n1778), .B2(n2257), .ZN(n1480)
         );
  OAI22_X1 U2160 ( .A1(n2236), .A2(n1775), .B1(n1774), .B2(n2257), .ZN(n1476)
         );
  OAI22_X1 U2161 ( .A1(n2236), .A2(n1771), .B1(n1770), .B2(n2258), .ZN(n1472)
         );
  OAI22_X1 U2162 ( .A1(n2236), .A2(n1778), .B1(n1777), .B2(n2257), .ZN(n1479)
         );
  OAI22_X1 U2163 ( .A1(n1988), .A2(n1770), .B1(n1769), .B2(n2258), .ZN(n1471)
         );
  OAI22_X1 U2164 ( .A1(n1988), .A2(n1774), .B1(n1773), .B2(n2257), .ZN(n1475)
         );
  OAI21_X1 U2165 ( .B1(n2233), .B2(n2109), .A(n2318), .ZN(n1338) );
  NOR2_X1 U2166 ( .A1(n420), .A2(n402), .ZN(n400) );
  OAI22_X1 U2167 ( .A1(n2100), .A2(n1696), .B1(n2251), .B2(n1695), .ZN(n1399)
         );
  XNOR2_X1 U2168 ( .A(b[5]), .B(n2292), .ZN(n1700) );
  XNOR2_X1 U2169 ( .A(b[1]), .B(n2292), .ZN(n1704) );
  XNOR2_X1 U2170 ( .A(b[7]), .B(n2292), .ZN(n1698) );
  XNOR2_X1 U2171 ( .A(b[3]), .B(n2292), .ZN(n1702) );
  XNOR2_X1 U2172 ( .A(b[9]), .B(n2292), .ZN(n1696) );
  XNOR2_X1 U2173 ( .A(b[23]), .B(n2292), .ZN(n1682) );
  NOR2_X1 U2174 ( .A1(n502), .A2(n495), .ZN(n489) );
  INV_X1 U2175 ( .A(n2295), .ZN(n2291) );
  AND2_X1 U2176 ( .A1(n2020), .A2(n1991), .ZN(n2182) );
  INV_X1 U2177 ( .A(n2311), .ZN(n2184) );
  INV_X1 U2178 ( .A(n2311), .ZN(n2183) );
  XNOR2_X1 U2179 ( .A(b[11]), .B(n2002), .ZN(n1669) );
  OR2_X1 U2180 ( .A1(n856), .A2(n2073), .ZN(n2185) );
  INV_X1 U2181 ( .A(n2008), .ZN(n2188) );
  NOR2_X1 U2182 ( .A1(n839), .A2(n856), .ZN(n513) );
  OR2_X1 U2183 ( .A1(n502), .A2(n2059), .ZN(n2186) );
  NOR2_X1 U2184 ( .A1(n821), .A2(n838), .ZN(n502) );
  INV_X1 U2185 ( .A(n674), .ZN(n2187) );
  INV_X1 U2186 ( .A(n2009), .ZN(n2189) );
  NOR2_X1 U2187 ( .A1(n941), .A2(n962), .ZN(n547) );
  NAND2_X1 U2188 ( .A1(n1939), .A2(n2312), .ZN(n1506) );
  OR2_X2 U2189 ( .A1(n788), .A2(n775), .ZN(n2190) );
  OAI21_X1 U2190 ( .B1(n2009), .B2(n2181), .A(n2317), .ZN(n1362) );
  INV_X1 U2191 ( .A(n1934), .ZN(n2274) );
  BUF_X2 U2192 ( .A(n285), .Z(n2193) );
  INV_X1 U2193 ( .A(n2138), .ZN(n2223) );
  INV_X1 U2194 ( .A(n802), .ZN(n803) );
  INV_X1 U2195 ( .A(n2140), .ZN(n2231) );
  OAI21_X1 U2196 ( .B1(n390), .B2(n384), .A(n387), .ZN(n383) );
  AOI21_X1 U2197 ( .B1(n401), .B2(n2120), .A(n394), .ZN(n390) );
  XNOR2_X1 U2198 ( .A(b[11]), .B(n2297), .ZN(n1719) );
  NOR2_X1 U2199 ( .A1(n919), .A2(n940), .ZN(n542) );
  CLKBUF_X1 U2200 ( .A(n505), .Z(n2194) );
  OR2_X1 U2201 ( .A1(n940), .A2(n1929), .ZN(n2195) );
  INV_X1 U2202 ( .A(n2281), .ZN(n2279) );
  INV_X1 U2203 ( .A(n2273), .ZN(n2268) );
  NAND2_X1 U2204 ( .A1(n588), .A2(n2115), .ZN(n582) );
  OAI22_X1 U2205 ( .A1(n2041), .A2(n1701), .B1(n1700), .B2(n2251), .ZN(n1404)
         );
  OAI22_X1 U2206 ( .A1(n2053), .A2(n1695), .B1(n1694), .B2(n2251), .ZN(n1398)
         );
  OAI22_X1 U2207 ( .A1(n2074), .A2(n1704), .B1(n2252), .B2(n1703), .ZN(n1407)
         );
  OAI22_X1 U2208 ( .A1(n2074), .A2(n1700), .B1(n2252), .B2(n1699), .ZN(n1403)
         );
  OAI22_X1 U2209 ( .A1(n2100), .A2(n1699), .B1(n1698), .B2(n2251), .ZN(n1402)
         );
  OAI22_X1 U2210 ( .A1(n2074), .A2(n1694), .B1(n2251), .B2(n1693), .ZN(n1397)
         );
  OAI22_X1 U2211 ( .A1(n2074), .A2(n1702), .B1(n2251), .B2(n1701), .ZN(n1405)
         );
  OAI22_X1 U2212 ( .A1(n2074), .A2(n1698), .B1(n2252), .B2(n1697), .ZN(n1401)
         );
  INV_X1 U2213 ( .A(n2055), .ZN(n555) );
  NOR2_X1 U2214 ( .A1(n563), .A2(n558), .ZN(n552) );
  OAI21_X1 U2215 ( .B1(n558), .B2(n564), .A(n559), .ZN(n553) );
  OAI22_X1 U2216 ( .A1(n2236), .A2(n2311), .B1(n1781), .B2(n2257), .ZN(n1193)
         );
  OAI22_X1 U2217 ( .A1(n2236), .A2(n1768), .B1(n1767), .B2(n2257), .ZN(n1469)
         );
  OAI22_X1 U2218 ( .A1(n2236), .A2(n1764), .B1(n1763), .B2(n2258), .ZN(n1465)
         );
  OAI22_X1 U2219 ( .A1(n2236), .A2(n1760), .B1(n1759), .B2(n2257), .ZN(n1461)
         );
  OAI22_X1 U2220 ( .A1(n2236), .A2(n1763), .B1(n1762), .B2(n2257), .ZN(n1464)
         );
  OAI22_X1 U2221 ( .A1(n2236), .A2(n1767), .B1(n1766), .B2(n2258), .ZN(n1468)
         );
  OAI22_X1 U2222 ( .A1(n2237), .A2(n1759), .B1(n1758), .B2(n2258), .ZN(n1460)
         );
  OAI22_X1 U2223 ( .A1(n2237), .A2(n1761), .B1(n1760), .B2(n2258), .ZN(n1462)
         );
  OAI22_X1 U2224 ( .A1(n2237), .A2(n1758), .B1(n1757), .B2(n2257), .ZN(n1459)
         );
  OAI22_X1 U2225 ( .A1(n1988), .A2(n1765), .B1(n1764), .B2(n2258), .ZN(n1466)
         );
  OAI22_X1 U2226 ( .A1(n1988), .A2(n1766), .B1(n1765), .B2(n2258), .ZN(n1467)
         );
  OAI22_X1 U2227 ( .A1(n2237), .A2(n1762), .B1(n1761), .B2(n2257), .ZN(n1463)
         );
  XNOR2_X1 U2228 ( .A(b[1]), .B(n2309), .ZN(n1779) );
  XNOR2_X1 U2229 ( .A(b[5]), .B(n2183), .ZN(n1775) );
  XNOR2_X1 U2230 ( .A(b[9]), .B(n2183), .ZN(n1771) );
  XNOR2_X1 U2231 ( .A(b[7]), .B(n2309), .ZN(n1773) );
  XNOR2_X1 U2232 ( .A(b[3]), .B(n2183), .ZN(n1777) );
  XNOR2_X1 U2233 ( .A(b[23]), .B(n2183), .ZN(n1757) );
  OAI22_X1 U2234 ( .A1(n1985), .A2(n1536), .B1(n2243), .B2(n1535), .ZN(n1245)
         );
  OAI22_X1 U2235 ( .A1(n1985), .A2(n1534), .B1(n2244), .B2(n1533), .ZN(n1243)
         );
  OAI22_X1 U2236 ( .A1(n2226), .A2(n1542), .B1(n2244), .B2(n1541), .ZN(n1251)
         );
  OAI22_X1 U2237 ( .A1(n2159), .A2(n1540), .B1(n2243), .B2(n1539), .ZN(n1249)
         );
  OAI21_X1 U2238 ( .B1(n2034), .B2(n1992), .A(n2323), .ZN(n1218) );
  INV_X1 U2239 ( .A(n502), .ZN(n668) );
  XNOR2_X1 U2240 ( .A(n2198), .B(n2083), .ZN(n953) );
  XNOR2_X1 U2241 ( .A(n1326), .B(n1392), .ZN(n2198) );
  NAND2_X1 U2242 ( .A1(n668), .A2(n2035), .ZN(n317) );
  INV_X1 U2243 ( .A(n503), .ZN(n501) );
  AOI21_X1 U2244 ( .B1(n359), .B2(n2126), .A(n350), .ZN(n348) );
  INV_X1 U2245 ( .A(n2131), .ZN(n2225) );
  AOI21_X1 U2246 ( .B1(n589), .B2(n2115), .A(n1969), .ZN(n583) );
  NAND2_X1 U2247 ( .A1(n1326), .A2(n1392), .ZN(n2199) );
  NAND2_X1 U2248 ( .A1(n1326), .A2(n961), .ZN(n2200) );
  NAND2_X1 U2249 ( .A1(n1392), .A2(n961), .ZN(n2201) );
  NAND3_X1 U2250 ( .A1(n2199), .A2(n2200), .A3(n2201), .ZN(n952) );
  NAND2_X1 U2251 ( .A1(n2040), .A2(n959), .ZN(n2202) );
  NAND2_X1 U2252 ( .A1(n972), .A2(n953), .ZN(n2203) );
  NAND2_X1 U2253 ( .A1(n959), .A2(n953), .ZN(n2204) );
  NAND3_X1 U2254 ( .A1(n2202), .A2(n2203), .A3(n2204), .ZN(n946) );
  OR2_X1 U2255 ( .A1(n2223), .A2(n1528), .ZN(n2205) );
  OR2_X1 U2256 ( .A1(n1527), .A2(n2240), .ZN(n2206) );
  NAND2_X1 U2257 ( .A1(n2205), .A2(n2206), .ZN(n1238) );
  XNOR2_X1 U2258 ( .A(n2262), .B(b[2]), .ZN(n1528) );
  XNOR2_X1 U2259 ( .A(b[3]), .B(n2262), .ZN(n1527) );
  CLKBUF_X1 U2260 ( .A(n2209), .Z(n2207) );
  OAI21_X1 U2261 ( .B1(n2145), .B2(n1989), .A(n2321), .ZN(n1266) );
  NOR2_X1 U2262 ( .A1(n983), .A2(n1002), .ZN(n563) );
  NAND2_X1 U2263 ( .A1(n983), .A2(n1002), .ZN(n564) );
  NAND2_X1 U2264 ( .A1(n2113), .A2(n461), .ZN(n313) );
  INV_X1 U2265 ( .A(n461), .ZN(n459) );
  NAND2_X1 U2266 ( .A1(n1003), .A2(n1020), .ZN(n570) );
  NOR2_X1 U2267 ( .A1(n1003), .A2(n1020), .ZN(n569) );
  INV_X1 U2268 ( .A(n2306), .ZN(n2303) );
  AOI21_X1 U2269 ( .B1(n511), .B2(n526), .A(n512), .ZN(n2209) );
  NAND2_X1 U2270 ( .A1(n1812), .A2(n1964), .ZN(n285) );
  INV_X1 U2271 ( .A(n285), .ZN(n2233) );
  INV_X1 U2272 ( .A(n547), .ZN(n674) );
  NOR2_X1 U2273 ( .A1(n554), .A2(n2187), .ZN(n545) );
  OAI21_X1 U2274 ( .B1(n555), .B2(n2187), .A(n550), .ZN(n546) );
  NAND2_X1 U2275 ( .A1(n919), .A2(n940), .ZN(n543) );
  NAND2_X1 U2276 ( .A1(n1932), .A2(n2114), .ZN(n571) );
  AOI21_X1 U2277 ( .B1(n2169), .B2(n2112), .A(n1970), .ZN(n572) );
  INV_X1 U2278 ( .A(n401), .ZN(n399) );
  OAI21_X1 U2279 ( .B1(n421), .B2(n402), .A(n405), .ZN(n401) );
  AOI21_X1 U2280 ( .B1(n595), .B2(n609), .A(n596), .ZN(n594) );
  OAI21_X1 U2281 ( .B1(n620), .B2(n610), .A(n611), .ZN(n609) );
  INV_X1 U2282 ( .A(n2137), .ZN(n2253) );
  OAI21_X1 U2283 ( .B1(n2143), .B2(n2137), .A(n2315), .ZN(n1410) );
  AOI21_X1 U2284 ( .B1(n511), .B2(n2019), .A(n512), .ZN(n506) );
  XNOR2_X1 U2285 ( .A(b[21]), .B(n1981), .ZN(n1534) );
  XNOR2_X1 U2286 ( .A(b[19]), .B(n1981), .ZN(n1536) );
  XNOR2_X1 U2287 ( .A(b[13]), .B(n1981), .ZN(n1542) );
  XNOR2_X1 U2288 ( .A(b[11]), .B(n1981), .ZN(n1544) );
  XNOR2_X1 U2289 ( .A(b[15]), .B(n1981), .ZN(n1540) );
  XNOR2_X1 U2290 ( .A(b[17]), .B(n1981), .ZN(n1538) );
  OAI21_X1 U2291 ( .B1(n456), .B2(n481), .A(n457), .ZN(n455) );
  AOI21_X1 U2292 ( .B1(n565), .B2(n1979), .A(n2055), .ZN(n551) );
  INV_X1 U2293 ( .A(n552), .ZN(n554) );
  NOR2_X1 U2294 ( .A1(n597), .A2(n599), .ZN(n595) );
  OAI21_X1 U2295 ( .B1(n600), .B2(n597), .A(n598), .ZN(n596) );
  NAND2_X1 U2296 ( .A1(n1099), .A2(n1110), .ZN(n598) );
  NOR2_X1 U2297 ( .A1(n1099), .A2(n1110), .ZN(n597) );
  NAND2_X1 U2298 ( .A1(n2180), .A2(n521), .ZN(n319) );
  INV_X1 U2299 ( .A(n521), .ZN(n519) );
  OAI21_X1 U2300 ( .B1(n2170), .B2(n2010), .A(n2324), .ZN(n1194) );
  NOR2_X1 U2301 ( .A1(n857), .A2(n876), .ZN(n520) );
  NAND2_X1 U2302 ( .A1(n857), .A2(n876), .ZN(n521) );
  INV_X1 U2303 ( .A(n2071), .ZN(n492) );
  XNOR2_X1 U2304 ( .A(b[17]), .B(n2025), .ZN(n1738) );
  XNOR2_X1 U2305 ( .A(n533), .B(n320), .ZN(product[26]) );
  NOR2_X1 U2306 ( .A1(n1085), .A2(n1098), .ZN(n592) );
  NAND2_X1 U2307 ( .A1(n701), .A2(n708), .ZN(n396) );
  XNOR2_X1 U2308 ( .A(b[19]), .B(n2279), .ZN(n1611) );
  XNOR2_X1 U2309 ( .A(b[21]), .B(n2279), .ZN(n1609) );
  XNOR2_X1 U2310 ( .A(b[11]), .B(n2279), .ZN(n1619) );
  XNOR2_X1 U2311 ( .A(b[13]), .B(n2279), .ZN(n1617) );
  XNOR2_X1 U2312 ( .A(b[17]), .B(n2279), .ZN(n1613) );
  XNOR2_X1 U2313 ( .A(b[15]), .B(n2279), .ZN(n1615) );
  INV_X1 U2314 ( .A(n400), .ZN(n398) );
  NAND2_X1 U2315 ( .A1(n400), .A2(n2120), .ZN(n389) );
  NAND2_X1 U2316 ( .A1(n426), .A2(n2167), .ZN(n420) );
  XNOR2_X1 U2317 ( .A(n522), .B(n319), .ZN(product[27]) );
  NAND2_X1 U2318 ( .A1(n2122), .A2(n2124), .ZN(n599) );
  XNOR2_X1 U2319 ( .A(n515), .B(n318), .ZN(product[28]) );
  NOR2_X1 U2320 ( .A1(n590), .A2(n592), .ZN(n588) );
  XNOR2_X1 U2321 ( .A(n504), .B(n317), .ZN(product[29]) );
  NAND2_X1 U2322 ( .A1(n332), .A2(n2128), .ZN(n326) );
  AOI21_X1 U2323 ( .B1(n2113), .B2(n472), .A(n459), .ZN(n457) );
  OAI22_X1 U2324 ( .A1(n2074), .A2(n1705), .B1(n1704), .B2(n2251), .ZN(n1408)
         );
  OAI22_X1 U2325 ( .A1(n2100), .A2(n1703), .B1(n1702), .B2(n2251), .ZN(n1406)
         );
  XNOR2_X1 U2326 ( .A(n486), .B(n315), .ZN(product[31]) );
  NAND2_X1 U2327 ( .A1(n1991), .A2(n525), .ZN(n505) );
  INV_X1 U2328 ( .A(n2008), .ZN(n2235) );
  OAI22_X1 U2329 ( .A1(n2188), .A2(n1671), .B1(n2250), .B2(n1670), .ZN(n1375)
         );
  OAI22_X1 U2330 ( .A1(n2188), .A2(n1672), .B1(n1671), .B2(n2250), .ZN(n1376)
         );
  OAI22_X1 U2331 ( .A1(n2234), .A2(n1676), .B1(n1675), .B2(n2250), .ZN(n1380)
         );
  OAI22_X1 U2332 ( .A1(n2234), .A2(n1669), .B1(n2250), .B2(n1668), .ZN(n1373)
         );
  OAI22_X1 U2333 ( .A1(n2188), .A2(n1679), .B1(n1978), .B2(n1678), .ZN(n1383)
         );
  OAI22_X1 U2334 ( .A1(n2234), .A2(n1670), .B1(n1669), .B2(n2250), .ZN(n1374)
         );
  NOR2_X1 U2335 ( .A1(n336), .A2(n334), .ZN(n332) );
  NAND2_X1 U2336 ( .A1(n356), .A2(n2126), .ZN(n347) );
  XOR2_X1 U2337 ( .A(n994), .B(n1217), .Z(n2210) );
  XOR2_X1 U2338 ( .A(n2026), .B(n2210), .Z(n973) );
  NAND2_X1 U2339 ( .A1(n2026), .A2(n994), .ZN(n2211) );
  NAND2_X1 U2340 ( .A1(n996), .A2(n1217), .ZN(n2212) );
  NAND2_X1 U2341 ( .A1(n994), .A2(n1217), .ZN(n2213) );
  NAND3_X1 U2342 ( .A1(n2211), .A2(n2212), .A3(n2213), .ZN(n972) );
  AND2_X1 U2343 ( .A1(n2219), .A2(n2220), .ZN(n2214) );
  OR2_X1 U2344 ( .A1(n2235), .A2(n1668), .ZN(n2216) );
  OR2_X1 U2345 ( .A1(n1667), .A2(n1978), .ZN(n2217) );
  NAND2_X1 U2346 ( .A1(n2216), .A2(n2217), .ZN(n1372) );
  OR2_X1 U2347 ( .A1(n897), .A2(n918), .ZN(n2218) );
  NOR2_X1 U2348 ( .A1(n2238), .A2(n2312), .ZN(n1217) );
  AND2_X1 U2349 ( .A1(n2219), .A2(n2220), .ZN(n301) );
  XNOR2_X1 U2350 ( .A(n2287), .B(b[12]), .ZN(n1668) );
  NOR2_X1 U2351 ( .A1(n571), .A2(n569), .ZN(n567) );
  INV_X1 U2352 ( .A(n2170), .ZN(n2222) );
  NAND2_X1 U2353 ( .A1(n2118), .A2(n418), .ZN(n309) );
  AOI21_X1 U2354 ( .B1(n333), .B2(n2128), .A(n2129), .ZN(n327) );
  OAI21_X1 U2355 ( .B1(n337), .B2(n334), .A(n335), .ZN(n333) );
  INV_X1 U2356 ( .A(n418), .ZN(n416) );
  NAND2_X1 U2357 ( .A1(n963), .A2(n982), .ZN(n559) );
  NAND2_X1 U2358 ( .A1(n666), .A2(n2190), .ZN(n467) );
  AOI21_X1 U2359 ( .B1(n2190), .B2(n483), .A(n472), .ZN(n468) );
  NAND2_X1 U2360 ( .A1(n2190), .A2(n2113), .ZN(n456) );
  NAND2_X1 U2361 ( .A1(n2218), .A2(n535), .ZN(n321) );
  INV_X1 U2362 ( .A(n526), .ZN(n524) );
  AOI21_X1 U2363 ( .B1(n526), .B2(n2180), .A(n519), .ZN(n517) );
  INV_X1 U2364 ( .A(n537), .ZN(n536) );
  NAND2_X1 U2365 ( .A1(n897), .A2(n918), .ZN(n535) );
  NAND2_X1 U2366 ( .A1(n2123), .A2(n378), .ZN(n305) );
  NAND2_X1 U2367 ( .A1(n382), .A2(n2123), .ZN(n371) );
  AOI21_X1 U2368 ( .B1(n383), .B2(n2123), .A(n376), .ZN(n372) );
  NAND2_X1 U2369 ( .A1(n2123), .A2(n2125), .ZN(n364) );
  NAND2_X1 U2370 ( .A1(n685), .A2(n688), .ZN(n369) );
  NOR2_X1 U2371 ( .A1(n542), .A2(n547), .ZN(n540) );
  OAI21_X1 U2372 ( .B1(n2158), .B2(n550), .A(n543), .ZN(n541) );
  XNOR2_X1 U2373 ( .A(b[21]), .B(n2268), .ZN(n1559) );
  XNOR2_X1 U2374 ( .A(b[19]), .B(n2268), .ZN(n1561) );
  XNOR2_X1 U2375 ( .A(b[15]), .B(n2268), .ZN(n1565) );
  XNOR2_X1 U2376 ( .A(b[17]), .B(n2268), .ZN(n1563) );
  XNOR2_X1 U2377 ( .A(b[11]), .B(n2268), .ZN(n1569) );
  XNOR2_X1 U2378 ( .A(b[13]), .B(n2268), .ZN(n1567) );
  NAND2_X1 U2379 ( .A1(n2190), .A2(n474), .ZN(n314) );
  INV_X1 U2380 ( .A(n474), .ZN(n472) );
  INV_X1 U2381 ( .A(n874), .ZN(n875) );
  INV_X1 U2382 ( .A(n2106), .ZN(n565) );
  AOI21_X1 U2383 ( .B1(n581), .B2(n567), .A(n568), .ZN(n566) );
  OAI21_X1 U2384 ( .B1(n572), .B2(n1948), .A(n570), .ZN(n568) );
  XNOR2_X1 U2385 ( .A(b[19]), .B(n2291), .ZN(n1686) );
  XNOR2_X1 U2386 ( .A(b[17]), .B(n2291), .ZN(n1688) );
  NOR2_X1 U2387 ( .A1(n918), .A2(n897), .ZN(n534) );
  NAND2_X1 U2388 ( .A1(n1171), .A2(n1174), .ZN(n634) );
  NOR2_X1 U2389 ( .A1(n1171), .A2(n1174), .ZN(n633) );
  OAI21_X1 U2390 ( .B1(n2052), .B2(n521), .A(n514), .ZN(n512) );
  NAND2_X1 U2391 ( .A1(n839), .A2(n856), .ZN(n514) );
  INV_X1 U2392 ( .A(n746), .ZN(n747) );
  NAND2_X1 U2393 ( .A1(n709), .A2(n716), .ZN(n409) );
  NOR2_X1 U2394 ( .A1(n2186), .A2(n480), .ZN(n478) );
  OAI21_X1 U2395 ( .B1(n492), .B2(n480), .A(n481), .ZN(n479) );
  INV_X1 U2396 ( .A(n480), .ZN(n666) );
  NOR2_X1 U2397 ( .A1(n456), .A2(n480), .ZN(n454) );
  NOR2_X2 U2398 ( .A1(n789), .A2(n804), .ZN(n480) );
  OAI21_X1 U2399 ( .B1(n594), .B2(n582), .A(n583), .ZN(n581) );
  XNOR2_X1 U2400 ( .A(n497), .B(n316), .ZN(product[30]) );
  AOI21_X1 U2401 ( .B1(n508), .B2(n465), .A(n466), .ZN(n464) );
  AOI21_X1 U2402 ( .B1(n508), .B2(n478), .A(n479), .ZN(n477) );
  AOI21_X1 U2403 ( .B1(n508), .B2(n668), .A(n501), .ZN(n499) );
  NAND2_X1 U2404 ( .A1(n1165), .A2(n1170), .ZN(n632) );
  OAI22_X1 U2405 ( .A1(n2189), .A2(n1678), .B1(n1677), .B2(n1978), .ZN(n1382)
         );
  OAI22_X1 U2406 ( .A1(n2235), .A2(n1674), .B1(n1673), .B2(n2250), .ZN(n1378)
         );
  OAI22_X1 U2407 ( .A1(n2189), .A2(n1680), .B1(n1679), .B2(n1978), .ZN(n1384)
         );
  OAI22_X1 U2408 ( .A1(n2189), .A2(n1673), .B1(n2250), .B2(n1672), .ZN(n1377)
         );
  OAI22_X1 U2409 ( .A1(n2234), .A2(n1675), .B1(n2250), .B2(n1674), .ZN(n1379)
         );
  OAI22_X1 U2410 ( .A1(n2188), .A2(n1677), .B1(n2250), .B2(n1676), .ZN(n1381)
         );
  INV_X1 U2411 ( .A(n2059), .ZN(n667) );
  OAI21_X1 U2412 ( .B1(n495), .B2(n503), .A(n496), .ZN(n490) );
  INV_X1 U2413 ( .A(n420), .ZN(n422) );
  NOR2_X1 U2414 ( .A1(n420), .A2(n347), .ZN(n345) );
  NAND2_X1 U2415 ( .A1(n749), .A2(n760), .ZN(n439) );
  OAI22_X1 U2416 ( .A1(n2100), .A2(n1697), .B1(n1696), .B2(n2251), .ZN(n1400)
         );
  INV_X1 U2417 ( .A(n2021), .ZN(n671) );
  INV_X1 U2418 ( .A(n2209), .ZN(n508) );
  INV_X1 U2419 ( .A(n428), .ZN(n661) );
  OAI21_X1 U2420 ( .B1(n428), .B2(n436), .A(n429), .ZN(n427) );
  NAND2_X1 U2421 ( .A1(n727), .A2(n736), .ZN(n429) );
  NOR2_X1 U2422 ( .A1(n727), .A2(n736), .ZN(n428) );
  OAI22_X1 U2423 ( .A1(n2056), .A2(n1613), .B1(n2157), .B2(n1612), .ZN(n1319)
         );
  OAI22_X1 U2424 ( .A1(n2057), .A2(n1615), .B1(n2248), .B2(n1614), .ZN(n1321)
         );
  OAI22_X1 U2425 ( .A1(n2232), .A2(n2281), .B1(n1631), .B2(n2157), .ZN(n1187)
         );
  OAI22_X1 U2426 ( .A1(n2056), .A2(n1612), .B1(n1611), .B2(n2157), .ZN(n1318)
         );
  OAI22_X1 U2427 ( .A1(n2232), .A2(n1617), .B1(n2248), .B2(n1616), .ZN(n1323)
         );
  OAI22_X1 U2428 ( .A1(n2232), .A2(n1614), .B1(n1613), .B2(n2157), .ZN(n1320)
         );
  OAI22_X1 U2429 ( .A1(n2057), .A2(n1611), .B1(n2248), .B2(n1610), .ZN(n1317)
         );
  OAI22_X1 U2430 ( .A1(n2231), .A2(n1618), .B1(n1617), .B2(n2157), .ZN(n1324)
         );
  OAI22_X1 U2431 ( .A1(n2056), .A2(n1608), .B1(n1607), .B2(n2157), .ZN(n746)
         );
  OAI22_X1 U2432 ( .A1(n2232), .A2(n1610), .B1(n1609), .B2(n2157), .ZN(n1316)
         );
  OAI22_X1 U2433 ( .A1(n2231), .A2(n1616), .B1(n1615), .B2(n2157), .ZN(n1322)
         );
  OAI22_X1 U2434 ( .A1(n2232), .A2(n1609), .B1(n2157), .B2(n1608), .ZN(n1315)
         );
  AOI21_X1 U2435 ( .B1(n508), .B2(n2031), .A(n2084), .ZN(n488) );
  NAND2_X1 U2436 ( .A1(n465), .A2(n2182), .ZN(n463) );
  NAND2_X1 U2437 ( .A1(n478), .A2(n2182), .ZN(n476) );
  NAND2_X1 U2438 ( .A1(n2182), .A2(n668), .ZN(n498) );
  NAND2_X1 U2439 ( .A1(n2182), .A2(n2031), .ZN(n487) );
  NAND2_X1 U2440 ( .A1(n877), .A2(n896), .ZN(n532) );
  NAND2_X1 U2441 ( .A1(n537), .A2(n450), .ZN(n2219) );
  INV_X1 U2442 ( .A(n451), .ZN(n2220) );
  OAI22_X1 U2443 ( .A1(n2100), .A2(n1683), .B1(n1682), .B2(n2251), .ZN(n2221)
         );
  NOR2_X1 U2444 ( .A1(n505), .A2(n452), .ZN(n450) );
  NAND2_X1 U2445 ( .A1(n694), .A2(n689), .ZN(n378) );
  XNOR2_X1 U2446 ( .A(n475), .B(n314), .ZN(product[32]) );
  NAND2_X1 U2447 ( .A1(n805), .A2(n820), .ZN(n496) );
  XNOR2_X1 U2448 ( .A(n437), .B(n311), .ZN(product[35]) );
  XNOR2_X1 U2449 ( .A(b[17]), .B(n2184), .ZN(n1763) );
  XNOR2_X1 U2450 ( .A(b[21]), .B(n2183), .ZN(n1759) );
  XNOR2_X1 U2451 ( .A(b[13]), .B(n2183), .ZN(n1767) );
  XNOR2_X1 U2452 ( .A(n430), .B(n310), .ZN(product[36]) );
  XNOR2_X1 U2453 ( .A(n419), .B(n309), .ZN(product[37]) );
  OAI22_X1 U2454 ( .A1(n2189), .A2(n1661), .B1(n1978), .B2(n1660), .ZN(n1365)
         );
  OAI22_X1 U2455 ( .A1(n2234), .A2(n1660), .B1(n1659), .B2(n1978), .ZN(n1364)
         );
  OAI22_X1 U2456 ( .A1(n2188), .A2(n1663), .B1(n1978), .B2(n1662), .ZN(n1367)
         );
  OAI22_X1 U2457 ( .A1(n2234), .A2(n1982), .B1(n1681), .B2(n1978), .ZN(n1189)
         );
  OAI22_X1 U2458 ( .A1(n2234), .A2(n1664), .B1(n1663), .B2(n1978), .ZN(n1368)
         );
  OAI22_X1 U2459 ( .A1(n2235), .A2(n1667), .B1(n2250), .B2(n1666), .ZN(n1371)
         );
  OAI22_X1 U2460 ( .A1(n2189), .A2(n1658), .B1(n1657), .B2(n2250), .ZN(n802)
         );
  OAI22_X1 U2461 ( .A1(n2189), .A2(n1665), .B1(n2250), .B2(n1664), .ZN(n1369)
         );
  OAI22_X1 U2462 ( .A1(n2235), .A2(n1662), .B1(n1661), .B2(n2250), .ZN(n1366)
         );
  OAI22_X1 U2463 ( .A1(n2235), .A2(n1666), .B1(n1665), .B2(n2250), .ZN(n1370)
         );
  OAI22_X1 U2464 ( .A1(n2188), .A2(n1659), .B1(n1978), .B2(n1658), .ZN(n1363)
         );
  OAI22_X1 U2465 ( .A1(n2155), .A2(n1570), .B1(n1569), .B2(n2245), .ZN(n1278)
         );
  OAI22_X1 U2466 ( .A1(n2156), .A2(n1571), .B1(n2245), .B2(n1570), .ZN(n1279)
         );
  OAI22_X1 U2467 ( .A1(n2156), .A2(n1575), .B1(n2246), .B2(n1574), .ZN(n1283)
         );
  OAI22_X1 U2468 ( .A1(n2156), .A2(n1580), .B1(n1579), .B2(n2245), .ZN(n1288)
         );
  OAI22_X1 U2469 ( .A1(n2156), .A2(n1579), .B1(n2246), .B2(n1578), .ZN(n1287)
         );
  OAI22_X1 U2470 ( .A1(n2154), .A2(n1569), .B1(n2246), .B2(n1568), .ZN(n1277)
         );
  OAI22_X1 U2471 ( .A1(n2155), .A2(n1578), .B1(n1577), .B2(n2245), .ZN(n1286)
         );
  OAI22_X1 U2472 ( .A1(n1573), .A2(n2227), .B1(n2245), .B2(n1572), .ZN(n1281)
         );
  OAI22_X1 U2473 ( .A1(n2227), .A2(n1577), .B1(n2245), .B2(n1576), .ZN(n1285)
         );
  OAI22_X1 U2474 ( .A1(n1572), .A2(n2227), .B1(n1571), .B2(n2246), .ZN(n1280)
         );
  OAI22_X1 U2475 ( .A1(n2227), .A2(n1574), .B1(n1573), .B2(n2245), .ZN(n1282)
         );
  OAI22_X1 U2476 ( .A1(n2227), .A2(n1576), .B1(n1575), .B2(n2246), .ZN(n1284)
         );
  OAI22_X1 U2477 ( .A1(n2160), .A2(n1535), .B1(n1534), .B2(n2244), .ZN(n1244)
         );
  OAI22_X1 U2478 ( .A1(n2160), .A2(n1537), .B1(n1536), .B2(n2243), .ZN(n1246)
         );
  OAI22_X1 U2479 ( .A1(n2160), .A2(n1544), .B1(n2243), .B2(n1543), .ZN(n1253)
         );
  OAI22_X1 U2480 ( .A1(n2159), .A2(n1543), .B1(n1542), .B2(n2244), .ZN(n1252)
         );
  OAI22_X1 U2481 ( .A1(n2160), .A2(n1539), .B1(n1538), .B2(n2243), .ZN(n1248)
         );
  OAI22_X1 U2482 ( .A1(n2226), .A2(n2000), .B1(n1556), .B2(n2244), .ZN(n1184)
         );
  OAI22_X1 U2483 ( .A1(n2226), .A2(n1546), .B1(n2244), .B2(n1545), .ZN(n1255)
         );
  OAI22_X1 U2484 ( .A1(n2160), .A2(n1552), .B1(n2243), .B2(n1551), .ZN(n1261)
         );
  OAI22_X1 U2485 ( .A1(n2160), .A2(n1555), .B1(n1554), .B2(n2243), .ZN(n1264)
         );
  OAI22_X1 U2486 ( .A1(n2226), .A2(n1533), .B1(n1532), .B2(n2244), .ZN(n692)
         );
  OAI22_X1 U2487 ( .A1(n1985), .A2(n1541), .B1(n1540), .B2(n2243), .ZN(n1250)
         );
  OAI22_X1 U2488 ( .A1(n2226), .A2(n1549), .B1(n1548), .B2(n2244), .ZN(n1258)
         );
  OAI22_X1 U2489 ( .A1(n2159), .A2(n1545), .B1(n1544), .B2(n2244), .ZN(n1254)
         );
  OAI22_X1 U2490 ( .A1(n2226), .A2(n1548), .B1(n2243), .B2(n1547), .ZN(n1257)
         );
  OAI22_X1 U2491 ( .A1(n2159), .A2(n1547), .B1(n1546), .B2(n2244), .ZN(n1256)
         );
  OAI22_X1 U2492 ( .A1(n2160), .A2(n1550), .B1(n2243), .B2(n1549), .ZN(n1259)
         );
  OAI22_X1 U2493 ( .A1(n2225), .A2(n1554), .B1(n2244), .B2(n1553), .ZN(n1263)
         );
  OAI22_X1 U2494 ( .A1(n2225), .A2(n1551), .B1(n1550), .B2(n2243), .ZN(n1260)
         );
  OAI22_X1 U2495 ( .A1(n1956), .A2(n1593), .B1(n1592), .B2(n2150), .ZN(n1300)
         );
  OAI22_X1 U2496 ( .A1(n2230), .A2(n1589), .B1(n1588), .B2(n2150), .ZN(n1296)
         );
  OAI22_X1 U2497 ( .A1(n1955), .A2(n1583), .B1(n1582), .B2(n2150), .ZN(n724)
         );
  OAI22_X1 U2498 ( .A1(n2230), .A2(n1585), .B1(n1584), .B2(n2150), .ZN(n1292)
         );
  OAI22_X1 U2499 ( .A1(n2230), .A2(n1591), .B1(n1590), .B2(n2150), .ZN(n1298)
         );
  OAI22_X1 U2500 ( .A1(n1956), .A2(n1587), .B1(n1586), .B2(n2150), .ZN(n1294)
         );
  OAI22_X1 U2501 ( .A1(n2230), .A2(n1934), .B1(n1606), .B2(n2150), .ZN(n1186)
         );
  OAI22_X1 U2502 ( .A1(n2152), .A2(n1753), .B1(n1752), .B2(n2256), .ZN(n1454)
         );
  OAI22_X1 U2503 ( .A1(n2152), .A2(n1747), .B1(n1746), .B2(n2256), .ZN(n1448)
         );
  OAI22_X1 U2504 ( .A1(n2153), .A2(n1750), .B1(n2255), .B2(n1749), .ZN(n1451)
         );
  OAI22_X1 U2505 ( .A1(n2152), .A2(n1749), .B1(n1748), .B2(n2256), .ZN(n1450)
         );
  OAI22_X1 U2506 ( .A1(n2152), .A2(n1745), .B1(n1744), .B2(n2255), .ZN(n1446)
         );
  OAI22_X1 U2507 ( .A1(n2152), .A2(n1748), .B1(n2255), .B2(n1747), .ZN(n1449)
         );
  OAI22_X1 U2508 ( .A1(n2152), .A2(n1744), .B1(n2255), .B2(n1743), .ZN(n1445)
         );
  OAI22_X1 U2509 ( .A1(n2153), .A2(n1746), .B1(n2255), .B2(n1745), .ZN(n1447)
         );
  OAI22_X1 U2510 ( .A1(n2011), .A2(n1754), .B1(n2256), .B2(n1753), .ZN(n1455)
         );
  OAI22_X1 U2511 ( .A1(n2153), .A2(n1752), .B1(n2255), .B2(n1751), .ZN(n1453)
         );
  OAI22_X1 U2512 ( .A1(n2153), .A2(n1751), .B1(n1750), .B2(n2255), .ZN(n1452)
         );
  OAI22_X1 U2513 ( .A1(n2153), .A2(n1755), .B1(n1754), .B2(n2256), .ZN(n1456)
         );
  XNOR2_X1 U2514 ( .A(b[13]), .B(n2002), .ZN(n1667) );
  XNOR2_X1 U2515 ( .A(b[21]), .B(n2287), .ZN(n1659) );
  XNOR2_X1 U2516 ( .A(b[15]), .B(n2289), .ZN(n1665) );
  XNOR2_X1 U2517 ( .A(b[19]), .B(n2289), .ZN(n1661) );
  XNOR2_X1 U2518 ( .A(b[17]), .B(n2287), .ZN(n1663) );
  INV_X1 U2519 ( .A(n345), .ZN(n343) );
  NAND2_X1 U2520 ( .A1(n345), .A2(n2127), .ZN(n336) );
  OAI22_X1 U2521 ( .A1(n2015), .A2(n1508), .B1(n1507), .B2(n2007), .ZN(n682)
         );
  OAI22_X1 U2522 ( .A1(n2014), .A2(n1513), .B1(n2241), .B2(n1512), .ZN(n1223)
         );
  OAI22_X1 U2523 ( .A1(n2014), .A2(n1518), .B1(n1517), .B2(n2241), .ZN(n1228)
         );
  OAI22_X1 U2524 ( .A1(n2014), .A2(n1515), .B1(n2241), .B2(n1514), .ZN(n1225)
         );
  OAI22_X1 U2525 ( .A1(n2015), .A2(n1514), .B1(n1513), .B2(n2007), .ZN(n1224)
         );
  OAI22_X1 U2526 ( .A1(n2014), .A2(n1509), .B1(n2007), .B2(n1508), .ZN(n1219)
         );
  OAI22_X1 U2527 ( .A1(n2015), .A2(n1511), .B1(n2241), .B2(n1510), .ZN(n1221)
         );
  OAI22_X1 U2528 ( .A1(n2014), .A2(n2264), .B1(n1531), .B2(n2241), .ZN(n1183)
         );
  OAI22_X1 U2529 ( .A1(n2014), .A2(n1517), .B1(n2007), .B2(n1516), .ZN(n1227)
         );
  OAI22_X1 U2530 ( .A1(n2015), .A2(n1510), .B1(n1509), .B2(n2007), .ZN(n1220)
         );
  OAI22_X1 U2531 ( .A1(n2014), .A2(n1516), .B1(n1515), .B2(n2241), .ZN(n1226)
         );
  OAI22_X1 U2532 ( .A1(n2014), .A2(n1512), .B1(n1511), .B2(n2007), .ZN(n1222)
         );
  XNOR2_X1 U2533 ( .A(b[13]), .B(n2304), .ZN(n1742) );
  XNOR2_X1 U2534 ( .A(b[19]), .B(n2305), .ZN(n1736) );
  XNOR2_X1 U2535 ( .A(b[21]), .B(n2304), .ZN(n1734) );
  XNOR2_X1 U2536 ( .A(b[11]), .B(n2025), .ZN(n1744) );
  XNOR2_X1 U2537 ( .A(b[15]), .B(n2304), .ZN(n1740) );
  NAND2_X1 U2538 ( .A1(n1071), .A2(n1084), .ZN(n591) );
  XNOR2_X1 U2539 ( .A(b[17]), .B(n2263), .ZN(n1513) );
  XNOR2_X1 U2540 ( .A(b[11]), .B(n2263), .ZN(n1519) );
  XNOR2_X1 U2541 ( .A(b[13]), .B(n2263), .ZN(n1517) );
  XNOR2_X1 U2542 ( .A(b[21]), .B(n1977), .ZN(n1509) );
  XNOR2_X1 U2543 ( .A(b[15]), .B(n2263), .ZN(n1515) );
  XNOR2_X1 U2544 ( .A(b[19]), .B(n2263), .ZN(n1511) );
  XNOR2_X1 U2545 ( .A(b[11]), .B(n2183), .ZN(n1769) );
  XNOR2_X1 U2546 ( .A(b[15]), .B(n2184), .ZN(n1765) );
  XNOR2_X1 U2547 ( .A(b[19]), .B(n2184), .ZN(n1761) );
  XNOR2_X1 U2548 ( .A(b[17]), .B(n2297), .ZN(n1713) );
  XNOR2_X1 U2549 ( .A(b[19]), .B(n2297), .ZN(n1711) );
  XNOR2_X1 U2550 ( .A(b[21]), .B(n2297), .ZN(n1709) );
  XNOR2_X1 U2551 ( .A(b[13]), .B(n2297), .ZN(n1717) );
  XNOR2_X1 U2552 ( .A(b[15]), .B(n2297), .ZN(n1715) );
  OAI22_X1 U2553 ( .A1(n1956), .A2(n1600), .B1(n2150), .B2(n1599), .ZN(n1307)
         );
  OAI22_X1 U2554 ( .A1(n1955), .A2(n1601), .B1(n1600), .B2(n2150), .ZN(n1308)
         );
  OAI22_X1 U2555 ( .A1(n1956), .A2(n1602), .B1(n2150), .B2(n1601), .ZN(n1309)
         );
  OAI22_X1 U2556 ( .A1(n2229), .A2(n1598), .B1(n2247), .B2(n1597), .ZN(n1305)
         );
  OAI22_X1 U2557 ( .A1(n2230), .A2(n1596), .B1(n2247), .B2(n1595), .ZN(n1303)
         );
  OAI22_X1 U2558 ( .A1(n2229), .A2(n1594), .B1(n2247), .B2(n1593), .ZN(n1301)
         );
  OAI22_X1 U2559 ( .A1(n2229), .A2(n1597), .B1(n1596), .B2(n2247), .ZN(n1304)
         );
  OAI22_X1 U2560 ( .A1(n2229), .A2(n1595), .B1(n1594), .B2(n2247), .ZN(n1302)
         );
  OAI22_X1 U2561 ( .A1(n1955), .A2(n1603), .B1(n1602), .B2(n2150), .ZN(n1310)
         );
  OAI22_X1 U2562 ( .A1(n1956), .A2(n1604), .B1(n2247), .B2(n1603), .ZN(n1311)
         );
  OAI22_X1 U2563 ( .A1(n2229), .A2(n1599), .B1(n1598), .B2(n2247), .ZN(n1306)
         );
  OAI22_X1 U2564 ( .A1(n1956), .A2(n1605), .B1(n1604), .B2(n2150), .ZN(n1312)
         );
  INV_X1 U2565 ( .A(n421), .ZN(n423) );
  OAI22_X1 U2566 ( .A1(n2193), .A2(n1637), .B1(n1636), .B2(n2037), .ZN(n1342)
         );
  OAI22_X1 U2567 ( .A1(n1993), .A2(n1636), .B1(n2036), .B2(n1635), .ZN(n1341)
         );
  OAI22_X1 U2568 ( .A1(n2193), .A2(n1634), .B1(n2036), .B2(n1633), .ZN(n1339)
         );
  OAI22_X1 U2569 ( .A1(n2193), .A2(n1635), .B1(n1634), .B2(n2037), .ZN(n1340)
         );
  INV_X1 U2570 ( .A(n772), .ZN(n773) );
  OAI22_X1 U2571 ( .A1(n2193), .A2(n1638), .B1(n2037), .B2(n1637), .ZN(n1343)
         );
  OAI22_X1 U2572 ( .A1(n2193), .A2(n1639), .B1(n1638), .B2(n2249), .ZN(n1344)
         );
  OAI22_X1 U2573 ( .A1(n1993), .A2(n1640), .B1(n2036), .B2(n1639), .ZN(n1345)
         );
  OAI22_X1 U2574 ( .A1(n2193), .A2(n1642), .B1(n2037), .B2(n1641), .ZN(n1347)
         );
  OAI22_X1 U2575 ( .A1(n1993), .A2(n1633), .B1(n1632), .B2(n2036), .ZN(n772)
         );
  OAI22_X1 U2576 ( .A1(n2208), .A2(n1641), .B1(n1640), .B2(n2249), .ZN(n1346)
         );
  OAI22_X1 U2577 ( .A1(n2193), .A2(n2284), .B1(n1656), .B2(n2249), .ZN(n1188)
         );
  OAI22_X1 U2578 ( .A1(n2208), .A2(n1643), .B1(n1642), .B2(n2249), .ZN(n1348)
         );
  XNOR2_X1 U2579 ( .A(n410), .B(n308), .ZN(product[38]) );
  NAND2_X1 U2580 ( .A1(n761), .A2(n774), .ZN(n461) );
  NAND2_X1 U2581 ( .A1(n540), .A2(n552), .ZN(n538) );
  AOI21_X1 U2582 ( .B1(n2072), .B2(n553), .A(n541), .ZN(n539) );
  OAI21_X1 U2583 ( .B1(n2001), .B2(n347), .A(n348), .ZN(n346) );
  OAI22_X1 U2584 ( .A1(n2130), .A2(n1483), .B1(n1482), .B2(n2239), .ZN(n676)
         );
  OAI22_X1 U2585 ( .A1(n1980), .A2(n1484), .B1(n2239), .B2(n1483), .ZN(n1195)
         );
  NAND2_X1 U2586 ( .A1(n717), .A2(n726), .ZN(n418) );
  OAI22_X1 U2587 ( .A1(n2130), .A2(n1485), .B1(n1484), .B2(n2238), .ZN(n1196)
         );
  OAI22_X1 U2588 ( .A1(n2130), .A2(n1491), .B1(n1490), .B2(n2238), .ZN(n1202)
         );
  OAI22_X1 U2589 ( .A1(n1980), .A2(n1486), .B1(n2239), .B2(n1485), .ZN(n1197)
         );
  OAI22_X1 U2590 ( .A1(n1980), .A2(n1488), .B1(n2239), .B2(n1487), .ZN(n1199)
         );
  OAI22_X1 U2591 ( .A1(n1980), .A2(n1490), .B1(n2238), .B2(n1489), .ZN(n1201)
         );
  OAI22_X1 U2592 ( .A1(n2130), .A2(n1487), .B1(n1486), .B2(n2238), .ZN(n1198)
         );
  OAI22_X1 U2593 ( .A1(n1980), .A2(n1492), .B1(n2238), .B2(n1491), .ZN(n1203)
         );
  OAI22_X1 U2594 ( .A1(n2130), .A2(n1493), .B1(n1492), .B2(n2239), .ZN(n1204)
         );
  OAI22_X1 U2595 ( .A1(n2222), .A2(n1938), .B1(n1506), .B2(n2238), .ZN(n1182)
         );
  OAI22_X1 U2596 ( .A1(n2130), .A2(n1489), .B1(n1488), .B2(n2238), .ZN(n1200)
         );
  OAI22_X1 U2597 ( .A1(n2011), .A2(n2306), .B1(n1756), .B2(n2255), .ZN(n1192)
         );
  OAI22_X1 U2598 ( .A1(n2152), .A2(n1738), .B1(n2256), .B2(n1737), .ZN(n1439)
         );
  OAI22_X1 U2599 ( .A1(n2152), .A2(n1741), .B1(n1740), .B2(n2256), .ZN(n1442)
         );
  OAI22_X1 U2600 ( .A1(n2153), .A2(n1740), .B1(n2255), .B2(n1739), .ZN(n1441)
         );
  INV_X1 U2601 ( .A(n916), .ZN(n917) );
  OAI22_X1 U2602 ( .A1(n2153), .A2(n1735), .B1(n1734), .B2(n2256), .ZN(n1436)
         );
  OAI22_X1 U2603 ( .A1(n2151), .A2(n1739), .B1(n1738), .B2(n2255), .ZN(n1440)
         );
  OAI22_X1 U2604 ( .A1(n2151), .A2(n1736), .B1(n2255), .B2(n1735), .ZN(n1437)
         );
  OAI22_X1 U2605 ( .A1(n2152), .A2(n1734), .B1(n2256), .B2(n1733), .ZN(n1435)
         );
  OAI22_X1 U2606 ( .A1(n2153), .A2(n1743), .B1(n1742), .B2(n2256), .ZN(n1444)
         );
  OAI22_X1 U2607 ( .A1(n2153), .A2(n1742), .B1(n2255), .B2(n1741), .ZN(n1443)
         );
  OAI22_X1 U2608 ( .A1(n2153), .A2(n1737), .B1(n1736), .B2(n2256), .ZN(n1438)
         );
  OAI22_X1 U2609 ( .A1(n2193), .A2(n1652), .B1(n2036), .B2(n1651), .ZN(n1357)
         );
  OAI22_X1 U2610 ( .A1(n2193), .A2(n1649), .B1(n1648), .B2(n2036), .ZN(n1354)
         );
  OAI22_X1 U2611 ( .A1(n1993), .A2(n1653), .B1(n1652), .B2(n2037), .ZN(n1358)
         );
  OAI22_X1 U2612 ( .A1(n1993), .A2(n1648), .B1(n2036), .B2(n1647), .ZN(n1353)
         );
  OAI22_X1 U2613 ( .A1(n1993), .A2(n1654), .B1(n2037), .B2(n1653), .ZN(n1359)
         );
  OAI22_X1 U2614 ( .A1(n1993), .A2(n1645), .B1(n1644), .B2(n2037), .ZN(n1350)
         );
  OAI22_X1 U2615 ( .A1(n1993), .A2(n1655), .B1(n1654), .B2(n2037), .ZN(n1360)
         );
  OAI22_X1 U2616 ( .A1(n2193), .A2(n1647), .B1(n1646), .B2(n2036), .ZN(n1352)
         );
  OAI22_X1 U2617 ( .A1(n1993), .A2(n1644), .B1(n2037), .B2(n1643), .ZN(n1349)
         );
  OAI22_X1 U2618 ( .A1(n1993), .A2(n1651), .B1(n1650), .B2(n2036), .ZN(n1356)
         );
  OAI22_X1 U2619 ( .A1(n2193), .A2(n1650), .B1(n2036), .B2(n1649), .ZN(n1355)
         );
  OAI22_X1 U2620 ( .A1(n2208), .A2(n1646), .B1(n2249), .B2(n1645), .ZN(n1351)
         );
  XNOR2_X1 U2621 ( .A(n397), .B(n307), .ZN(product[39]) );
  XNOR2_X1 U2622 ( .A(n2016), .B(n1237), .ZN(n939) );
  OR2_X1 U2623 ( .A1(n1215), .A2(n1237), .ZN(n938) );
  XNOR2_X1 U2624 ( .A(n388), .B(n306), .ZN(product[40]) );
  NAND2_X1 U2625 ( .A1(n775), .A2(n788), .ZN(n474) );
  XNOR2_X1 U2626 ( .A(n379), .B(n305), .ZN(product[41]) );
  OAI22_X1 U2627 ( .A1(n2015), .A2(n1522), .B1(n1521), .B2(n2007), .ZN(n1232)
         );
  OAI22_X1 U2628 ( .A1(n2014), .A2(n1519), .B1(n2241), .B2(n1518), .ZN(n1229)
         );
  OAI22_X1 U2629 ( .A1(n2015), .A2(n1521), .B1(n2007), .B2(n1520), .ZN(n1231)
         );
  OAI22_X1 U2630 ( .A1(n2014), .A2(n1520), .B1(n1519), .B2(n2007), .ZN(n1230)
         );
  OAI22_X1 U2631 ( .A1(n2013), .A2(n1525), .B1(n2007), .B2(n1524), .ZN(n1235)
         );
  OAI22_X1 U2632 ( .A1(n2223), .A2(n1524), .B1(n1523), .B2(n2241), .ZN(n1234)
         );
  OAI22_X1 U2633 ( .A1(n2223), .A2(n1526), .B1(n1525), .B2(n2240), .ZN(n1236)
         );
  OAI22_X1 U2634 ( .A1(n2013), .A2(n1523), .B1(n2007), .B2(n1522), .ZN(n1233)
         );
  OAI22_X1 U2635 ( .A1(n2223), .A2(n1529), .B1(n2240), .B2(n1528), .ZN(n1239)
         );
  OAI22_X1 U2636 ( .A1(n2223), .A2(n1527), .B1(n2240), .B2(n1526), .ZN(n1237)
         );
  XNOR2_X1 U2637 ( .A(b[13]), .B(n2291), .ZN(n1692) );
  XNOR2_X1 U2638 ( .A(b[21]), .B(n2291), .ZN(n1684) );
  XNOR2_X1 U2639 ( .A(b[11]), .B(n2291), .ZN(n1694) );
  XNOR2_X1 U2640 ( .A(b[15]), .B(n2291), .ZN(n1690) );
  XNOR2_X1 U2641 ( .A(n370), .B(n304), .ZN(product[42]) );
  OAI22_X1 U2642 ( .A1(n2147), .A2(n1931), .B1(n1731), .B2(n2254), .ZN(n1191)
         );
  OAI22_X1 U2643 ( .A1(n2006), .A2(n1718), .B1(n1717), .B2(n2253), .ZN(n1420)
         );
  OAI22_X1 U2644 ( .A1(n2149), .A2(n1717), .B1(n2253), .B2(n1716), .ZN(n1419)
         );
  OAI22_X1 U2645 ( .A1(n2147), .A2(n1713), .B1(n2254), .B2(n1712), .ZN(n1415)
         );
  OAI22_X1 U2646 ( .A1(n2148), .A2(n1715), .B1(n2253), .B2(n1714), .ZN(n1417)
         );
  OAI22_X1 U2647 ( .A1(n2148), .A2(n1709), .B1(n2253), .B2(n1708), .ZN(n1411)
         );
  OAI22_X1 U2648 ( .A1(n2149), .A2(n1716), .B1(n1715), .B2(n2254), .ZN(n1418)
         );
  OAI22_X1 U2649 ( .A1(n2149), .A2(n1708), .B1(n1707), .B2(n2253), .ZN(n874)
         );
  OAI22_X1 U2650 ( .A1(n2148), .A2(n1710), .B1(n1709), .B2(n2254), .ZN(n1412)
         );
  OAI22_X1 U2651 ( .A1(n2085), .A2(n1712), .B1(n1711), .B2(n2254), .ZN(n1414)
         );
  OAI22_X1 U2652 ( .A1(n2085), .A2(n1714), .B1(n1713), .B2(n2253), .ZN(n1416)
         );
  INV_X1 U2653 ( .A(n346), .ZN(n344) );
  AOI21_X1 U2654 ( .B1(n346), .B2(n2127), .A(n339), .ZN(n337) );
  XNOR2_X1 U2655 ( .A(b[17]), .B(n2277), .ZN(n1588) );
  XNOR2_X1 U2656 ( .A(b[15]), .B(n2277), .ZN(n1590) );
  XNOR2_X1 U2657 ( .A(b[13]), .B(n2275), .ZN(n1592) );
  XNOR2_X1 U2658 ( .A(b[21]), .B(n2274), .ZN(n1584) );
  XNOR2_X1 U2659 ( .A(b[19]), .B(n2275), .ZN(n1586) );
  XNOR2_X1 U2660 ( .A(b[11]), .B(n2277), .ZN(n1594) );
  XNOR2_X1 U2661 ( .A(n353), .B(n303), .ZN(product[43]) );
  OAI22_X1 U2662 ( .A1(n1980), .A2(n1497), .B1(n1496), .B2(n2239), .ZN(n1208)
         );
  OAI22_X1 U2663 ( .A1(n2130), .A2(n1496), .B1(n2238), .B2(n1495), .ZN(n1207)
         );
  OAI22_X1 U2664 ( .A1(n2130), .A2(n1502), .B1(n2238), .B2(n1501), .ZN(n1213)
         );
  OAI22_X1 U2665 ( .A1(n1980), .A2(n1495), .B1(n1494), .B2(n2238), .ZN(n1206)
         );
  OAI22_X1 U2666 ( .A1(n2130), .A2(n1501), .B1(n1500), .B2(n2239), .ZN(n1212)
         );
  OAI22_X1 U2667 ( .A1(n2130), .A2(n1494), .B1(n2239), .B2(n1493), .ZN(n1205)
         );
  OAI22_X1 U2668 ( .A1(n2222), .A2(n1503), .B1(n1502), .B2(n2239), .ZN(n1214)
         );
  OAI22_X1 U2669 ( .A1(n1980), .A2(n1500), .B1(n2238), .B2(n1499), .ZN(n1211)
         );
  OAI22_X1 U2670 ( .A1(n1980), .A2(n1504), .B1(n2238), .B2(n1503), .ZN(n1215)
         );
  OAI22_X1 U2671 ( .A1(n2222), .A2(n1499), .B1(n1498), .B2(n2239), .ZN(n1210)
         );
  OAI22_X1 U2672 ( .A1(n2222), .A2(n1505), .B1(n1504), .B2(n2239), .ZN(n1216)
         );
  OAI22_X1 U2673 ( .A1(n1980), .A2(n1498), .B1(n2238), .B2(n1497), .ZN(n1209)
         );
  OAI22_X1 U2674 ( .A1(n2225), .A2(n1553), .B1(n1552), .B2(n2244), .ZN(n1262)
         );
  OAI22_X1 U2675 ( .A1(n2223), .A2(n1530), .B1(n2241), .B2(n1529), .ZN(n1240)
         );
  OAI21_X1 U2676 ( .B1(n566), .B2(n538), .A(n539), .ZN(n537) );
  OAI22_X1 U2677 ( .A1(n2232), .A2(n1620), .B1(n1619), .B2(n2248), .ZN(n1326)
         );
  OAI22_X1 U2678 ( .A1(n2057), .A2(n1626), .B1(n1625), .B2(n2248), .ZN(n1332)
         );
  OAI22_X1 U2679 ( .A1(n2057), .A2(n1623), .B1(n2248), .B2(n1622), .ZN(n1329)
         );
  OAI22_X1 U2680 ( .A1(n2056), .A2(n1630), .B1(n1629), .B2(n2157), .ZN(n1336)
         );
  OAI22_X1 U2681 ( .A1(n2056), .A2(n1625), .B1(n2248), .B2(n1624), .ZN(n1331)
         );
  OAI22_X1 U2682 ( .A1(n2057), .A2(n1629), .B1(n2248), .B2(n1628), .ZN(n1335)
         );
  OAI22_X1 U2683 ( .A1(n2231), .A2(n1621), .B1(n2248), .B2(n1620), .ZN(n1327)
         );
  OAI22_X1 U2684 ( .A1(n2056), .A2(n1619), .B1(n2248), .B2(n1618), .ZN(n1325)
         );
  OAI22_X1 U2685 ( .A1(n2057), .A2(n1624), .B1(n1623), .B2(n2248), .ZN(n1330)
         );
  OAI22_X1 U2686 ( .A1(n2232), .A2(n1627), .B1(n2248), .B2(n1626), .ZN(n1333)
         );
  OAI22_X1 U2687 ( .A1(n2057), .A2(n1622), .B1(n1621), .B2(n2248), .ZN(n1328)
         );
  XNOR2_X1 U2688 ( .A(b[19]), .B(n1954), .ZN(n1636) );
  XNOR2_X1 U2689 ( .A(b[21]), .B(n1954), .ZN(n1634) );
  OAI22_X1 U2690 ( .A1(n2231), .A2(n1628), .B1(n1627), .B2(n2157), .ZN(n1334)
         );
  XNOR2_X1 U2691 ( .A(b[11]), .B(n1954), .ZN(n1644) );
  XNOR2_X1 U2692 ( .A(b[17]), .B(n1954), .ZN(n1638) );
  XNOR2_X1 U2693 ( .A(b[15]), .B(n1954), .ZN(n1640) );
  XNOR2_X1 U2694 ( .A(b[13]), .B(n1954), .ZN(n1642) );
  NAND2_X1 U2695 ( .A1(n489), .A2(n454), .ZN(n452) );
  AOI21_X1 U2696 ( .B1(n490), .B2(n454), .A(n455), .ZN(n453) );
  OAI22_X1 U2697 ( .A1(n2051), .A2(n1733), .B1(n1732), .B2(n2256), .ZN(n916)
         );
  OAI21_X1 U2698 ( .B1(n506), .B2(n452), .A(n453), .ZN(n451) );
  XNOR2_X1 U2699 ( .A(n462), .B(n313), .ZN(product[33]) );
  XOR2_X1 U2700 ( .A(n1975), .B(n321), .Z(product[25]) );
  OAI21_X1 U2701 ( .B1(n1975), .B2(n516), .A(n517), .ZN(n515) );
  OAI21_X1 U2702 ( .B1(n1974), .B2(n523), .A(n524), .ZN(n522) );
  OAI21_X1 U2703 ( .B1(n1976), .B2(n463), .A(n464), .ZN(n462) );
  OAI21_X1 U2704 ( .B1(n1974), .B2(n534), .A(n2060), .ZN(n533) );
  OAI21_X1 U2705 ( .B1(n1976), .B2(n476), .A(n477), .ZN(n475) );
  OAI21_X1 U2706 ( .B1(n1976), .B2(n487), .A(n488), .ZN(n486) );
  OAI21_X1 U2707 ( .B1(n1975), .B2(n498), .A(n499), .ZN(n497) );
  OAI21_X1 U2708 ( .B1(n1974), .B2(n2194), .A(n2207), .ZN(n504) );
  OAI22_X1 U2709 ( .A1(n2006), .A2(n1727), .B1(n2254), .B2(n1726), .ZN(n1429)
         );
  OAI22_X1 U2710 ( .A1(n1933), .A2(n1720), .B1(n1719), .B2(n2253), .ZN(n1422)
         );
  OAI22_X1 U2711 ( .A1(n1933), .A2(n1721), .B1(n2254), .B2(n1720), .ZN(n1423)
         );
  OAI22_X1 U2712 ( .A1(n1933), .A2(n1726), .B1(n1725), .B2(n2254), .ZN(n1428)
         );
  OAI22_X1 U2713 ( .A1(n2147), .A2(n1730), .B1(n1729), .B2(n2253), .ZN(n1432)
         );
  OAI22_X1 U2714 ( .A1(n1933), .A2(n1725), .B1(n2254), .B2(n1724), .ZN(n1427)
         );
  OAI22_X1 U2715 ( .A1(n2147), .A2(n1723), .B1(n2253), .B2(n1722), .ZN(n1425)
         );
  OAI22_X1 U2716 ( .A1(n2147), .A2(n1728), .B1(n1727), .B2(n2253), .ZN(n1430)
         );
  OAI22_X1 U2717 ( .A1(n1933), .A2(n1722), .B1(n1721), .B2(n2254), .ZN(n1424)
         );
  OAI22_X1 U2718 ( .A1(n2147), .A2(n1729), .B1(n2254), .B2(n1728), .ZN(n1431)
         );
  OAI22_X1 U2719 ( .A1(n2147), .A2(n1719), .B1(n2254), .B2(n1718), .ZN(n1421)
         );
  OAI22_X1 U2720 ( .A1(n2149), .A2(n1724), .B1(n1723), .B2(n2253), .ZN(n1426)
         );
  INV_X1 U2721 ( .A(n325), .ZN(product[47]) );
  AOI21_X1 U2722 ( .B1(n423), .B2(n356), .A(n359), .ZN(n355) );
  NAND2_X1 U2723 ( .A1(n422), .A2(n356), .ZN(n354) );
  OAI22_X1 U2724 ( .A1(n2155), .A2(n1563), .B1(n2246), .B2(n1562), .ZN(n1271)
         );
  OAI22_X1 U2725 ( .A1(n2155), .A2(n1566), .B1(n1565), .B2(n2246), .ZN(n1274)
         );
  OAI22_X1 U2726 ( .A1(n2156), .A2(n1561), .B1(n2245), .B2(n1560), .ZN(n1269)
         );
  OAI22_X1 U2727 ( .A1(n2155), .A2(n1567), .B1(n2245), .B2(n1566), .ZN(n1275)
         );
  OAI22_X1 U2728 ( .A1(n2155), .A2(n1564), .B1(n1563), .B2(n2245), .ZN(n1272)
         );
  OAI22_X1 U2729 ( .A1(n2156), .A2(n1560), .B1(n1559), .B2(n2245), .ZN(n1268)
         );
  OAI22_X1 U2730 ( .A1(n2156), .A2(n1990), .B1(n1581), .B2(n2245), .ZN(n1185)
         );
  OAI22_X1 U2731 ( .A1(n2156), .A2(n1559), .B1(n2246), .B2(n1558), .ZN(n1267)
         );
  OAI22_X1 U2732 ( .A1(n2155), .A2(n1565), .B1(n2246), .B2(n1564), .ZN(n1273)
         );
  INV_X1 U2733 ( .A(n706), .ZN(n707) );
  OAI22_X1 U2734 ( .A1(n2155), .A2(n1562), .B1(n1561), .B2(n2245), .ZN(n1270)
         );
  OAI22_X1 U2735 ( .A1(n2154), .A2(n1568), .B1(n1567), .B2(n2245), .ZN(n1276)
         );
  OAI22_X1 U2736 ( .A1(n2227), .A2(n1558), .B1(n1557), .B2(n2246), .ZN(n706)
         );
  XNOR2_X1 U2737 ( .A(n342), .B(n302), .ZN(product[44]) );
  OAI21_X1 U2738 ( .B1(n2107), .B2(n326), .A(n327), .ZN(n325) );
  OAI21_X1 U2739 ( .B1(n2214), .B2(n411), .A(n412), .ZN(n410) );
  OAI21_X1 U2740 ( .B1(n2215), .B2(n431), .A(n432), .ZN(n430) );
  OAI21_X1 U2741 ( .B1(n2215), .B2(n354), .A(n355), .ZN(n353) );
  OAI21_X1 U2742 ( .B1(n2108), .B2(n420), .A(n2001), .ZN(n419) );
  OAI21_X1 U2743 ( .B1(n2214), .B2(n398), .A(n399), .ZN(n397) );
  OAI21_X1 U2744 ( .B1(n2215), .B2(n438), .A(n439), .ZN(n437) );
  OAI21_X1 U2745 ( .B1(n301), .B2(n343), .A(n344), .ZN(n342) );
  OAI21_X1 U2746 ( .B1(n2214), .B2(n389), .A(n390), .ZN(n388) );
  OAI21_X1 U2747 ( .B1(n301), .B2(n371), .A(n372), .ZN(n370) );
  OAI21_X1 U2748 ( .B1(n301), .B2(n380), .A(n381), .ZN(n379) );
  OAI22_X1 U2749 ( .A1(n2100), .A2(n1691), .B1(n1690), .B2(n2251), .ZN(n1394)
         );
  OAI22_X1 U2750 ( .A1(n2074), .A2(n1686), .B1(n2251), .B2(n1685), .ZN(n1389)
         );
  OAI22_X1 U2751 ( .A1(n2074), .A2(n1689), .B1(n1688), .B2(n2251), .ZN(n1392)
         );
  OAI22_X1 U2752 ( .A1(n2100), .A2(n1690), .B1(n2252), .B2(n1689), .ZN(n1393)
         );
  OAI22_X1 U2753 ( .A1(n2100), .A2(n1687), .B1(n1686), .B2(n2252), .ZN(n1390)
         );
  OAI22_X1 U2754 ( .A1(n2074), .A2(n1692), .B1(n2252), .B2(n1691), .ZN(n1395)
         );
  OAI22_X1 U2755 ( .A1(n2100), .A2(n1685), .B1(n1684), .B2(n2252), .ZN(n1388)
         );
  OAI22_X1 U2756 ( .A1(n2074), .A2(n1688), .B1(n2251), .B2(n1687), .ZN(n1391)
         );
  INV_X1 U2757 ( .A(n836), .ZN(n837) );
  OAI22_X1 U2758 ( .A1(n2074), .A2(n1684), .B1(n2251), .B2(n1683), .ZN(n1387)
         );
  OAI22_X1 U2759 ( .A1(n2041), .A2(n2295), .B1(n1706), .B2(n2251), .ZN(n1190)
         );
  OAI22_X1 U2760 ( .A1(n2074), .A2(n1693), .B1(n1692), .B2(n2251), .ZN(n1396)
         );
  OAI22_X1 U2761 ( .A1(n2100), .A2(n1683), .B1(n1682), .B2(n2252), .ZN(n836)
         );
  INV_X2 U2762 ( .A(n2134), .ZN(n2230) );
  INV_X2 U2763 ( .A(n2168), .ZN(n2251) );
  INV_X2 U2764 ( .A(n2264), .ZN(n2263) );
  INV_X2 U2765 ( .A(n2273), .ZN(n2270) );
  INV_X2 U2766 ( .A(n2281), .ZN(n2280) );
  INV_X2 U2767 ( .A(n2296), .ZN(n2293) );
  INV_X1 U2768 ( .A(n2197), .ZN(n2244) );
  INV_X1 U2769 ( .A(n2192), .ZN(n2246) );
  INV_X1 U2770 ( .A(n2267), .ZN(n2266) );
  INV_X1 U2771 ( .A(a[19]), .ZN(n2267) );
  INV_X1 U2772 ( .A(n2273), .ZN(n2271) );
  INV_X1 U2773 ( .A(a[17]), .ZN(n2272) );
  INV_X1 U2774 ( .A(a[17]), .ZN(n2273) );
  INV_X1 U2775 ( .A(n2278), .ZN(n2277) );
  INV_X1 U2776 ( .A(a[15]), .ZN(n2278) );
  INV_X1 U2777 ( .A(a[13]), .ZN(n2281) );
  INV_X1 U2778 ( .A(a[11]), .ZN(n2284) );
  INV_X1 U2779 ( .A(a[11]), .ZN(n2285) );
  INV_X1 U2780 ( .A(n1982), .ZN(n2289) );
  INV_X1 U2781 ( .A(a[9]), .ZN(n2290) );
  INV_X1 U2782 ( .A(n2296), .ZN(n2294) );
  INV_X1 U2783 ( .A(a[7]), .ZN(n2295) );
  INV_X1 U2784 ( .A(a[7]), .ZN(n2296) );
  INV_X1 U2785 ( .A(n2302), .ZN(n2300) );
  INV_X1 U2786 ( .A(a[5]), .ZN(n2301) );
  INV_X1 U2787 ( .A(a[5]), .ZN(n2302) );
  INV_X1 U2788 ( .A(n2307), .ZN(n2305) );
  INV_X1 U2789 ( .A(a[3]), .ZN(n2306) );
  INV_X1 U2790 ( .A(a[3]), .ZN(n2307) );
  INV_X1 U2791 ( .A(n2311), .ZN(n2309) );
  INV_X1 U2792 ( .A(a[1]), .ZN(n2310) );
  INV_X1 U2793 ( .A(a[1]), .ZN(n2311) );
  INV_X2 U2794 ( .A(b[0]), .ZN(n2312) );
endmodule


module iir_filter_DW01_add_2 ( A, B, SUM, CI, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n17,
         n19, n21, n22, n23, n25, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n66, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n165, n167, n169, n170, n173, n243, n244, n245, n246,
         n247;

  NOR2_X1 U192 ( .A1(A[13]), .A2(B[13]), .ZN(n103) );
  OR2_X1 U193 ( .A1(A[15]), .A2(B[15]), .ZN(n243) );
  BUF_X2 U194 ( .A(n76), .Z(n1) );
  OR2_X1 U195 ( .A1(A[22]), .A2(B[22]), .ZN(n244) );
  OR2_X1 U196 ( .A1(A[11]), .A2(B[11]), .ZN(n245) );
  NOR2_X1 U197 ( .A1(A[16]), .A2(B[16]), .ZN(n74) );
  NOR2_X1 U198 ( .A1(A[14]), .A2(B[14]), .ZN(n92) );
  INV_X1 U199 ( .A(n47), .ZN(n45) );
  INV_X1 U200 ( .A(n49), .ZN(n47) );
  INV_X1 U201 ( .A(n99), .ZN(n97) );
  NAND2_X1 U202 ( .A1(n47), .A2(n31), .ZN(n29) );
  OR2_X1 U203 ( .A1(n49), .A2(n22), .ZN(n246) );
  NAND2_X1 U204 ( .A1(n115), .A2(n97), .ZN(n95) );
  NAND2_X1 U205 ( .A1(n88), .A2(n115), .ZN(n86) );
  INV_X1 U206 ( .A(n116), .ZN(n114) );
  INV_X1 U207 ( .A(n48), .ZN(n46) );
  AOI21_X1 U208 ( .B1(n116), .B2(n97), .A(n98), .ZN(n96) );
  INV_X1 U209 ( .A(n100), .ZN(n98) );
  INV_X1 U210 ( .A(n115), .ZN(n113) );
  INV_X1 U211 ( .A(n69), .ZN(n63) );
  INV_X1 U212 ( .A(n66), .ZN(n64) );
  INV_X1 U213 ( .A(n118), .ZN(n116) );
  NOR2_X1 U214 ( .A1(n99), .A2(n90), .ZN(n88) );
  AOI21_X1 U215 ( .B1(n48), .B2(n31), .A(n34), .ZN(n30) );
  INV_X1 U216 ( .A(n117), .ZN(n115) );
  INV_X1 U217 ( .A(n50), .ZN(n48) );
  INV_X1 U218 ( .A(n102), .ZN(n100) );
  INV_X1 U219 ( .A(n32), .ZN(n31) );
  INV_X1 U220 ( .A(n33), .ZN(n32) );
  INV_X1 U221 ( .A(n68), .ZN(n66) );
  INV_X1 U222 ( .A(n70), .ZN(n68) );
  NAND2_X1 U223 ( .A1(n115), .A2(n108), .ZN(n106) );
  NAND2_X1 U224 ( .A1(n69), .A2(n58), .ZN(n56) );
  AOI21_X1 U225 ( .B1(n51), .B2(n70), .A(n52), .ZN(n50) );
  OAI21_X1 U226 ( .B1(n35), .B2(n43), .A(n36), .ZN(n34) );
  OAI21_X1 U227 ( .B1(n71), .B2(n75), .A(n72), .ZN(n70) );
  XNOR2_X1 U228 ( .A(n28), .B(n3), .ZN(SUM[22]) );
  NAND2_X1 U229 ( .A1(n244), .A2(n27), .ZN(n3) );
  OAI21_X1 U230 ( .B1(n1), .B2(n29), .A(n30), .ZN(n28) );
  AOI21_X1 U231 ( .B1(n137), .B2(n77), .A(n78), .ZN(n76) );
  NOR2_X1 U232 ( .A1(n117), .A2(n79), .ZN(n77) );
  NOR2_X1 U233 ( .A1(n128), .A2(n121), .ZN(n119) );
  OAI21_X1 U234 ( .B1(n103), .B2(n111), .A(n104), .ZN(n102) );
  AOI21_X1 U235 ( .B1(n119), .B2(n131), .A(n120), .ZN(n118) );
  INV_X1 U236 ( .A(n137), .ZN(n136) );
  AOI21_X1 U237 ( .B1(n88), .B2(n116), .A(n89), .ZN(n87) );
  OAI21_X1 U238 ( .B1(n100), .B2(n90), .A(n93), .ZN(n89) );
  AOI21_X1 U239 ( .B1(n66), .B2(n58), .A(n59), .ZN(n57) );
  INV_X1 U240 ( .A(n61), .ZN(n59) );
  AOI21_X1 U241 ( .B1(n116), .B2(n108), .A(n109), .ZN(n107) );
  INV_X1 U242 ( .A(n111), .ZN(n109) );
  AOI21_X1 U243 ( .B1(n131), .B2(n126), .A(n127), .ZN(n125) );
  INV_X1 U244 ( .A(n129), .ZN(n127) );
  NOR2_X1 U245 ( .A1(n60), .A2(n53), .ZN(n51) );
  XOR2_X1 U246 ( .A(n1), .B(n9), .Z(SUM[16]) );
  NAND2_X1 U247 ( .A1(n170), .A2(n75), .ZN(n9) );
  INV_X1 U248 ( .A(n74), .ZN(n170) );
  INV_X1 U249 ( .A(n60), .ZN(n58) );
  OAI21_X1 U250 ( .B1(n1), .B2(n38), .A(n39), .ZN(n37) );
  NAND2_X1 U251 ( .A1(n47), .A2(n40), .ZN(n38) );
  AOI21_X1 U252 ( .B1(n48), .B2(n40), .A(n41), .ZN(n39) );
  INV_X1 U253 ( .A(n42), .ZN(n40) );
  XNOR2_X1 U254 ( .A(n73), .B(n8), .ZN(SUM[17]) );
  NAND2_X1 U255 ( .A1(n169), .A2(n72), .ZN(n8) );
  OAI21_X1 U256 ( .B1(n1), .B2(n74), .A(n75), .ZN(n73) );
  XNOR2_X1 U257 ( .A(n62), .B(n7), .ZN(SUM[18]) );
  NAND2_X1 U258 ( .A1(n58), .A2(n61), .ZN(n7) );
  OAI21_X1 U259 ( .B1(n1), .B2(n63), .A(n64), .ZN(n62) );
  XNOR2_X1 U260 ( .A(n55), .B(n6), .ZN(SUM[19]) );
  NAND2_X1 U261 ( .A1(n167), .A2(n54), .ZN(n6) );
  OAI21_X1 U262 ( .B1(n1), .B2(n56), .A(n57), .ZN(n55) );
  XNOR2_X1 U263 ( .A(n44), .B(n5), .ZN(SUM[20]) );
  NAND2_X1 U264 ( .A1(n40), .A2(n43), .ZN(n5) );
  OAI21_X1 U265 ( .B1(n1), .B2(n45), .A(n46), .ZN(n44) );
  XNOR2_X1 U266 ( .A(n85), .B(n10), .ZN(SUM[15]) );
  NAND2_X1 U267 ( .A1(n243), .A2(n84), .ZN(n10) );
  OAI21_X1 U268 ( .B1(n136), .B2(n86), .A(n87), .ZN(n85) );
  XNOR2_X1 U269 ( .A(n123), .B(n14), .ZN(SUM[11]) );
  NAND2_X1 U270 ( .A1(n245), .A2(n122), .ZN(n14) );
  OAI21_X1 U271 ( .B1(n136), .B2(n124), .A(n125), .ZN(n123) );
  XNOR2_X1 U272 ( .A(n112), .B(n13), .ZN(SUM[12]) );
  NAND2_X1 U273 ( .A1(n108), .A2(n111), .ZN(n13) );
  OAI21_X1 U274 ( .B1(n136), .B2(n113), .A(n114), .ZN(n112) );
  XNOR2_X1 U275 ( .A(n105), .B(n12), .ZN(SUM[13]) );
  NAND2_X1 U276 ( .A1(n173), .A2(n104), .ZN(n12) );
  OAI21_X1 U277 ( .B1(n136), .B2(n106), .A(n107), .ZN(n105) );
  INV_X1 U278 ( .A(n103), .ZN(n173) );
  XNOR2_X1 U279 ( .A(n94), .B(n11), .ZN(SUM[14]) );
  NAND2_X1 U280 ( .A1(n91), .A2(n93), .ZN(n11) );
  OAI21_X1 U281 ( .B1(n136), .B2(n95), .A(n96), .ZN(n94) );
  NAND2_X1 U282 ( .A1(n130), .A2(n119), .ZN(n117) );
  NAND2_X1 U283 ( .A1(n130), .A2(n126), .ZN(n124) );
  INV_X1 U284 ( .A(n128), .ZN(n126) );
  INV_X1 U285 ( .A(n91), .ZN(n90) );
  INV_X1 U286 ( .A(n92), .ZN(n91) );
  INV_X1 U287 ( .A(n43), .ZN(n41) );
  INV_X1 U288 ( .A(n21), .ZN(n19) );
  OAI21_X1 U289 ( .B1(n50), .B2(n22), .A(n23), .ZN(n21) );
  AOI21_X1 U290 ( .B1(n34), .B2(n244), .A(n25), .ZN(n23) );
  INV_X1 U291 ( .A(n27), .ZN(n25) );
  NOR2_X1 U292 ( .A1(n134), .A2(n132), .ZN(n130) );
  NOR2_X1 U293 ( .A1(A[8]), .A2(B[8]), .ZN(n134) );
  NOR2_X1 U294 ( .A1(A[20]), .A2(B[20]), .ZN(n42) );
  OAI21_X1 U295 ( .B1(n132), .B2(n135), .A(n133), .ZN(n131) );
  NAND2_X1 U296 ( .A1(A[8]), .A2(B[8]), .ZN(n135) );
  NAND2_X1 U297 ( .A1(A[9]), .A2(B[9]), .ZN(n133) );
  OAI21_X1 U298 ( .B1(n152), .B2(n138), .A(n139), .ZN(n137) );
  AOI21_X1 U299 ( .B1(n153), .B2(n159), .A(n154), .ZN(n152) );
  AOI21_X1 U300 ( .B1(n140), .B2(n147), .A(n141), .ZN(n139) );
  NAND2_X1 U301 ( .A1(n146), .A2(n140), .ZN(n138) );
  NOR2_X1 U302 ( .A1(A[11]), .A2(B[11]), .ZN(n121) );
  NOR2_X1 U303 ( .A1(A[17]), .A2(B[17]), .ZN(n71) );
  NOR2_X1 U304 ( .A1(A[9]), .A2(B[9]), .ZN(n132) );
  NOR2_X1 U305 ( .A1(A[18]), .A2(B[18]), .ZN(n60) );
  NOR2_X1 U306 ( .A1(A[7]), .A2(B[7]), .ZN(n142) );
  NOR2_X1 U307 ( .A1(A[3]), .A2(B[3]), .ZN(n155) );
  NOR2_X1 U308 ( .A1(A[5]), .A2(B[5]), .ZN(n148) );
  NOR2_X1 U309 ( .A1(n144), .A2(n142), .ZN(n140) );
  NOR2_X1 U310 ( .A1(A[6]), .A2(B[6]), .ZN(n144) );
  NOR2_X1 U311 ( .A1(A[12]), .A2(B[12]), .ZN(n110) );
  NOR2_X1 U312 ( .A1(A[15]), .A2(B[15]), .ZN(n83) );
  NOR2_X1 U313 ( .A1(A[10]), .A2(B[10]), .ZN(n128) );
  OAI21_X1 U314 ( .B1(n148), .B2(n151), .A(n149), .ZN(n147) );
  NAND2_X1 U315 ( .A1(A[4]), .A2(B[4]), .ZN(n151) );
  NAND2_X1 U316 ( .A1(A[5]), .A2(B[5]), .ZN(n149) );
  NAND2_X1 U317 ( .A1(A[16]), .A2(B[16]), .ZN(n75) );
  OAI21_X1 U318 ( .B1(n142), .B2(n145), .A(n143), .ZN(n141) );
  NAND2_X1 U319 ( .A1(A[6]), .A2(B[6]), .ZN(n145) );
  NAND2_X1 U320 ( .A1(A[7]), .A2(B[7]), .ZN(n143) );
  OAI21_X1 U321 ( .B1(n155), .B2(n158), .A(n156), .ZN(n154) );
  NAND2_X1 U322 ( .A1(A[3]), .A2(B[3]), .ZN(n156) );
  NAND2_X1 U323 ( .A1(A[2]), .A2(B[2]), .ZN(n158) );
  NOR2_X1 U324 ( .A1(A[19]), .A2(B[19]), .ZN(n53) );
  NAND2_X1 U325 ( .A1(A[18]), .A2(B[18]), .ZN(n61) );
  NAND2_X1 U326 ( .A1(A[14]), .A2(B[14]), .ZN(n93) );
  NOR2_X1 U327 ( .A1(A[21]), .A2(B[21]), .ZN(n35) );
  NAND2_X1 U328 ( .A1(A[12]), .A2(B[12]), .ZN(n111) );
  NAND2_X1 U329 ( .A1(A[20]), .A2(B[20]), .ZN(n43) );
  NOR2_X1 U330 ( .A1(n157), .A2(n155), .ZN(n153) );
  NOR2_X1 U331 ( .A1(A[2]), .A2(B[2]), .ZN(n157) );
  NOR2_X1 U332 ( .A1(n150), .A2(n148), .ZN(n146) );
  NOR2_X1 U333 ( .A1(A[4]), .A2(B[4]), .ZN(n150) );
  NAND2_X1 U334 ( .A1(A[13]), .A2(B[13]), .ZN(n104) );
  NAND2_X1 U335 ( .A1(A[21]), .A2(B[21]), .ZN(n36) );
  NAND2_X1 U336 ( .A1(A[19]), .A2(B[19]), .ZN(n54) );
  NAND2_X1 U337 ( .A1(A[10]), .A2(B[10]), .ZN(n129) );
  NAND2_X1 U338 ( .A1(A[22]), .A2(B[22]), .ZN(n27) );
  NAND2_X1 U339 ( .A1(A[17]), .A2(B[17]), .ZN(n72) );
  NAND2_X1 U340 ( .A1(A[11]), .A2(B[11]), .ZN(n122) );
  NAND2_X1 U341 ( .A1(A[15]), .A2(B[15]), .ZN(n84) );
  OAI21_X1 U342 ( .B1(n160), .B2(n162), .A(n161), .ZN(n159) );
  NAND2_X1 U343 ( .A1(A[1]), .A2(B[1]), .ZN(n161) );
  NOR2_X1 U344 ( .A1(A[1]), .A2(B[1]), .ZN(n160) );
  NAND2_X1 U345 ( .A1(A[0]), .A2(B[0]), .ZN(n162) );
  XNOR2_X1 U346 ( .A(n17), .B(n2), .ZN(SUM[23]) );
  NAND2_X1 U347 ( .A1(n247), .A2(n16), .ZN(n2) );
  OAI21_X1 U348 ( .B1(n1), .B2(n246), .A(n19), .ZN(n17) );
  NAND2_X1 U349 ( .A1(A[23]), .A2(B[23]), .ZN(n16) );
  OR2_X1 U350 ( .A1(A[23]), .A2(B[23]), .ZN(n247) );
  XNOR2_X1 U351 ( .A(n37), .B(n4), .ZN(SUM[21]) );
  NAND2_X1 U352 ( .A1(n165), .A2(n36), .ZN(n4) );
  OAI21_X1 U353 ( .B1(n118), .B2(n79), .A(n80), .ZN(n78) );
  NOR2_X1 U354 ( .A1(n110), .A2(n103), .ZN(n101) );
  NAND2_X1 U355 ( .A1(n101), .A2(n81), .ZN(n79) );
  INV_X1 U356 ( .A(n101), .ZN(n99) );
  INV_X1 U357 ( .A(n110), .ZN(n108) );
  NOR2_X1 U358 ( .A1(n92), .A2(n83), .ZN(n81) );
  OAI21_X1 U359 ( .B1(n83), .B2(n93), .A(n84), .ZN(n82) );
  AOI21_X1 U360 ( .B1(n81), .B2(n102), .A(n82), .ZN(n80) );
  NAND2_X1 U361 ( .A1(n33), .A2(n244), .ZN(n22) );
  NOR2_X1 U362 ( .A1(n42), .A2(n35), .ZN(n33) );
  INV_X1 U363 ( .A(n53), .ZN(n167) );
  OAI21_X1 U364 ( .B1(n53), .B2(n61), .A(n54), .ZN(n52) );
  INV_X1 U365 ( .A(n35), .ZN(n165) );
  NAND2_X1 U366 ( .A1(n69), .A2(n51), .ZN(n49) );
  INV_X1 U367 ( .A(n71), .ZN(n169) );
  NOR2_X1 U368 ( .A1(n74), .A2(n71), .ZN(n69) );
  OAI21_X1 U369 ( .B1(n121), .B2(n129), .A(n122), .ZN(n120) );
endmodule


module iir_filter_DW01_sub_1 ( A, B, DIFF, CI, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n17,
         n19, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n84, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n137, n138,
         n139, n141, n143, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, B_0_, n238,
         n239;
  assign DIFF[0] = B_0_;
  assign B_0_ = B[0];

  NOR2_X1 U188 ( .A1(n152), .A2(A[19]), .ZN(n42) );
  NOR2_X1 U189 ( .A1(n154), .A2(A[17]), .ZN(n60) );
  NOR2_X1 U190 ( .A1(n156), .A2(A[15]), .ZN(n78) );
  NOR2_X1 U191 ( .A1(n157), .A2(A[14]), .ZN(n89) );
  NOR2_X1 U192 ( .A1(n160), .A2(A[11]), .ZN(n103) );
  NOR2_X1 U193 ( .A1(n158), .A2(A[13]), .ZN(n92) );
  NOR2_X1 U194 ( .A1(n150), .A2(A[21]), .ZN(n25) );
  INV_X1 U195 ( .A(n65), .ZN(n63) );
  NAND2_X1 U196 ( .A1(n65), .A2(n47), .ZN(n45) );
  INV_X1 U197 ( .A(n50), .ZN(n48) );
  NOR2_X1 U198 ( .A1(n126), .A2(n121), .ZN(n120) );
  INV_X1 U199 ( .A(n67), .ZN(n65) );
  INV_X1 U200 ( .A(n114), .ZN(n113) );
  NAND2_X1 U201 ( .A1(n38), .A2(n65), .ZN(n36) );
  INV_X1 U202 ( .A(n127), .ZN(n126) );
  NAND2_X1 U203 ( .A1(n113), .A2(n106), .ZN(n105) );
  INV_X1 U204 ( .A(n133), .ZN(n132) );
  INV_X1 U205 ( .A(n49), .ZN(n47) );
  INV_X1 U206 ( .A(n66), .ZN(n64) );
  INV_X1 U207 ( .A(n87), .ZN(n81) );
  INV_X1 U208 ( .A(n84), .ZN(n82) );
  INV_X1 U209 ( .A(n95), .ZN(n94) );
  AOI21_X1 U210 ( .B1(n27), .B2(n95), .A(n28), .ZN(n1) );
  NOR2_X1 U211 ( .A1(n67), .A2(n29), .ZN(n27) );
  INV_X1 U212 ( .A(n68), .ZN(n66) );
  NOR2_X1 U213 ( .A1(n128), .A2(n133), .ZN(n127) );
  NAND2_X1 U214 ( .A1(n131), .A2(n129), .ZN(n128) );
  INV_X1 U215 ( .A(B[3]), .ZN(n129) );
  NOR2_X1 U216 ( .A1(n109), .A2(B[10]), .ZN(n106) );
  XOR2_X1 U217 ( .A(n126), .B(B[4]), .Z(DIFF[4]) );
  XOR2_X1 U218 ( .A(n111), .B(B[9]), .Z(DIFF[9]) );
  NAND2_X1 U219 ( .A1(n113), .A2(n112), .ZN(n111) );
  XOR2_X1 U220 ( .A(n118), .B(B[7]), .Z(DIFF[7]) );
  NAND2_X1 U221 ( .A1(n120), .A2(n119), .ZN(n118) );
  XOR2_X1 U222 ( .A(n130), .B(B[3]), .Z(DIFF[3]) );
  NAND2_X1 U223 ( .A1(n132), .A2(n131), .ZN(n130) );
  XOR2_X1 U224 ( .A(n107), .B(B[10]), .Z(DIFF[10]) );
  NAND2_X1 U225 ( .A1(n113), .A2(n108), .ZN(n107) );
  INV_X1 U226 ( .A(n109), .ZN(n108) );
  XNOR2_X1 U227 ( .A(n113), .B(B[8]), .ZN(DIFF[8]) );
  XNOR2_X1 U228 ( .A(B[2]), .B(n132), .ZN(DIFF[2]) );
  XNOR2_X1 U229 ( .A(n120), .B(B[6]), .ZN(DIFF[6]) );
  XNOR2_X1 U230 ( .A(n123), .B(B[5]), .ZN(DIFF[5]) );
  NOR2_X1 U231 ( .A1(n126), .A2(n124), .ZN(n123) );
  INV_X1 U232 ( .A(n125), .ZN(n124) );
  NAND2_X1 U233 ( .A1(n87), .A2(n69), .ZN(n67) );
  NAND2_X1 U234 ( .A1(n125), .A2(n122), .ZN(n121) );
  INV_X1 U235 ( .A(B[5]), .ZN(n122) );
  NAND2_X1 U236 ( .A1(n51), .A2(n31), .ZN(n29) );
  NAND2_X1 U237 ( .A1(n112), .A2(n110), .ZN(n109) );
  INV_X1 U238 ( .A(B[9]), .ZN(n110) );
  NAND2_X1 U239 ( .A1(n134), .A2(n135), .ZN(n133) );
  INV_X1 U240 ( .A(B[1]), .ZN(n134) );
  NAND2_X1 U241 ( .A1(n115), .A2(n127), .ZN(n114) );
  NOR2_X1 U242 ( .A1(n121), .A2(n116), .ZN(n115) );
  NAND2_X1 U243 ( .A1(n119), .A2(n117), .ZN(n116) );
  INV_X1 U244 ( .A(B[7]), .ZN(n117) );
  INV_X1 U245 ( .A(B[6]), .ZN(n119) );
  INV_X1 U246 ( .A(B[8]), .ZN(n112) );
  INV_X1 U247 ( .A(B[2]), .ZN(n131) );
  INV_X1 U248 ( .A(B[4]), .ZN(n125) );
  INV_X1 U249 ( .A(n86), .ZN(n84) );
  INV_X1 U250 ( .A(n88), .ZN(n86) );
  INV_X1 U251 ( .A(n51), .ZN(n49) );
  NAND2_X1 U252 ( .A1(n65), .A2(n58), .ZN(n56) );
  NAND2_X1 U253 ( .A1(n87), .A2(n76), .ZN(n74) );
  XNOR2_X1 U254 ( .A(B[1]), .B(n135), .ZN(DIFF[1]) );
  NOR2_X1 U255 ( .A1(n60), .A2(n53), .ZN(n51) );
  NOR2_X1 U256 ( .A1(n42), .A2(n33), .ZN(n31) );
  AOI21_X1 U257 ( .B1(n69), .B2(n88), .A(n70), .ZN(n68) );
  OAI21_X1 U258 ( .B1(n89), .B2(n93), .A(n90), .ZN(n88) );
  OAI21_X1 U259 ( .B1(n96), .B2(n114), .A(n97), .ZN(n95) );
  NAND2_X1 U260 ( .A1(n98), .A2(n106), .ZN(n96) );
  NOR2_X1 U261 ( .A1(n92), .A2(n89), .ZN(n87) );
  AOI21_X1 U262 ( .B1(n66), .B2(n58), .A(n59), .ZN(n57) );
  INV_X1 U263 ( .A(n61), .ZN(n59) );
  AOI21_X1 U264 ( .B1(n84), .B2(n76), .A(n77), .ZN(n75) );
  INV_X1 U265 ( .A(n79), .ZN(n77) );
  XOR2_X1 U266 ( .A(n94), .B(n12), .Z(DIFF[13]) );
  NAND2_X1 U267 ( .A1(n146), .A2(n93), .ZN(n12) );
  INV_X1 U268 ( .A(n92), .ZN(n146) );
  XNOR2_X1 U269 ( .A(n24), .B(n3), .ZN(DIFF[22]) );
  NAND2_X1 U270 ( .A1(n137), .A2(n23), .ZN(n3) );
  INV_X1 U271 ( .A(n22), .ZN(n137) );
  XNOR2_X1 U272 ( .A(n91), .B(n11), .ZN(DIFF[14]) );
  NAND2_X1 U273 ( .A1(n145), .A2(n90), .ZN(n11) );
  OAI21_X1 U274 ( .B1(n94), .B2(n92), .A(n93), .ZN(n91) );
  INV_X1 U275 ( .A(n89), .ZN(n145) );
  XNOR2_X1 U276 ( .A(n44), .B(n6), .ZN(DIFF[19]) );
  NAND2_X1 U277 ( .A1(n41), .A2(n43), .ZN(n6) );
  XNOR2_X1 U278 ( .A(n102), .B(n13), .ZN(DIFF[12]) );
  NAND2_X1 U279 ( .A1(n147), .A2(n101), .ZN(n13) );
  OAI21_X1 U280 ( .B1(n105), .B2(n103), .A(n104), .ZN(n102) );
  XNOR2_X1 U281 ( .A(n17), .B(n2), .ZN(DIFF[23]) );
  NAND2_X1 U282 ( .A1(n239), .A2(n16), .ZN(n2) );
  NAND2_X1 U283 ( .A1(n161), .A2(B[23]), .ZN(n16) );
  XNOR2_X1 U284 ( .A(n35), .B(n5), .ZN(DIFF[20]) );
  NAND2_X1 U285 ( .A1(n139), .A2(n34), .ZN(n5) );
  OAI21_X1 U286 ( .B1(n36), .B2(n94), .A(n37), .ZN(n35) );
  INV_X1 U287 ( .A(n33), .ZN(n139) );
  XNOR2_X1 U288 ( .A(n55), .B(n7), .ZN(DIFF[18]) );
  NAND2_X1 U289 ( .A1(n141), .A2(n54), .ZN(n7) );
  OAI21_X1 U290 ( .B1(n94), .B2(n56), .A(n57), .ZN(n55) );
  XNOR2_X1 U291 ( .A(n62), .B(n8), .ZN(DIFF[17]) );
  NAND2_X1 U292 ( .A1(n58), .A2(n61), .ZN(n8) );
  OAI21_X1 U293 ( .B1(n94), .B2(n63), .A(n64), .ZN(n62) );
  XNOR2_X1 U294 ( .A(n73), .B(n9), .ZN(DIFF[16]) );
  NAND2_X1 U295 ( .A1(n143), .A2(n72), .ZN(n9) );
  OAI21_X1 U296 ( .B1(n94), .B2(n74), .A(n75), .ZN(n73) );
  XNOR2_X1 U297 ( .A(n80), .B(n10), .ZN(DIFF[15]) );
  NAND2_X1 U298 ( .A1(n76), .A2(n79), .ZN(n10) );
  OAI21_X1 U299 ( .B1(n94), .B2(n81), .A(n82), .ZN(n80) );
  INV_X1 U300 ( .A(n60), .ZN(n58) );
  INV_X1 U301 ( .A(n78), .ZN(n76) );
  INV_X1 U302 ( .A(B[16]), .ZN(n155) );
  INV_X1 U303 ( .A(B[15]), .ZN(n156) );
  INV_X1 U304 ( .A(B[13]), .ZN(n158) );
  INV_X1 U305 ( .A(B[11]), .ZN(n160) );
  INV_X1 U306 ( .A(B[21]), .ZN(n150) );
  INV_X1 U307 ( .A(B[12]), .ZN(n159) );
  INV_X1 U308 ( .A(B[20]), .ZN(n151) );
  INV_X1 U309 ( .A(B[22]), .ZN(n149) );
  INV_X1 U310 ( .A(B_0_), .ZN(n135) );
  XOR2_X1 U311 ( .A(n105), .B(n14), .Z(DIFF[11]) );
  NAND2_X1 U312 ( .A1(n148), .A2(n104), .ZN(n14) );
  INV_X1 U313 ( .A(n103), .ZN(n148) );
  INV_X1 U314 ( .A(n21), .ZN(n19) );
  NAND2_X1 U315 ( .A1(n138), .A2(n26), .ZN(n4) );
  INV_X1 U316 ( .A(n25), .ZN(n138) );
  OR2_X1 U317 ( .A1(n25), .A2(n22), .ZN(n238) );
  OR2_X1 U318 ( .A1(n161), .A2(B[23]), .ZN(n239) );
  INV_X1 U319 ( .A(n41), .ZN(n40) );
  INV_X1 U320 ( .A(n42), .ZN(n41) );
  NOR2_X1 U321 ( .A1(n153), .A2(A[18]), .ZN(n53) );
  NOR2_X1 U322 ( .A1(n149), .A2(A[22]), .ZN(n22) );
  NOR2_X1 U323 ( .A1(n151), .A2(A[20]), .ZN(n33) );
  NOR2_X1 U324 ( .A1(n155), .A2(A[16]), .ZN(n71) );
  NAND2_X1 U325 ( .A1(n149), .A2(A[22]), .ZN(n23) );
  NAND2_X1 U326 ( .A1(n158), .A2(A[13]), .ZN(n93) );
  NAND2_X1 U327 ( .A1(n154), .A2(A[17]), .ZN(n61) );
  NAND2_X1 U328 ( .A1(n156), .A2(A[15]), .ZN(n79) );
  NAND2_X1 U329 ( .A1(n160), .A2(A[11]), .ZN(n104) );
  NAND2_X1 U330 ( .A1(n157), .A2(A[14]), .ZN(n90) );
  NAND2_X1 U331 ( .A1(n152), .A2(A[19]), .ZN(n43) );
  NAND2_X1 U332 ( .A1(n150), .A2(A[21]), .ZN(n26) );
  NAND2_X1 U333 ( .A1(n151), .A2(A[20]), .ZN(n34) );
  NAND2_X1 U334 ( .A1(n155), .A2(A[16]), .ZN(n72) );
  NAND2_X1 U335 ( .A1(n153), .A2(A[18]), .ZN(n54) );
  NAND2_X1 U336 ( .A1(n159), .A2(A[12]), .ZN(n101) );
  INV_X1 U337 ( .A(A[22]), .ZN(n161) );
  INV_X1 U338 ( .A(B[14]), .ZN(n157) );
  OAI21_X1 U339 ( .B1(n22), .B2(n26), .A(n23), .ZN(n21) );
  INV_X1 U340 ( .A(B[18]), .ZN(n153) );
  OAI21_X1 U341 ( .B1(n94), .B2(n45), .A(n46), .ZN(n44) );
  AOI21_X1 U342 ( .B1(n66), .B2(n47), .A(n48), .ZN(n46) );
  INV_X1 U343 ( .A(n52), .ZN(n50) );
  AOI21_X1 U344 ( .B1(n31), .B2(n52), .A(n32), .ZN(n30) );
  INV_X1 U345 ( .A(n99), .ZN(n97) );
  OAI21_X1 U346 ( .B1(n100), .B2(n104), .A(n101), .ZN(n99) );
  NOR2_X1 U347 ( .A1(n103), .A2(n100), .ZN(n98) );
  INV_X1 U348 ( .A(n100), .ZN(n147) );
  NOR2_X1 U349 ( .A1(n159), .A2(A[12]), .ZN(n100) );
  XOR2_X1 U350 ( .A(n1), .B(n4), .Z(DIFF[21]) );
  OAI21_X1 U351 ( .B1(n33), .B2(n43), .A(n34), .ZN(n32) );
  INV_X1 U352 ( .A(B[17]), .ZN(n154) );
  AOI21_X1 U353 ( .B1(n38), .B2(n66), .A(n39), .ZN(n37) );
  OAI21_X1 U354 ( .B1(n50), .B2(n40), .A(n43), .ZN(n39) );
  NOR2_X1 U355 ( .A1(n49), .A2(n40), .ZN(n38) );
  INV_X1 U356 ( .A(B[19]), .ZN(n152) );
  OAI21_X1 U357 ( .B1(n68), .B2(n29), .A(n30), .ZN(n28) );
  NOR2_X1 U358 ( .A1(n78), .A2(n71), .ZN(n69) );
  OAI21_X1 U359 ( .B1(n71), .B2(n79), .A(n72), .ZN(n70) );
  INV_X1 U360 ( .A(n71), .ZN(n143) );
  OAI21_X1 U361 ( .B1(n53), .B2(n61), .A(n54), .ZN(n52) );
  INV_X1 U362 ( .A(n53), .ZN(n141) );
  OAI21_X1 U363 ( .B1(n1), .B2(n25), .A(n26), .ZN(n24) );
  OAI21_X1 U364 ( .B1(n1), .B2(n238), .A(n19), .ZN(n17) );
endmodule


module iir_filter_DW01_add_1 ( A, B, SUM, CI, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n27, n28, n30, n32, n33, n34,
         n36, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n145, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n190, n193, n195, n197, n198, n199, n201,
         n203, n205, n206, n207, n208, n209, n211, n212, n213, n293, n295,
         n296, n297;

  OR2_X1 U242 ( .A1(A[22]), .A2(B[22]), .ZN(n293) );
  AND2_X1 U243 ( .A1(n295), .A2(n190), .ZN(SUM[0]) );
  OR2_X1 U244 ( .A1(A[0]), .A2(B[0]), .ZN(n295) );
  NOR2_X1 U245 ( .A1(A[4]), .A2(B[4]), .ZN(n174) );
  NOR2_X1 U246 ( .A1(A[14]), .A2(B[14]), .ZN(n103) );
  NOR2_X1 U247 ( .A1(A[10]), .A2(B[10]), .ZN(n139) );
  NOR2_X1 U248 ( .A1(A[12]), .A2(B[12]), .ZN(n121) );
  NOR2_X1 U249 ( .A1(A[5]), .A2(B[5]), .ZN(n169) );
  NOR2_X1 U250 ( .A1(A[13]), .A2(B[13]), .ZN(n114) );
  NOR2_X1 U251 ( .A1(A[15]), .A2(B[15]), .ZN(n94) );
  NOR2_X1 U252 ( .A1(A[7]), .A2(B[7]), .ZN(n161) );
  NOR2_X1 U253 ( .A1(A[8]), .A2(B[8]), .ZN(n153) );
  NOR2_X1 U254 ( .A1(A[2]), .A2(B[2]), .ZN(n183) );
  NOR2_X1 U255 ( .A1(A[6]), .A2(B[6]), .ZN(n164) );
  NOR2_X1 U256 ( .A1(A[1]), .A2(B[1]), .ZN(n187) );
  NOR2_X1 U257 ( .A1(A[18]), .A2(B[18]), .ZN(n71) );
  NOR2_X1 U258 ( .A1(A[20]), .A2(B[20]), .ZN(n53) );
  NOR2_X1 U259 ( .A1(A[17]), .A2(B[17]), .ZN(n82) );
  NOR2_X1 U260 ( .A1(A[19]), .A2(B[19]), .ZN(n64) );
  NOR2_X1 U261 ( .A1(A[21]), .A2(B[21]), .ZN(n46) );
  NOR2_X1 U262 ( .A1(A[16]), .A2(B[16]), .ZN(n85) );
  NAND2_X1 U263 ( .A1(n126), .A2(n108), .ZN(n106) );
  INV_X1 U264 ( .A(n126), .ZN(n124) );
  INV_X1 U265 ( .A(n58), .ZN(n56) );
  AOI21_X1 U266 ( .B1(n127), .B2(n108), .A(n109), .ZN(n107) );
  INV_X1 U267 ( .A(n111), .ZN(n109) );
  INV_X1 U268 ( .A(n128), .ZN(n126) );
  INV_X1 U269 ( .A(n60), .ZN(n58) );
  INV_X1 U270 ( .A(n110), .ZN(n108) );
  NAND2_X1 U271 ( .A1(n99), .A2(n126), .ZN(n97) );
  NAND2_X1 U272 ( .A1(n58), .A2(n42), .ZN(n40) );
  INV_X1 U273 ( .A(n127), .ZN(n125) );
  INV_X1 U274 ( .A(n59), .ZN(n57) );
  OR2_X1 U275 ( .A1(n60), .A2(n33), .ZN(n296) );
  INV_X1 U276 ( .A(n148), .ZN(n142) );
  INV_X1 U277 ( .A(n76), .ZN(n74) );
  INV_X1 U278 ( .A(n145), .ZN(n143) );
  INV_X1 U279 ( .A(n77), .ZN(n75) );
  INV_X1 U280 ( .A(n156), .ZN(n155) );
  BUF_X1 U281 ( .A(n87), .Z(n1) );
  AOI21_X1 U282 ( .B1(n156), .B2(n88), .A(n89), .ZN(n87) );
  NOR2_X1 U283 ( .A1(n128), .A2(n90), .ZN(n88) );
  OAI21_X1 U284 ( .B1(n129), .B2(n90), .A(n91), .ZN(n89) );
  AOI21_X1 U285 ( .B1(n176), .B2(n167), .A(n168), .ZN(n166) );
  NOR2_X1 U286 ( .A1(n110), .A2(n101), .ZN(n99) );
  AOI21_X1 U287 ( .B1(n59), .B2(n42), .A(n45), .ZN(n41) );
  NAND2_X1 U288 ( .A1(n148), .A2(n130), .ZN(n128) );
  INV_X1 U289 ( .A(n129), .ZN(n127) );
  INV_X1 U290 ( .A(n147), .ZN(n145) );
  INV_X1 U291 ( .A(n149), .ZN(n147) );
  INV_X1 U292 ( .A(n61), .ZN(n59) );
  NAND2_X1 U293 ( .A1(n112), .A2(n92), .ZN(n90) );
  INV_X1 U294 ( .A(n177), .ZN(n176) );
  NAND2_X1 U295 ( .A1(n80), .A2(n62), .ZN(n60) );
  NAND2_X1 U296 ( .A1(n44), .A2(n293), .ZN(n33) );
  INV_X1 U297 ( .A(n113), .ZN(n111) );
  INV_X1 U298 ( .A(n112), .ZN(n110) );
  INV_X1 U299 ( .A(n186), .ZN(n185) );
  INV_X1 U300 ( .A(n43), .ZN(n42) );
  INV_X1 U301 ( .A(n44), .ZN(n43) );
  INV_X1 U302 ( .A(n79), .ZN(n77) );
  INV_X1 U303 ( .A(n81), .ZN(n79) );
  INV_X1 U304 ( .A(n78), .ZN(n76) );
  INV_X1 U305 ( .A(n80), .ZN(n78) );
  NAND2_X1 U306 ( .A1(n126), .A2(n119), .ZN(n117) );
  NAND2_X1 U307 ( .A1(n58), .A2(n51), .ZN(n49) );
  NAND2_X1 U308 ( .A1(n76), .A2(n69), .ZN(n67) );
  NAND2_X1 U309 ( .A1(n148), .A2(n137), .ZN(n135) );
  XOR2_X1 U310 ( .A(n166), .B(n19), .Z(SUM[6]) );
  NAND2_X1 U311 ( .A1(n208), .A2(n165), .ZN(n19) );
  INV_X1 U312 ( .A(n164), .ZN(n208) );
  XOR2_X1 U313 ( .A(n155), .B(n17), .Z(SUM[8]) );
  NAND2_X1 U314 ( .A1(n206), .A2(n154), .ZN(n17) );
  INV_X1 U315 ( .A(n153), .ZN(n206) );
  XOR2_X1 U316 ( .A(n171), .B(n20), .Z(SUM[5]) );
  NAND2_X1 U317 ( .A1(n209), .A2(n170), .ZN(n20) );
  AOI21_X1 U318 ( .B1(n176), .B2(n172), .A(n173), .ZN(n171) );
  INV_X1 U319 ( .A(n169), .ZN(n209) );
  XOR2_X1 U320 ( .A(n185), .B(n23), .Z(SUM[2]) );
  NAND2_X1 U321 ( .A1(n212), .A2(n184), .ZN(n23) );
  INV_X1 U322 ( .A(n183), .ZN(n212) );
  XOR2_X1 U323 ( .A(n24), .B(n190), .Z(SUM[1]) );
  NAND2_X1 U324 ( .A1(n213), .A2(n188), .ZN(n24) );
  INV_X1 U325 ( .A(n187), .ZN(n213) );
  XNOR2_X1 U326 ( .A(n141), .B(n15), .ZN(SUM[10]) );
  NAND2_X1 U327 ( .A1(n137), .A2(n140), .ZN(n15) );
  OAI21_X1 U328 ( .B1(n155), .B2(n142), .A(n143), .ZN(n141) );
  XNOR2_X1 U329 ( .A(n163), .B(n18), .ZN(SUM[7]) );
  NAND2_X1 U330 ( .A1(n207), .A2(n162), .ZN(n18) );
  OAI21_X1 U331 ( .B1(n166), .B2(n164), .A(n165), .ZN(n163) );
  INV_X1 U332 ( .A(n161), .ZN(n207) );
  XNOR2_X1 U333 ( .A(n152), .B(n16), .ZN(SUM[9]) );
  NAND2_X1 U334 ( .A1(n205), .A2(n151), .ZN(n16) );
  OAI21_X1 U335 ( .B1(n155), .B2(n153), .A(n154), .ZN(n152) );
  INV_X1 U336 ( .A(n150), .ZN(n205) );
  XNOR2_X1 U337 ( .A(n182), .B(n22), .ZN(SUM[3]) );
  NAND2_X1 U338 ( .A1(n211), .A2(n181), .ZN(n22) );
  OAI21_X1 U339 ( .B1(n185), .B2(n183), .A(n184), .ZN(n182) );
  XNOR2_X1 U340 ( .A(n176), .B(n21), .ZN(SUM[4]) );
  NAND2_X1 U341 ( .A1(n172), .A2(n175), .ZN(n21) );
  NAND2_X1 U342 ( .A1(n197), .A2(n83), .ZN(n8) );
  XNOR2_X1 U343 ( .A(n66), .B(n6), .ZN(SUM[19]) );
  NAND2_X1 U344 ( .A1(n195), .A2(n65), .ZN(n6) );
  OAI21_X1 U345 ( .B1(n1), .B2(n67), .A(n68), .ZN(n66) );
  XNOR2_X1 U346 ( .A(n105), .B(n11), .ZN(SUM[14]) );
  NAND2_X1 U347 ( .A1(n102), .A2(n104), .ZN(n11) );
  OAI21_X1 U348 ( .B1(n155), .B2(n106), .A(n107), .ZN(n105) );
  AOI21_X1 U349 ( .B1(n130), .B2(n149), .A(n131), .ZN(n129) );
  AOI21_X1 U350 ( .B1(n62), .B2(n81), .A(n63), .ZN(n61) );
  OAI21_X1 U351 ( .B1(n64), .B2(n72), .A(n65), .ZN(n63) );
  AOI21_X1 U352 ( .B1(n178), .B2(n186), .A(n179), .ZN(n177) );
  OAI21_X1 U353 ( .B1(n114), .B2(n122), .A(n115), .ZN(n113) );
  OAI21_X1 U354 ( .B1(n82), .B2(n86), .A(n83), .ZN(n81) );
  OAI21_X1 U355 ( .B1(n187), .B2(n190), .A(n188), .ZN(n186) );
  OAI21_X1 U356 ( .B1(n169), .B2(n175), .A(n170), .ZN(n168) );
  OAI21_X1 U357 ( .B1(n177), .B2(n157), .A(n158), .ZN(n156) );
  NAND2_X1 U358 ( .A1(n167), .A2(n159), .ZN(n157) );
  AOI21_X1 U359 ( .B1(n159), .B2(n168), .A(n160), .ZN(n158) );
  NOR2_X1 U360 ( .A1(n164), .A2(n161), .ZN(n159) );
  OAI21_X1 U361 ( .B1(n46), .B2(n54), .A(n47), .ZN(n45) );
  NAND2_X1 U362 ( .A1(n69), .A2(n72), .ZN(n7) );
  OAI21_X1 U363 ( .B1(n1), .B2(n74), .A(n75), .ZN(n73) );
  NOR2_X1 U364 ( .A1(n174), .A2(n169), .ZN(n167) );
  NOR2_X1 U365 ( .A1(n71), .A2(n64), .ZN(n62) );
  NOR2_X1 U366 ( .A1(n103), .A2(n94), .ZN(n92) );
  NOR2_X1 U367 ( .A1(n121), .A2(n114), .ZN(n112) );
  NOR2_X1 U368 ( .A1(n85), .A2(n82), .ZN(n80) );
  NOR2_X1 U369 ( .A1(n53), .A2(n46), .ZN(n44) );
  AOI21_X1 U370 ( .B1(n92), .B2(n113), .A(n93), .ZN(n91) );
  OAI21_X1 U371 ( .B1(n94), .B2(n104), .A(n95), .ZN(n93) );
  AOI21_X1 U372 ( .B1(n99), .B2(n127), .A(n100), .ZN(n98) );
  OAI21_X1 U373 ( .B1(n111), .B2(n101), .A(n104), .ZN(n100) );
  AOI21_X1 U374 ( .B1(n127), .B2(n119), .A(n120), .ZN(n118) );
  INV_X1 U375 ( .A(n122), .ZN(n120) );
  AOI21_X1 U376 ( .B1(n145), .B2(n137), .A(n138), .ZN(n136) );
  INV_X1 U377 ( .A(n140), .ZN(n138) );
  AOI21_X1 U378 ( .B1(n59), .B2(n51), .A(n52), .ZN(n50) );
  INV_X1 U379 ( .A(n54), .ZN(n52) );
  AOI21_X1 U380 ( .B1(n77), .B2(n69), .A(n70), .ZN(n68) );
  INV_X1 U381 ( .A(n72), .ZN(n70) );
  OAI21_X1 U382 ( .B1(n161), .B2(n165), .A(n162), .ZN(n160) );
  INV_X1 U383 ( .A(n121), .ZN(n119) );
  INV_X1 U384 ( .A(n53), .ZN(n51) );
  INV_X1 U385 ( .A(n71), .ZN(n69) );
  INV_X1 U386 ( .A(n139), .ZN(n137) );
  XOR2_X1 U387 ( .A(n1), .B(n9), .Z(SUM[16]) );
  NAND2_X1 U388 ( .A1(n198), .A2(n86), .ZN(n9) );
  INV_X1 U389 ( .A(n85), .ZN(n198) );
  XNOR2_X1 U390 ( .A(n96), .B(n10), .ZN(SUM[15]) );
  NAND2_X1 U391 ( .A1(n199), .A2(n95), .ZN(n10) );
  OAI21_X1 U392 ( .B1(n155), .B2(n97), .A(n98), .ZN(n96) );
  XNOR2_X1 U393 ( .A(n116), .B(n12), .ZN(SUM[13]) );
  NAND2_X1 U394 ( .A1(n201), .A2(n115), .ZN(n12) );
  OAI21_X1 U395 ( .B1(n155), .B2(n117), .A(n118), .ZN(n116) );
  XNOR2_X1 U396 ( .A(n134), .B(n14), .ZN(SUM[11]) );
  NAND2_X1 U397 ( .A1(n203), .A2(n133), .ZN(n14) );
  OAI21_X1 U398 ( .B1(n155), .B2(n135), .A(n136), .ZN(n134) );
  XNOR2_X1 U399 ( .A(n48), .B(n4), .ZN(SUM[21]) );
  NAND2_X1 U400 ( .A1(n193), .A2(n47), .ZN(n4) );
  OAI21_X1 U401 ( .B1(n1), .B2(n49), .A(n50), .ZN(n48) );
  XNOR2_X1 U402 ( .A(n123), .B(n13), .ZN(SUM[12]) );
  NAND2_X1 U403 ( .A1(n119), .A2(n122), .ZN(n13) );
  OAI21_X1 U404 ( .B1(n155), .B2(n124), .A(n125), .ZN(n123) );
  INV_X1 U405 ( .A(n174), .ZN(n172) );
  INV_X1 U406 ( .A(n102), .ZN(n101) );
  INV_X1 U407 ( .A(n103), .ZN(n102) );
  XNOR2_X1 U408 ( .A(n55), .B(n5), .ZN(SUM[20]) );
  NAND2_X1 U409 ( .A1(n51), .A2(n54), .ZN(n5) );
  OAI21_X1 U410 ( .B1(n1), .B2(n56), .A(n57), .ZN(n55) );
  XNOR2_X1 U411 ( .A(n39), .B(n3), .ZN(SUM[22]) );
  NAND2_X1 U412 ( .A1(n293), .A2(n38), .ZN(n3) );
  OAI21_X1 U413 ( .B1(n1), .B2(n40), .A(n41), .ZN(n39) );
  INV_X1 U414 ( .A(n94), .ZN(n199) );
  INV_X1 U415 ( .A(n114), .ZN(n201) );
  INV_X1 U416 ( .A(n46), .ZN(n193) );
  INV_X1 U417 ( .A(n64), .ZN(n195) );
  INV_X1 U418 ( .A(n82), .ZN(n197) );
  INV_X1 U419 ( .A(n175), .ZN(n173) );
  INV_X1 U420 ( .A(n32), .ZN(n30) );
  OAI21_X1 U421 ( .B1(n61), .B2(n33), .A(n34), .ZN(n32) );
  AOI21_X1 U422 ( .B1(n45), .B2(n293), .A(n36), .ZN(n34) );
  INV_X1 U423 ( .A(n38), .ZN(n36) );
  INV_X1 U424 ( .A(n132), .ZN(n203) );
  XNOR2_X1 U425 ( .A(n28), .B(n2), .ZN(SUM[23]) );
  NAND2_X1 U426 ( .A1(n297), .A2(n27), .ZN(n2) );
  OAI21_X1 U427 ( .B1(n1), .B2(n296), .A(n30), .ZN(n28) );
  NAND2_X1 U428 ( .A1(A[23]), .A2(B[23]), .ZN(n27) );
  NOR2_X1 U429 ( .A1(A[9]), .A2(B[9]), .ZN(n150) );
  NOR2_X1 U430 ( .A1(A[11]), .A2(B[11]), .ZN(n132) );
  NAND2_X1 U431 ( .A1(A[4]), .A2(B[4]), .ZN(n175) );
  NAND2_X1 U432 ( .A1(A[12]), .A2(B[12]), .ZN(n122) );
  NAND2_X1 U433 ( .A1(A[18]), .A2(B[18]), .ZN(n72) );
  NAND2_X1 U434 ( .A1(A[6]), .A2(B[6]), .ZN(n165) );
  NAND2_X1 U435 ( .A1(A[14]), .A2(B[14]), .ZN(n104) );
  NAND2_X1 U436 ( .A1(A[20]), .A2(B[20]), .ZN(n54) );
  NAND2_X1 U437 ( .A1(A[0]), .A2(B[0]), .ZN(n190) );
  NAND2_X1 U438 ( .A1(A[16]), .A2(B[16]), .ZN(n86) );
  NAND2_X1 U439 ( .A1(A[10]), .A2(B[10]), .ZN(n140) );
  NAND2_X1 U440 ( .A1(A[2]), .A2(B[2]), .ZN(n184) );
  NAND2_X1 U441 ( .A1(A[8]), .A2(B[8]), .ZN(n154) );
  NAND2_X1 U442 ( .A1(A[22]), .A2(B[22]), .ZN(n38) );
  NAND2_X1 U443 ( .A1(A[1]), .A2(B[1]), .ZN(n188) );
  NAND2_X1 U444 ( .A1(A[5]), .A2(B[5]), .ZN(n170) );
  NAND2_X1 U445 ( .A1(A[7]), .A2(B[7]), .ZN(n162) );
  NAND2_X1 U446 ( .A1(A[13]), .A2(B[13]), .ZN(n115) );
  NAND2_X1 U447 ( .A1(A[15]), .A2(B[15]), .ZN(n95) );
  NAND2_X1 U448 ( .A1(A[17]), .A2(B[17]), .ZN(n83) );
  NAND2_X1 U449 ( .A1(A[19]), .A2(B[19]), .ZN(n65) );
  NAND2_X1 U450 ( .A1(A[21]), .A2(B[21]), .ZN(n47) );
  NAND2_X1 U451 ( .A1(A[11]), .A2(B[11]), .ZN(n133) );
  NAND2_X1 U452 ( .A1(A[9]), .A2(B[9]), .ZN(n151) );
  NAND2_X1 U453 ( .A1(A[3]), .A2(B[3]), .ZN(n181) );
  OR2_X1 U454 ( .A1(A[23]), .A2(B[23]), .ZN(n297) );
  NOR2_X1 U455 ( .A1(n139), .A2(n132), .ZN(n130) );
  OAI21_X1 U456 ( .B1(n132), .B2(n140), .A(n133), .ZN(n131) );
  NOR2_X1 U457 ( .A1(A[3]), .A2(B[3]), .ZN(n180) );
  OAI21_X1 U458 ( .B1(n180), .B2(n184), .A(n181), .ZN(n179) );
  NOR2_X1 U459 ( .A1(n183), .A2(n180), .ZN(n178) );
  INV_X1 U460 ( .A(n180), .ZN(n211) );
  XNOR2_X1 U461 ( .A(n73), .B(n7), .ZN(SUM[18]) );
  NOR2_X1 U462 ( .A1(n153), .A2(n150), .ZN(n148) );
  OAI21_X1 U463 ( .B1(n150), .B2(n154), .A(n151), .ZN(n149) );
  XNOR2_X1 U464 ( .A(n84), .B(n8), .ZN(SUM[17]) );
  OAI21_X1 U465 ( .B1(n1), .B2(n85), .A(n86), .ZN(n84) );
endmodule


module iir_filter_DW01_add_6 ( A, B, SUM, CI, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n27, n28, n30, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n145, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n190, n192, n193, n195, n197,
         n198, n199, n201, n203, n205, n206, n207, n208, n209, n211, n212,
         n213, n294, n295, n296;

  AND2_X1 U242 ( .A1(n294), .A2(n190), .ZN(SUM[0]) );
  INV_X2 U243 ( .A(n156), .ZN(n155) );
  NOR2_X1 U244 ( .A1(A[4]), .A2(B[4]), .ZN(n174) );
  NOR2_X1 U245 ( .A1(A[20]), .A2(B[20]), .ZN(n53) );
  NOR2_X1 U246 ( .A1(A[18]), .A2(B[18]), .ZN(n71) );
  NOR2_X1 U247 ( .A1(A[10]), .A2(B[10]), .ZN(n139) );
  NOR2_X1 U248 ( .A1(A[14]), .A2(B[14]), .ZN(n103) );
  NOR2_X1 U249 ( .A1(A[12]), .A2(B[12]), .ZN(n121) );
  NOR2_X1 U250 ( .A1(A[7]), .A2(B[7]), .ZN(n161) );
  NOR2_X1 U251 ( .A1(A[5]), .A2(B[5]), .ZN(n169) );
  NOR2_X1 U252 ( .A1(A[21]), .A2(B[21]), .ZN(n46) );
  NOR2_X1 U253 ( .A1(A[3]), .A2(B[3]), .ZN(n180) );
  NOR2_X1 U254 ( .A1(A[19]), .A2(B[19]), .ZN(n64) );
  NOR2_X1 U255 ( .A1(A[17]), .A2(B[17]), .ZN(n82) );
  NOR2_X1 U256 ( .A1(A[11]), .A2(B[11]), .ZN(n132) );
  NOR2_X1 U257 ( .A1(A[15]), .A2(B[15]), .ZN(n94) );
  NOR2_X1 U258 ( .A1(A[13]), .A2(B[13]), .ZN(n114) );
  NOR2_X1 U259 ( .A1(A[6]), .A2(B[6]), .ZN(n164) );
  NOR2_X1 U260 ( .A1(A[2]), .A2(B[2]), .ZN(n183) );
  NOR2_X1 U261 ( .A1(A[16]), .A2(B[16]), .ZN(n85) );
  NOR2_X1 U262 ( .A1(A[8]), .A2(B[8]), .ZN(n153) );
  NOR2_X1 U263 ( .A1(A[1]), .A2(B[1]), .ZN(n187) );
  NOR2_X1 U264 ( .A1(A[22]), .A2(B[22]), .ZN(n37) );
  OR2_X1 U265 ( .A1(A[0]), .A2(B[0]), .ZN(n294) );
  NAND2_X1 U266 ( .A1(n126), .A2(n108), .ZN(n106) );
  INV_X1 U267 ( .A(n126), .ZN(n124) );
  INV_X1 U268 ( .A(n58), .ZN(n56) );
  AOI21_X1 U269 ( .B1(n127), .B2(n108), .A(n109), .ZN(n107) );
  INV_X1 U270 ( .A(n111), .ZN(n109) );
  INV_X1 U271 ( .A(n128), .ZN(n126) );
  INV_X1 U272 ( .A(n60), .ZN(n58) );
  INV_X1 U273 ( .A(n110), .ZN(n108) );
  NAND2_X1 U274 ( .A1(n99), .A2(n126), .ZN(n97) );
  NAND2_X1 U275 ( .A1(n58), .A2(n42), .ZN(n40) );
  INV_X1 U276 ( .A(n127), .ZN(n125) );
  INV_X1 U277 ( .A(n59), .ZN(n57) );
  OR2_X1 U278 ( .A1(n60), .A2(n33), .ZN(n295) );
  INV_X1 U279 ( .A(n148), .ZN(n142) );
  INV_X1 U280 ( .A(n76), .ZN(n74) );
  INV_X1 U281 ( .A(n77), .ZN(n75) );
  INV_X1 U282 ( .A(n145), .ZN(n143) );
  AOI21_X1 U283 ( .B1(n176), .B2(n167), .A(n168), .ZN(n166) );
  NOR2_X1 U284 ( .A1(n110), .A2(n101), .ZN(n99) );
  BUF_X1 U285 ( .A(n87), .Z(n1) );
  AOI21_X1 U286 ( .B1(n156), .B2(n88), .A(n89), .ZN(n87) );
  NOR2_X1 U287 ( .A1(n128), .A2(n90), .ZN(n88) );
  OAI21_X1 U288 ( .B1(n129), .B2(n90), .A(n91), .ZN(n89) );
  AOI21_X1 U289 ( .B1(n59), .B2(n42), .A(n45), .ZN(n41) );
  INV_X1 U290 ( .A(n129), .ZN(n127) );
  NAND2_X1 U291 ( .A1(n148), .A2(n130), .ZN(n128) );
  INV_X1 U292 ( .A(n61), .ZN(n59) );
  NAND2_X1 U293 ( .A1(n112), .A2(n92), .ZN(n90) );
  NAND2_X1 U294 ( .A1(n80), .A2(n62), .ZN(n60) );
  NAND2_X1 U295 ( .A1(n44), .A2(n35), .ZN(n33) );
  INV_X1 U296 ( .A(n177), .ZN(n176) );
  INV_X1 U297 ( .A(n113), .ZN(n111) );
  INV_X1 U298 ( .A(n112), .ZN(n110) );
  INV_X1 U299 ( .A(n186), .ZN(n185) );
  INV_X1 U300 ( .A(n147), .ZN(n145) );
  INV_X1 U301 ( .A(n149), .ZN(n147) );
  INV_X1 U302 ( .A(n43), .ZN(n42) );
  INV_X1 U303 ( .A(n44), .ZN(n43) );
  INV_X1 U304 ( .A(n79), .ZN(n77) );
  INV_X1 U305 ( .A(n81), .ZN(n79) );
  INV_X1 U306 ( .A(n78), .ZN(n76) );
  INV_X1 U307 ( .A(n80), .ZN(n78) );
  NAND2_X1 U308 ( .A1(n126), .A2(n119), .ZN(n117) );
  NAND2_X1 U309 ( .A1(n148), .A2(n137), .ZN(n135) );
  NAND2_X1 U310 ( .A1(n58), .A2(n51), .ZN(n49) );
  NAND2_X1 U311 ( .A1(n76), .A2(n69), .ZN(n67) );
  XOR2_X1 U312 ( .A(n1), .B(n9), .Z(SUM[16]) );
  NAND2_X1 U313 ( .A1(n198), .A2(n86), .ZN(n9) );
  INV_X1 U314 ( .A(n85), .ZN(n198) );
  XOR2_X1 U315 ( .A(n155), .B(n17), .Z(SUM[8]) );
  NAND2_X1 U316 ( .A1(n206), .A2(n154), .ZN(n17) );
  INV_X1 U317 ( .A(n153), .ZN(n206) );
  XOR2_X1 U318 ( .A(n166), .B(n19), .Z(SUM[6]) );
  NAND2_X1 U319 ( .A1(n208), .A2(n165), .ZN(n19) );
  INV_X1 U320 ( .A(n164), .ZN(n208) );
  XOR2_X1 U321 ( .A(n171), .B(n20), .Z(SUM[5]) );
  NAND2_X1 U322 ( .A1(n209), .A2(n170), .ZN(n20) );
  AOI21_X1 U323 ( .B1(n176), .B2(n172), .A(n173), .ZN(n171) );
  INV_X1 U324 ( .A(n169), .ZN(n209) );
  XOR2_X1 U325 ( .A(n24), .B(n190), .Z(SUM[1]) );
  NAND2_X1 U326 ( .A1(n213), .A2(n188), .ZN(n24) );
  INV_X1 U327 ( .A(n187), .ZN(n213) );
  OAI21_X1 U328 ( .B1(n150), .B2(n154), .A(n151), .ZN(n149) );
  XNOR2_X1 U329 ( .A(n163), .B(n18), .ZN(SUM[7]) );
  NAND2_X1 U330 ( .A1(n207), .A2(n162), .ZN(n18) );
  OAI21_X1 U331 ( .B1(n166), .B2(n164), .A(n165), .ZN(n163) );
  INV_X1 U332 ( .A(n161), .ZN(n207) );
  XNOR2_X1 U333 ( .A(n182), .B(n22), .ZN(SUM[3]) );
  OAI21_X1 U334 ( .B1(n185), .B2(n183), .A(n184), .ZN(n182) );
  NAND2_X1 U335 ( .A1(n211), .A2(n181), .ZN(n22) );
  INV_X1 U336 ( .A(n180), .ZN(n211) );
  XNOR2_X1 U337 ( .A(n73), .B(n7), .ZN(SUM[18]) );
  NAND2_X1 U338 ( .A1(n69), .A2(n72), .ZN(n7) );
  OAI21_X1 U339 ( .B1(n1), .B2(n74), .A(n75), .ZN(n73) );
  XNOR2_X1 U340 ( .A(n105), .B(n11), .ZN(SUM[14]) );
  NAND2_X1 U341 ( .A1(n102), .A2(n104), .ZN(n11) );
  OAI21_X1 U342 ( .B1(n155), .B2(n106), .A(n107), .ZN(n105) );
  XNOR2_X1 U343 ( .A(n116), .B(n12), .ZN(SUM[13]) );
  NAND2_X1 U344 ( .A1(n201), .A2(n115), .ZN(n12) );
  OAI21_X1 U345 ( .B1(n155), .B2(n117), .A(n118), .ZN(n116) );
  INV_X1 U346 ( .A(n114), .ZN(n201) );
  XNOR2_X1 U347 ( .A(n141), .B(n15), .ZN(SUM[10]) );
  NAND2_X1 U348 ( .A1(n137), .A2(n140), .ZN(n15) );
  OAI21_X1 U349 ( .B1(n155), .B2(n142), .A(n143), .ZN(n141) );
  XNOR2_X1 U350 ( .A(n48), .B(n4), .ZN(SUM[21]) );
  NAND2_X1 U351 ( .A1(n193), .A2(n47), .ZN(n4) );
  OAI21_X1 U352 ( .B1(n1), .B2(n49), .A(n50), .ZN(n48) );
  INV_X1 U353 ( .A(n46), .ZN(n193) );
  XNOR2_X1 U354 ( .A(n66), .B(n6), .ZN(SUM[19]) );
  NAND2_X1 U355 ( .A1(n195), .A2(n65), .ZN(n6) );
  OAI21_X1 U356 ( .B1(n1), .B2(n67), .A(n68), .ZN(n66) );
  INV_X1 U357 ( .A(n64), .ZN(n195) );
  XNOR2_X1 U358 ( .A(n176), .B(n21), .ZN(SUM[4]) );
  NAND2_X1 U359 ( .A1(n172), .A2(n175), .ZN(n21) );
  NOR2_X1 U360 ( .A1(n153), .A2(n150), .ZN(n148) );
  XNOR2_X1 U361 ( .A(n123), .B(n13), .ZN(SUM[12]) );
  NAND2_X1 U362 ( .A1(n119), .A2(n122), .ZN(n13) );
  OAI21_X1 U363 ( .B1(n155), .B2(n124), .A(n125), .ZN(n123) );
  XNOR2_X1 U364 ( .A(n55), .B(n5), .ZN(SUM[20]) );
  NAND2_X1 U365 ( .A1(n51), .A2(n54), .ZN(n5) );
  OAI21_X1 U366 ( .B1(n1), .B2(n56), .A(n57), .ZN(n55) );
  XNOR2_X1 U367 ( .A(n134), .B(n14), .ZN(SUM[11]) );
  NAND2_X1 U368 ( .A1(n203), .A2(n133), .ZN(n14) );
  OAI21_X1 U369 ( .B1(n155), .B2(n135), .A(n136), .ZN(n134) );
  INV_X1 U370 ( .A(n132), .ZN(n203) );
  XNOR2_X1 U371 ( .A(n96), .B(n10), .ZN(SUM[15]) );
  NAND2_X1 U372 ( .A1(n199), .A2(n95), .ZN(n10) );
  OAI21_X1 U373 ( .B1(n155), .B2(n97), .A(n98), .ZN(n96) );
  INV_X1 U374 ( .A(n94), .ZN(n199) );
  XNOR2_X1 U375 ( .A(n84), .B(n8), .ZN(SUM[17]) );
  NAND2_X1 U376 ( .A1(n197), .A2(n83), .ZN(n8) );
  OAI21_X1 U377 ( .B1(n1), .B2(n85), .A(n86), .ZN(n84) );
  INV_X1 U378 ( .A(n82), .ZN(n197) );
  XNOR2_X1 U379 ( .A(n152), .B(n16), .ZN(SUM[9]) );
  NAND2_X1 U380 ( .A1(n205), .A2(n151), .ZN(n16) );
  OAI21_X1 U381 ( .B1(n155), .B2(n153), .A(n154), .ZN(n152) );
  XNOR2_X1 U382 ( .A(n39), .B(n3), .ZN(SUM[22]) );
  NAND2_X1 U383 ( .A1(n192), .A2(n38), .ZN(n3) );
  OAI21_X1 U384 ( .B1(n1), .B2(n40), .A(n41), .ZN(n39) );
  INV_X1 U385 ( .A(n37), .ZN(n192) );
  AOI21_X1 U386 ( .B1(n62), .B2(n81), .A(n63), .ZN(n61) );
  OAI21_X1 U387 ( .B1(n64), .B2(n72), .A(n65), .ZN(n63) );
  AOI21_X1 U388 ( .B1(n130), .B2(n149), .A(n131), .ZN(n129) );
  OAI21_X1 U389 ( .B1(n132), .B2(n140), .A(n133), .ZN(n131) );
  AOI21_X1 U390 ( .B1(n178), .B2(n186), .A(n179), .ZN(n177) );
  NOR2_X1 U391 ( .A1(n183), .A2(n180), .ZN(n178) );
  OAI21_X1 U392 ( .B1(n180), .B2(n184), .A(n181), .ZN(n179) );
  OAI21_X1 U393 ( .B1(n114), .B2(n122), .A(n115), .ZN(n113) );
  OAI21_X1 U394 ( .B1(n82), .B2(n86), .A(n83), .ZN(n81) );
  OAI21_X1 U395 ( .B1(n187), .B2(n190), .A(n188), .ZN(n186) );
  OAI21_X1 U396 ( .B1(n169), .B2(n175), .A(n170), .ZN(n168) );
  OAI21_X1 U397 ( .B1(n46), .B2(n54), .A(n47), .ZN(n45) );
  NOR2_X1 U398 ( .A1(n174), .A2(n169), .ZN(n167) );
  NOR2_X1 U399 ( .A1(n139), .A2(n132), .ZN(n130) );
  NOR2_X1 U400 ( .A1(n71), .A2(n64), .ZN(n62) );
  NOR2_X1 U401 ( .A1(n103), .A2(n94), .ZN(n92) );
  NOR2_X1 U402 ( .A1(n85), .A2(n82), .ZN(n80) );
  NOR2_X1 U403 ( .A1(n121), .A2(n114), .ZN(n112) );
  NOR2_X1 U404 ( .A1(n53), .A2(n46), .ZN(n44) );
  OAI21_X1 U405 ( .B1(n177), .B2(n157), .A(n158), .ZN(n156) );
  NAND2_X1 U406 ( .A1(n167), .A2(n159), .ZN(n157) );
  AOI21_X1 U407 ( .B1(n159), .B2(n168), .A(n160), .ZN(n158) );
  NOR2_X1 U408 ( .A1(n164), .A2(n161), .ZN(n159) );
  AOI21_X1 U409 ( .B1(n92), .B2(n113), .A(n93), .ZN(n91) );
  OAI21_X1 U410 ( .B1(n94), .B2(n104), .A(n95), .ZN(n93) );
  AOI21_X1 U411 ( .B1(n99), .B2(n127), .A(n100), .ZN(n98) );
  OAI21_X1 U412 ( .B1(n111), .B2(n101), .A(n104), .ZN(n100) );
  AOI21_X1 U413 ( .B1(n127), .B2(n119), .A(n120), .ZN(n118) );
  INV_X1 U414 ( .A(n122), .ZN(n120) );
  AOI21_X1 U415 ( .B1(n145), .B2(n137), .A(n138), .ZN(n136) );
  INV_X1 U416 ( .A(n140), .ZN(n138) );
  AOI21_X1 U417 ( .B1(n59), .B2(n51), .A(n52), .ZN(n50) );
  INV_X1 U418 ( .A(n54), .ZN(n52) );
  AOI21_X1 U419 ( .B1(n77), .B2(n69), .A(n70), .ZN(n68) );
  INV_X1 U420 ( .A(n72), .ZN(n70) );
  OAI21_X1 U421 ( .B1(n161), .B2(n165), .A(n162), .ZN(n160) );
  INV_X1 U422 ( .A(n121), .ZN(n119) );
  INV_X1 U423 ( .A(n139), .ZN(n137) );
  INV_X1 U424 ( .A(n53), .ZN(n51) );
  INV_X1 U425 ( .A(n71), .ZN(n69) );
  INV_X1 U426 ( .A(n37), .ZN(n35) );
  INV_X1 U427 ( .A(n174), .ZN(n172) );
  INV_X1 U428 ( .A(n102), .ZN(n101) );
  INV_X1 U429 ( .A(n103), .ZN(n102) );
  XOR2_X1 U430 ( .A(n185), .B(n23), .Z(SUM[2]) );
  NAND2_X1 U431 ( .A1(n212), .A2(n184), .ZN(n23) );
  INV_X1 U432 ( .A(n183), .ZN(n212) );
  INV_X1 U433 ( .A(n175), .ZN(n173) );
  INV_X1 U434 ( .A(n32), .ZN(n30) );
  OAI21_X1 U435 ( .B1(n61), .B2(n33), .A(n34), .ZN(n32) );
  AOI21_X1 U436 ( .B1(n45), .B2(n35), .A(n36), .ZN(n34) );
  INV_X1 U437 ( .A(n38), .ZN(n36) );
  XNOR2_X1 U438 ( .A(n28), .B(n2), .ZN(SUM[23]) );
  NAND2_X1 U439 ( .A1(n296), .A2(n27), .ZN(n2) );
  OAI21_X1 U440 ( .B1(n1), .B2(n295), .A(n30), .ZN(n28) );
  NAND2_X1 U441 ( .A1(A[23]), .A2(B[23]), .ZN(n27) );
  NOR2_X1 U442 ( .A1(A[9]), .A2(B[9]), .ZN(n150) );
  NAND2_X1 U443 ( .A1(A[10]), .A2(B[10]), .ZN(n140) );
  NAND2_X1 U444 ( .A1(A[4]), .A2(B[4]), .ZN(n175) );
  NAND2_X1 U445 ( .A1(A[12]), .A2(B[12]), .ZN(n122) );
  NAND2_X1 U446 ( .A1(A[18]), .A2(B[18]), .ZN(n72) );
  NAND2_X1 U447 ( .A1(A[20]), .A2(B[20]), .ZN(n54) );
  NAND2_X1 U448 ( .A1(A[2]), .A2(B[2]), .ZN(n184) );
  NAND2_X1 U449 ( .A1(A[6]), .A2(B[6]), .ZN(n165) );
  NAND2_X1 U450 ( .A1(A[16]), .A2(B[16]), .ZN(n86) );
  NAND2_X1 U451 ( .A1(A[14]), .A2(B[14]), .ZN(n104) );
  NAND2_X1 U452 ( .A1(A[0]), .A2(B[0]), .ZN(n190) );
  NAND2_X1 U453 ( .A1(A[8]), .A2(B[8]), .ZN(n154) );
  NAND2_X1 U454 ( .A1(A[22]), .A2(B[22]), .ZN(n38) );
  NAND2_X1 U455 ( .A1(A[11]), .A2(B[11]), .ZN(n133) );
  NAND2_X1 U456 ( .A1(A[1]), .A2(B[1]), .ZN(n188) );
  NAND2_X1 U457 ( .A1(A[3]), .A2(B[3]), .ZN(n181) );
  NAND2_X1 U458 ( .A1(A[5]), .A2(B[5]), .ZN(n170) );
  NAND2_X1 U459 ( .A1(A[7]), .A2(B[7]), .ZN(n162) );
  NAND2_X1 U460 ( .A1(A[13]), .A2(B[13]), .ZN(n115) );
  NAND2_X1 U461 ( .A1(A[17]), .A2(B[17]), .ZN(n83) );
  NAND2_X1 U462 ( .A1(A[19]), .A2(B[19]), .ZN(n65) );
  NAND2_X1 U463 ( .A1(A[21]), .A2(B[21]), .ZN(n47) );
  NAND2_X1 U464 ( .A1(A[15]), .A2(B[15]), .ZN(n95) );
  NAND2_X1 U465 ( .A1(A[9]), .A2(B[9]), .ZN(n151) );
  OR2_X1 U466 ( .A1(A[23]), .A2(B[23]), .ZN(n296) );
  INV_X1 U467 ( .A(n150), .ZN(n205) );
endmodule


module iir_filter_DW01_add_5 ( A, B, SUM, CI, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n27, n28, n30, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n77,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n145, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n190, n192, n193, n195, n197, n198, n199, n201,
         n203, n205, n206, n207, n208, n209, n211, n212, n213, n294, n295,
         n296, n297;

  NOR2_X2 U242 ( .A1(A[3]), .A2(B[3]), .ZN(n180) );
  AOI21_X1 U243 ( .B1(n178), .B2(n186), .A(n179), .ZN(n177) );
  AND2_X1 U244 ( .A1(n295), .A2(n190), .ZN(SUM[0]) );
  OAI21_X1 U245 ( .B1(n177), .B2(n157), .A(n158), .ZN(n294) );
  INV_X2 U246 ( .A(n294), .ZN(n155) );
  NOR2_X1 U247 ( .A1(A[4]), .A2(B[4]), .ZN(n174) );
  NOR2_X1 U248 ( .A1(A[20]), .A2(B[20]), .ZN(n53) );
  NOR2_X1 U249 ( .A1(A[18]), .A2(B[18]), .ZN(n71) );
  NOR2_X1 U250 ( .A1(A[10]), .A2(B[10]), .ZN(n139) );
  NOR2_X1 U251 ( .A1(A[14]), .A2(B[14]), .ZN(n103) );
  NOR2_X1 U252 ( .A1(A[12]), .A2(B[12]), .ZN(n121) );
  NOR2_X1 U253 ( .A1(A[7]), .A2(B[7]), .ZN(n161) );
  NOR2_X1 U254 ( .A1(A[21]), .A2(B[21]), .ZN(n46) );
  NOR2_X1 U255 ( .A1(A[19]), .A2(B[19]), .ZN(n64) );
  NOR2_X1 U256 ( .A1(A[17]), .A2(B[17]), .ZN(n82) );
  NOR2_X1 U257 ( .A1(A[15]), .A2(B[15]), .ZN(n94) );
  NOR2_X1 U258 ( .A1(A[6]), .A2(B[6]), .ZN(n164) );
  NOR2_X1 U259 ( .A1(A[2]), .A2(B[2]), .ZN(n183) );
  NOR2_X1 U260 ( .A1(A[16]), .A2(B[16]), .ZN(n85) );
  NOR2_X1 U261 ( .A1(A[8]), .A2(B[8]), .ZN(n153) );
  NOR2_X1 U262 ( .A1(A[1]), .A2(B[1]), .ZN(n187) );
  NOR2_X1 U263 ( .A1(A[22]), .A2(B[22]), .ZN(n37) );
  OR2_X1 U264 ( .A1(A[0]), .A2(B[0]), .ZN(n295) );
  NAND2_X1 U265 ( .A1(n126), .A2(n108), .ZN(n106) );
  INV_X1 U266 ( .A(n126), .ZN(n124) );
  INV_X1 U267 ( .A(n58), .ZN(n56) );
  AOI21_X1 U268 ( .B1(n127), .B2(n108), .A(n109), .ZN(n107) );
  INV_X1 U269 ( .A(n111), .ZN(n109) );
  INV_X1 U270 ( .A(n128), .ZN(n126) );
  INV_X1 U271 ( .A(n60), .ZN(n58) );
  INV_X1 U272 ( .A(n110), .ZN(n108) );
  NAND2_X1 U273 ( .A1(n99), .A2(n126), .ZN(n97) );
  NAND2_X1 U274 ( .A1(n58), .A2(n42), .ZN(n40) );
  INV_X1 U275 ( .A(n127), .ZN(n125) );
  INV_X1 U276 ( .A(n59), .ZN(n57) );
  OR2_X1 U277 ( .A1(n60), .A2(n33), .ZN(n296) );
  INV_X1 U278 ( .A(n148), .ZN(n142) );
  INV_X1 U279 ( .A(n80), .ZN(n74) );
  INV_X1 U280 ( .A(n145), .ZN(n143) );
  INV_X1 U281 ( .A(n77), .ZN(n75) );
  BUF_X1 U282 ( .A(n87), .Z(n1) );
  NOR2_X1 U283 ( .A1(n128), .A2(n90), .ZN(n88) );
  OAI21_X1 U284 ( .B1(n129), .B2(n90), .A(n91), .ZN(n89) );
  AOI21_X1 U285 ( .B1(n176), .B2(n167), .A(n168), .ZN(n166) );
  NOR2_X1 U286 ( .A1(n110), .A2(n101), .ZN(n99) );
  AOI21_X1 U287 ( .B1(n59), .B2(n42), .A(n45), .ZN(n41) );
  NAND2_X1 U288 ( .A1(n112), .A2(n92), .ZN(n90) );
  NAND2_X1 U289 ( .A1(n148), .A2(n130), .ZN(n128) );
  INV_X1 U290 ( .A(n129), .ZN(n127) );
  INV_X1 U291 ( .A(n113), .ZN(n111) );
  INV_X1 U292 ( .A(n112), .ZN(n110) );
  INV_X1 U293 ( .A(n61), .ZN(n59) );
  NAND2_X1 U294 ( .A1(n80), .A2(n62), .ZN(n60) );
  NAND2_X1 U295 ( .A1(n44), .A2(n35), .ZN(n33) );
  INV_X1 U296 ( .A(n177), .ZN(n176) );
  INV_X1 U297 ( .A(n186), .ZN(n185) );
  INV_X1 U298 ( .A(n147), .ZN(n145) );
  INV_X1 U299 ( .A(n149), .ZN(n147) );
  INV_X1 U300 ( .A(n43), .ZN(n42) );
  INV_X1 U301 ( .A(n44), .ZN(n43) );
  INV_X1 U302 ( .A(n79), .ZN(n77) );
  INV_X1 U303 ( .A(n81), .ZN(n79) );
  NAND2_X1 U304 ( .A1(n58), .A2(n51), .ZN(n49) );
  NAND2_X1 U305 ( .A1(n80), .A2(n69), .ZN(n67) );
  NAND2_X1 U306 ( .A1(n126), .A2(n119), .ZN(n117) );
  NAND2_X1 U307 ( .A1(n148), .A2(n137), .ZN(n135) );
  XOR2_X1 U308 ( .A(n1), .B(n9), .Z(SUM[16]) );
  NAND2_X1 U309 ( .A1(n198), .A2(n86), .ZN(n9) );
  INV_X1 U310 ( .A(n85), .ZN(n198) );
  XOR2_X1 U311 ( .A(n155), .B(n17), .Z(SUM[8]) );
  NAND2_X1 U312 ( .A1(n206), .A2(n154), .ZN(n17) );
  INV_X1 U313 ( .A(n153), .ZN(n206) );
  XOR2_X1 U314 ( .A(n166), .B(n19), .Z(SUM[6]) );
  NAND2_X1 U315 ( .A1(n208), .A2(n165), .ZN(n19) );
  INV_X1 U316 ( .A(n164), .ZN(n208) );
  XOR2_X1 U317 ( .A(n185), .B(n23), .Z(SUM[2]) );
  NAND2_X1 U318 ( .A1(n212), .A2(n184), .ZN(n23) );
  INV_X1 U319 ( .A(n183), .ZN(n212) );
  XOR2_X1 U320 ( .A(n171), .B(n20), .Z(SUM[5]) );
  NAND2_X1 U321 ( .A1(n209), .A2(n170), .ZN(n20) );
  AOI21_X1 U322 ( .B1(n176), .B2(n172), .A(n173), .ZN(n171) );
  XNOR2_X1 U323 ( .A(n163), .B(n18), .ZN(SUM[7]) );
  NAND2_X1 U324 ( .A1(n207), .A2(n162), .ZN(n18) );
  OAI21_X1 U325 ( .B1(n166), .B2(n164), .A(n165), .ZN(n163) );
  INV_X1 U326 ( .A(n161), .ZN(n207) );
  XNOR2_X1 U327 ( .A(n73), .B(n7), .ZN(SUM[18]) );
  NAND2_X1 U328 ( .A1(n69), .A2(n72), .ZN(n7) );
  OAI21_X1 U329 ( .B1(n1), .B2(n74), .A(n75), .ZN(n73) );
  XNOR2_X1 U330 ( .A(n48), .B(n4), .ZN(SUM[21]) );
  NAND2_X1 U331 ( .A1(n193), .A2(n47), .ZN(n4) );
  OAI21_X1 U332 ( .B1(n1), .B2(n49), .A(n50), .ZN(n48) );
  INV_X1 U333 ( .A(n46), .ZN(n193) );
  XNOR2_X1 U334 ( .A(n66), .B(n6), .ZN(SUM[19]) );
  NAND2_X1 U335 ( .A1(n195), .A2(n65), .ZN(n6) );
  OAI21_X1 U336 ( .B1(n1), .B2(n67), .A(n68), .ZN(n66) );
  INV_X1 U337 ( .A(n64), .ZN(n195) );
  XNOR2_X1 U338 ( .A(n105), .B(n11), .ZN(SUM[14]) );
  NAND2_X1 U339 ( .A1(n102), .A2(n104), .ZN(n11) );
  OAI21_X1 U340 ( .B1(n155), .B2(n106), .A(n107), .ZN(n105) );
  XNOR2_X1 U341 ( .A(n116), .B(n12), .ZN(SUM[13]) );
  NAND2_X1 U342 ( .A1(n201), .A2(n115), .ZN(n12) );
  OAI21_X1 U343 ( .B1(n155), .B2(n117), .A(n118), .ZN(n116) );
  INV_X1 U344 ( .A(n114), .ZN(n201) );
  XNOR2_X1 U345 ( .A(n141), .B(n15), .ZN(SUM[10]) );
  NAND2_X1 U346 ( .A1(n137), .A2(n140), .ZN(n15) );
  OAI21_X1 U347 ( .B1(n155), .B2(n142), .A(n143), .ZN(n141) );
  XNOR2_X1 U348 ( .A(n176), .B(n21), .ZN(SUM[4]) );
  NAND2_X1 U349 ( .A1(n172), .A2(n175), .ZN(n21) );
  OAI21_X1 U350 ( .B1(n150), .B2(n154), .A(n151), .ZN(n149) );
  OAI21_X1 U351 ( .B1(n169), .B2(n175), .A(n170), .ZN(n168) );
  NOR2_X1 U352 ( .A1(n174), .A2(n169), .ZN(n167) );
  XNOR2_X1 U353 ( .A(n123), .B(n13), .ZN(SUM[12]) );
  NAND2_X1 U354 ( .A1(n119), .A2(n122), .ZN(n13) );
  OAI21_X1 U355 ( .B1(n155), .B2(n124), .A(n125), .ZN(n123) );
  XNOR2_X1 U356 ( .A(n55), .B(n5), .ZN(SUM[20]) );
  NAND2_X1 U357 ( .A1(n51), .A2(n54), .ZN(n5) );
  OAI21_X1 U358 ( .B1(n1), .B2(n56), .A(n57), .ZN(n55) );
  XNOR2_X1 U359 ( .A(n134), .B(n14), .ZN(SUM[11]) );
  NAND2_X1 U360 ( .A1(n203), .A2(n133), .ZN(n14) );
  OAI21_X1 U361 ( .B1(n155), .B2(n135), .A(n136), .ZN(n134) );
  XNOR2_X1 U362 ( .A(n96), .B(n10), .ZN(SUM[15]) );
  NAND2_X1 U363 ( .A1(n199), .A2(n95), .ZN(n10) );
  OAI21_X1 U364 ( .B1(n155), .B2(n97), .A(n98), .ZN(n96) );
  INV_X1 U365 ( .A(n94), .ZN(n199) );
  XNOR2_X1 U366 ( .A(n84), .B(n8), .ZN(SUM[17]) );
  NAND2_X1 U367 ( .A1(n197), .A2(n83), .ZN(n8) );
  OAI21_X1 U368 ( .B1(n1), .B2(n85), .A(n86), .ZN(n84) );
  INV_X1 U369 ( .A(n82), .ZN(n197) );
  XNOR2_X1 U370 ( .A(n152), .B(n16), .ZN(SUM[9]) );
  NAND2_X1 U371 ( .A1(n205), .A2(n151), .ZN(n16) );
  OAI21_X1 U372 ( .B1(n155), .B2(n153), .A(n154), .ZN(n152) );
  XNOR2_X1 U373 ( .A(n39), .B(n3), .ZN(SUM[22]) );
  NAND2_X1 U374 ( .A1(n192), .A2(n38), .ZN(n3) );
  OAI21_X1 U375 ( .B1(n1), .B2(n40), .A(n41), .ZN(n39) );
  INV_X1 U376 ( .A(n37), .ZN(n192) );
  AOI21_X1 U377 ( .B1(n130), .B2(n149), .A(n131), .ZN(n129) );
  NOR2_X1 U378 ( .A1(n183), .A2(n180), .ZN(n178) );
  AOI21_X1 U379 ( .B1(n62), .B2(n81), .A(n63), .ZN(n61) );
  OAI21_X1 U380 ( .B1(n64), .B2(n72), .A(n65), .ZN(n63) );
  OAI21_X1 U381 ( .B1(n82), .B2(n86), .A(n83), .ZN(n81) );
  OAI21_X1 U382 ( .B1(n187), .B2(n190), .A(n188), .ZN(n186) );
  OAI21_X1 U383 ( .B1(n46), .B2(n54), .A(n47), .ZN(n45) );
  NOR2_X1 U384 ( .A1(n71), .A2(n64), .ZN(n62) );
  NOR2_X1 U385 ( .A1(n103), .A2(n94), .ZN(n92) );
  AOI21_X1 U386 ( .B1(n92), .B2(n113), .A(n93), .ZN(n91) );
  OAI21_X1 U387 ( .B1(n94), .B2(n104), .A(n95), .ZN(n93) );
  NOR2_X1 U388 ( .A1(n85), .A2(n82), .ZN(n80) );
  NOR2_X1 U389 ( .A1(n53), .A2(n46), .ZN(n44) );
  AOI21_X1 U390 ( .B1(n99), .B2(n127), .A(n100), .ZN(n98) );
  OAI21_X1 U391 ( .B1(n111), .B2(n101), .A(n104), .ZN(n100) );
  AOI21_X1 U392 ( .B1(n127), .B2(n119), .A(n120), .ZN(n118) );
  INV_X1 U393 ( .A(n122), .ZN(n120) );
  AOI21_X1 U394 ( .B1(n145), .B2(n137), .A(n138), .ZN(n136) );
  INV_X1 U395 ( .A(n140), .ZN(n138) );
  AOI21_X1 U396 ( .B1(n59), .B2(n51), .A(n52), .ZN(n50) );
  INV_X1 U397 ( .A(n54), .ZN(n52) );
  AOI21_X1 U398 ( .B1(n77), .B2(n69), .A(n70), .ZN(n68) );
  INV_X1 U399 ( .A(n72), .ZN(n70) );
  NAND2_X1 U400 ( .A1(n167), .A2(n159), .ZN(n157) );
  AOI21_X1 U401 ( .B1(n159), .B2(n168), .A(n160), .ZN(n158) );
  NOR2_X1 U402 ( .A1(n164), .A2(n161), .ZN(n159) );
  OAI21_X1 U403 ( .B1(n161), .B2(n165), .A(n162), .ZN(n160) );
  INV_X1 U404 ( .A(n53), .ZN(n51) );
  INV_X1 U405 ( .A(n71), .ZN(n69) );
  INV_X1 U406 ( .A(n121), .ZN(n119) );
  INV_X1 U407 ( .A(n139), .ZN(n137) );
  INV_X1 U408 ( .A(n37), .ZN(n35) );
  INV_X1 U409 ( .A(n174), .ZN(n172) );
  INV_X1 U410 ( .A(n102), .ZN(n101) );
  INV_X1 U411 ( .A(n103), .ZN(n102) );
  XNOR2_X1 U412 ( .A(n182), .B(n22), .ZN(SUM[3]) );
  OAI21_X1 U413 ( .B1(n185), .B2(n183), .A(n184), .ZN(n182) );
  NAND2_X1 U414 ( .A1(n211), .A2(n181), .ZN(n22) );
  INV_X1 U415 ( .A(n180), .ZN(n211) );
  XOR2_X1 U416 ( .A(n24), .B(n190), .Z(SUM[1]) );
  NAND2_X1 U417 ( .A1(n213), .A2(n188), .ZN(n24) );
  INV_X1 U418 ( .A(n187), .ZN(n213) );
  INV_X1 U419 ( .A(n175), .ZN(n173) );
  INV_X1 U420 ( .A(n32), .ZN(n30) );
  OAI21_X1 U421 ( .B1(n61), .B2(n33), .A(n34), .ZN(n32) );
  AOI21_X1 U422 ( .B1(n45), .B2(n35), .A(n36), .ZN(n34) );
  INV_X1 U423 ( .A(n38), .ZN(n36) );
  XNOR2_X1 U424 ( .A(n28), .B(n2), .ZN(SUM[23]) );
  NAND2_X1 U425 ( .A1(n297), .A2(n27), .ZN(n2) );
  OAI21_X1 U426 ( .B1(n1), .B2(n296), .A(n30), .ZN(n28) );
  NAND2_X1 U427 ( .A1(A[23]), .A2(B[23]), .ZN(n27) );
  NOR2_X1 U428 ( .A1(A[5]), .A2(B[5]), .ZN(n169) );
  NOR2_X1 U429 ( .A1(A[13]), .A2(B[13]), .ZN(n114) );
  NAND2_X1 U430 ( .A1(A[18]), .A2(B[18]), .ZN(n72) );
  NAND2_X1 U431 ( .A1(A[6]), .A2(B[6]), .ZN(n165) );
  NAND2_X1 U432 ( .A1(A[16]), .A2(B[16]), .ZN(n86) );
  NAND2_X1 U433 ( .A1(A[14]), .A2(B[14]), .ZN(n104) );
  NAND2_X1 U434 ( .A1(A[20]), .A2(B[20]), .ZN(n54) );
  NAND2_X1 U435 ( .A1(A[0]), .A2(B[0]), .ZN(n190) );
  NAND2_X1 U436 ( .A1(A[4]), .A2(B[4]), .ZN(n175) );
  NAND2_X1 U437 ( .A1(A[8]), .A2(B[8]), .ZN(n154) );
  NAND2_X1 U438 ( .A1(A[10]), .A2(B[10]), .ZN(n140) );
  NAND2_X1 U439 ( .A1(A[12]), .A2(B[12]), .ZN(n122) );
  NAND2_X1 U440 ( .A1(A[2]), .A2(B[2]), .ZN(n184) );
  NAND2_X1 U441 ( .A1(A[22]), .A2(B[22]), .ZN(n38) );
  NAND2_X1 U442 ( .A1(A[1]), .A2(B[1]), .ZN(n188) );
  NAND2_X1 U443 ( .A1(A[7]), .A2(B[7]), .ZN(n162) );
  NAND2_X1 U444 ( .A1(A[15]), .A2(B[15]), .ZN(n95) );
  NAND2_X1 U445 ( .A1(A[17]), .A2(B[17]), .ZN(n83) );
  NAND2_X1 U446 ( .A1(A[19]), .A2(B[19]), .ZN(n65) );
  NAND2_X1 U447 ( .A1(A[21]), .A2(B[21]), .ZN(n47) );
  NAND2_X1 U448 ( .A1(A[3]), .A2(B[3]), .ZN(n181) );
  NAND2_X1 U449 ( .A1(A[13]), .A2(B[13]), .ZN(n115) );
  NAND2_X1 U450 ( .A1(A[5]), .A2(B[5]), .ZN(n170) );
  NAND2_X1 U451 ( .A1(A[9]), .A2(B[9]), .ZN(n151) );
  NAND2_X1 U452 ( .A1(A[11]), .A2(B[11]), .ZN(n133) );
  OR2_X1 U453 ( .A1(A[23]), .A2(B[23]), .ZN(n297) );
  AOI21_X1 U454 ( .B1(n294), .B2(n88), .A(n89), .ZN(n87) );
  INV_X1 U455 ( .A(n169), .ZN(n209) );
  NOR2_X1 U456 ( .A1(n121), .A2(n114), .ZN(n112) );
  OAI21_X1 U457 ( .B1(n114), .B2(n122), .A(n115), .ZN(n113) );
  NOR2_X1 U458 ( .A1(A[11]), .A2(B[11]), .ZN(n132) );
  OAI21_X1 U459 ( .B1(n132), .B2(n140), .A(n133), .ZN(n131) );
  NOR2_X1 U460 ( .A1(n139), .A2(n132), .ZN(n130) );
  INV_X1 U461 ( .A(n132), .ZN(n203) );
  NOR2_X1 U462 ( .A1(A[9]), .A2(B[9]), .ZN(n150) );
  NOR2_X1 U463 ( .A1(n153), .A2(n150), .ZN(n148) );
  INV_X1 U464 ( .A(n150), .ZN(n205) );
  OAI21_X1 U465 ( .B1(n180), .B2(n184), .A(n181), .ZN(n179) );
endmodule


module iir_filter ( clk, rst_n, vIn, dIn, coeffs_fb, coeffs_ff, dOut, vOut );
  input [11:0] dIn;
  input [47:0] coeffs_fb;
  input [95:0] coeffs_ff;
  output [11:0] dOut;
  input clk, rst_n, vIn;
  output vOut;
  wire   delayed_controls_0__1_, delayed_controls_1__0_,
         delayed_controls_1__1_, delayed_controls_2__0_, DP_y_0_, DP_y_1_,
         DP_y_2_, DP_y_3_, DP_y_4_, DP_y_5_, DP_y_6_, DP_y_7_, DP_y_8_,
         DP_y_9_, DP_y_10_, DP_y_11_, DP_y_23, DP_sw1_0_, DP_sw1_1_, DP_sw1_2_,
         DP_sw1_3_, DP_sw1_4_, DP_sw1_5_, DP_sw1_6_, DP_sw1_7_, DP_sw1_8_,
         DP_sw1_9_, DP_sw1_10_, DP_sw1_11_, DP_sw1_12_, DP_sw1_13_, DP_sw1_14_,
         DP_sw1_15_, DP_sw1_16_, DP_sw1_17_, DP_sw1_18_, DP_sw1_19_,
         DP_sw1_20_, DP_sw1_21_, DP_sw1_22_, DP_sw1_23_, DP_sw0_0_, DP_sw0_1_,
         DP_sw0_2_, DP_sw0_3_, DP_sw0_4_, DP_sw0_5_, DP_sw0_6_, DP_sw0_7_,
         DP_sw0_8_, DP_sw0_9_, DP_sw0_10_, DP_sw0_11_, DP_sw0_12_, DP_sw0_13_,
         DP_sw0_14_, DP_sw0_15_, DP_sw0_16_, DP_sw0_17_, DP_sw0_18_,
         DP_sw0_19_, DP_sw0_20_, DP_sw0_21_, DP_sw0_22_, DP_sw0_23_, DP_w_0_,
         DP_w_1_, DP_w_2_, DP_w_3_, DP_w_4_, DP_w_5_, DP_w_6_, DP_w_7_,
         DP_w_8_, DP_w_9_, DP_w_10_, DP_w_11_, DP_w_12_, DP_w_13_, DP_w_14_,
         DP_w_15_, DP_w_16_, DP_w_17_, DP_w_18_, DP_w_19_, DP_w_20_, DP_w_21_,
         DP_w_22_, DP_w_23_, CU_nextState_0_, n280, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n529, n531, n533,
         n535, n537, n539, n541, n543, n545, n547, n549, n551, n553, n555,
         n557, n559, n561, n563, n565, n567, n569, n571, n573, n575, DP_fb_9_,
         DP_fb_8_, DP_fb_7_, DP_fb_6_, DP_fb_5_, DP_fb_4_, DP_fb_3_, DP_fb_2_,
         DP_fb_23_, DP_fb_22_, DP_fb_21_, DP_fb_20_, DP_fb_1_, DP_fb_19_,
         DP_fb_18_, DP_fb_17_, DP_fb_16_, DP_fb_15_, DP_fb_14_, DP_fb_13_,
         DP_fb_12_, DP_fb_11_, DP_fb_10_, DP_fb_0_, DP_ff_part_9_,
         DP_ff_part_8_, DP_ff_part_7_, DP_ff_part_6_, DP_ff_part_5_,
         DP_ff_part_4_, DP_ff_part_3_, DP_ff_part_2_, DP_ff_part_23_,
         DP_ff_part_22_, DP_ff_part_21_, DP_ff_part_20_, DP_ff_part_1_,
         DP_ff_part_19_, DP_ff_part_18_, DP_ff_part_17_, DP_ff_part_16_,
         DP_ff_part_15_, DP_ff_part_14_, DP_ff_part_13_, DP_ff_part_12_,
         DP_ff_part_11_, DP_ff_part_10_, DP_ff_part_0_, DP_ff_9_, DP_ff_8_,
         DP_ff_7_, DP_ff_6_, DP_ff_5_, DP_ff_4_, DP_ff_3_, DP_ff_2_, DP_ff_23_,
         DP_ff_22_, DP_ff_21_, DP_ff_20_, DP_ff_1_, DP_ff_19_, DP_ff_18_,
         DP_ff_17_, DP_ff_16_, DP_ff_15_, DP_ff_14_, DP_ff_13_, DP_ff_12_,
         DP_ff_11_, DP_ff_10_, DP_ff_0_, n997, n998, n1000, n1001, n1004,
         n1005, n1006, n1007, n1008, n1009, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1034, n1037, n1038, n1040, n1041, n1042, n1043, n1044, n1045,
         n1047, n1048, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1084, n1085, n1086, n1087, n1089, n1090, n1091, n1092,
         n1094, n1095, n1096, n1097, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1137,
         n1138, n1139, n1140, n1141, n1142, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471;
  wire   [0:23] DP_pipe13;
  wire   [0:23] DP_pipe0_coeff_pipe03;
  wire   [0:23] DP_pipe12;
  wire   [0:23] DP_pipe0_coeff_pipe02;
  wire   [0:23] DP_pipe11;
  wire   [0:23] DP_pipe0_coeff_pipe01;
  wire   [0:23] DP_pipe10;
  wire   [0:23] DP_pipe0_coeff_pipe00;
  wire   [0:23] DP_pipe03;
  wire   [0:23] DP_pipe02;
  wire   [0:23] DP_pipe01;
  wire   [0:23] DP_pipe00;
  wire   [0:23] DP_ret1;
  wire   [0:23] DP_sw1_coeff_ret1;
  wire   [0:23] DP_ret0;
  wire   [0:23] DP_sw0_coeff_ret0;
  wire   [95:0] DP_coeffs_ff_int;
  wire   [47:0] DP_coeffs_fb_int;
  wire   [0:11] DP_x;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154;

  DFFR_X1 DP_reg_in_Q_reg_0_ ( .D(n1268), .CK(clk), .RN(n1173), .Q(DP_x[0]) );
  DFFR_X1 DP_reg_in_Q_reg_1_ ( .D(n1269), .CK(clk), .RN(n1173), .Q(DP_x[1]) );
  DFFR_X1 DP_reg_in_Q_reg_2_ ( .D(n1270), .CK(clk), .RN(n1173), .Q(DP_x[2]) );
  DFFR_X1 DP_reg_in_Q_reg_3_ ( .D(n1271), .CK(clk), .RN(n1173), .Q(DP_x[3]) );
  DFFR_X1 DP_reg_in_Q_reg_4_ ( .D(n1272), .CK(clk), .RN(n1173), .Q(DP_x[4]) );
  DFFR_X1 DP_reg_in_Q_reg_5_ ( .D(n1273), .CK(clk), .RN(n1173), .Q(DP_x[5]) );
  DFFR_X1 DP_reg_in_Q_reg_6_ ( .D(n1274), .CK(clk), .RN(n1173), .Q(DP_x[6]) );
  DFFR_X1 DP_reg_in_Q_reg_7_ ( .D(n1275), .CK(clk), .RN(n1173), .Q(DP_x[7]) );
  DFFR_X1 DP_reg_in_Q_reg_8_ ( .D(n1276), .CK(clk), .RN(n1173), .Q(DP_x[8]) );
  DFFR_X1 DP_reg_in_Q_reg_9_ ( .D(n1277), .CK(clk), .RN(n1173), .Q(DP_x[9]) );
  DFFR_X1 DP_reg_in_Q_reg_10_ ( .D(n1278), .CK(clk), .RN(n1173), .Q(DP_x[10])
         );
  DFFR_X1 DP_reg_in_Q_reg_11_ ( .D(n1279), .CK(clk), .RN(n1173), .Q(DP_x[11])
         );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_0_ ( .D(n1280), .CK(clk), .RN(n1174), .Q(
        DP_coeffs_fb_int[23]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_1_ ( .D(n1281), .CK(clk), .RN(n1174), .Q(
        DP_coeffs_fb_int[22]), .QN(n1107) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_2_ ( .D(n1282), .CK(clk), .RN(n1174), .Q(
        DP_coeffs_fb_int[21]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_3_ ( .D(n1283), .CK(clk), .RN(n1174), .Q(
        DP_coeffs_fb_int[20]), .QN(n1078) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_4_ ( .D(n1284), .CK(clk), .RN(n1174), .Q(
        DP_coeffs_fb_int[19]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_5_ ( .D(n1285), .CK(clk), .RN(n1174), .Q(
        DP_coeffs_fb_int[18]), .QN(n1105) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_6_ ( .D(n1286), .CK(clk), .RN(n1174), .Q(
        DP_coeffs_fb_int[17]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_7_ ( .D(n1287), .CK(clk), .RN(n1174), .Q(
        DP_coeffs_fb_int[16]), .QN(n1042) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_8_ ( .D(n1288), .CK(clk), .RN(n1174), .Q(
        DP_coeffs_fb_int[15]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_9_ ( .D(n1289), .CK(clk), .RN(n1174), .Q(
        DP_coeffs_fb_int[14]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_10_ ( .D(n1290), .CK(clk), .RN(n1174), .Q(
        DP_coeffs_fb_int[13]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_11_ ( .D(n1291), .CK(clk), .RN(n1174), .Q(
        DP_coeffs_fb_int[12]), .QN(n1086) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_12_ ( .D(n1292), .CK(clk), .RN(n1175), .Q(
        DP_coeffs_fb_int[11]), .QN(n1062) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_13_ ( .D(n1293), .CK(clk), .RN(n1175), .Q(
        DP_coeffs_fb_int[10]), .QN(n1031) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_14_ ( .D(n1294), .CK(clk), .RN(n1175), .Q(
        DP_coeffs_fb_int[9]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_15_ ( .D(n1295), .CK(clk), .RN(n1175), .Q(
        DP_coeffs_fb_int[8]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_16_ ( .D(n1296), .CK(clk), .RN(n1175), .Q(
        DP_coeffs_fb_int[7]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_17_ ( .D(n1297), .CK(clk), .RN(n1175), .Q(
        DP_coeffs_fb_int[6]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_18_ ( .D(n1298), .CK(clk), .RN(n1175), .Q(
        DP_coeffs_fb_int[5]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_19_ ( .D(n1299), .CK(clk), .RN(n1175), .Q(
        DP_coeffs_fb_int[4]), .QN(n1089) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_20_ ( .D(n1300), .CK(clk), .RN(n1175), .Q(
        DP_coeffs_fb_int[3]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_21_ ( .D(n1301), .CK(clk), .RN(n1175), .Q(
        DP_coeffs_fb_int[2]), .QN(n1099) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_22_ ( .D(n1302), .CK(clk), .RN(n1175), .Q(
        DP_coeffs_fb_int[1]) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_23_ ( .D(n1303), .CK(clk), .RN(n1175), .Q(
        DP_coeffs_fb_int[0]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_0_ ( .D(n1304), .CK(clk), .RN(n1176), .Q(
        DP_coeffs_fb_int[47]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_1_ ( .D(n1305), .CK(clk), .RN(n1176), .Q(
        DP_coeffs_fb_int[46]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_2_ ( .D(n1306), .CK(clk), .RN(n1176), .Q(
        DP_coeffs_fb_int[45]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_3_ ( .D(n1307), .CK(clk), .RN(n1176), .Q(
        DP_coeffs_fb_int[44]), .QN(n1037) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_4_ ( .D(n1308), .CK(clk), .RN(n1176), .Q(
        DP_coeffs_fb_int[43]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_5_ ( .D(n1309), .CK(clk), .RN(n1176), .Q(
        DP_coeffs_fb_int[42]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_6_ ( .D(n1310), .CK(clk), .RN(n1176), .Q(
        DP_coeffs_fb_int[41]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_7_ ( .D(n1311), .CK(clk), .RN(n1176), .Q(
        DP_coeffs_fb_int[40]), .QN(n1084) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_8_ ( .D(n1312), .CK(clk), .RN(n1176), .Q(
        DP_coeffs_fb_int[39]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_9_ ( .D(n1313), .CK(clk), .RN(n1176), .Q(
        DP_coeffs_fb_int[38]), .QN(n1139) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_10_ ( .D(n1314), .CK(clk), .RN(n1176), .Q(
        DP_coeffs_fb_int[37]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_11_ ( .D(n1315), .CK(clk), .RN(n1176), .Q(
        DP_coeffs_fb_int[36]), .QN(n1004) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_12_ ( .D(n1316), .CK(clk), .RN(n1177), .Q(
        DP_coeffs_fb_int[35]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_13_ ( .D(n1317), .CK(clk), .RN(n1177), .Q(
        DP_coeffs_fb_int[34]), .QN(n1008) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_14_ ( .D(n1318), .CK(clk), .RN(n1177), .Q(
        DP_coeffs_fb_int[33]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_15_ ( .D(n1319), .CK(clk), .RN(n1177), .Q(
        DP_coeffs_fb_int[32]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_16_ ( .D(n1320), .CK(clk), .RN(n1177), .Q(
        DP_coeffs_fb_int[31]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_17_ ( .D(n1321), .CK(clk), .RN(n1177), .Q(
        DP_coeffs_fb_int[30]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_18_ ( .D(n1322), .CK(clk), .RN(n1177), .Q(
        DP_coeffs_fb_int[29]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_19_ ( .D(n1323), .CK(clk), .RN(n1177), .Q(
        DP_coeffs_fb_int[28]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_20_ ( .D(n1324), .CK(clk), .RN(n1177), .Q(
        DP_coeffs_fb_int[27]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_21_ ( .D(n1325), .CK(clk), .RN(n1177), .Q(
        DP_coeffs_fb_int[26]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_22_ ( .D(n1326), .CK(clk), .RN(n1177), .Q(
        DP_coeffs_fb_int[25]) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_23_ ( .D(n1327), .CK(clk), .RN(n1177), .Q(
        DP_coeffs_fb_int[24]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_0_ ( .D(n1328), .CK(clk), .RN(n1178), .Q(
        DP_coeffs_ff_int[23]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_1_ ( .D(n1329), .CK(clk), .RN(n1178), .Q(
        DP_coeffs_ff_int[22]), .QN(n1137) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_2_ ( .D(n1330), .CK(clk), .RN(n1178), .Q(
        DP_coeffs_ff_int[21]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_3_ ( .D(n1331), .CK(clk), .RN(n1178), .Q(
        DP_coeffs_ff_int[20]), .QN(n997) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_4_ ( .D(n1332), .CK(clk), .RN(n1178), .Q(
        DP_coeffs_ff_int[19]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_5_ ( .D(n1333), .CK(clk), .RN(n1178), .Q(
        DP_coeffs_ff_int[18]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_6_ ( .D(n1334), .CK(clk), .RN(n1178), .Q(
        DP_coeffs_ff_int[17]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_7_ ( .D(n1335), .CK(clk), .RN(n1178), .Q(
        DP_coeffs_ff_int[16]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_8_ ( .D(n1336), .CK(clk), .RN(n1178), .Q(
        DP_coeffs_ff_int[15]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_9_ ( .D(n1337), .CK(clk), .RN(n1178), .Q(
        DP_coeffs_ff_int[14]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_10_ ( .D(n1338), .CK(clk), .RN(n1178), .Q(
        DP_coeffs_ff_int[13]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_11_ ( .D(n1339), .CK(clk), .RN(n1178), .Q(
        DP_coeffs_ff_int[12]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_12_ ( .D(n1340), .CK(clk), .RN(n1179), .Q(
        DP_coeffs_ff_int[11]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_13_ ( .D(n1341), .CK(clk), .RN(n1179), .Q(
        DP_coeffs_ff_int[10]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_14_ ( .D(n1342), .CK(clk), .RN(n1179), .Q(
        DP_coeffs_ff_int[9]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_15_ ( .D(n1343), .CK(clk), .RN(n1179), .Q(
        DP_coeffs_ff_int[8]), .QN(n1076) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_16_ ( .D(n1344), .CK(clk), .RN(n1179), .Q(
        DP_coeffs_ff_int[7]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_17_ ( .D(n1345), .CK(clk), .RN(n1179), .Q(
        DP_coeffs_ff_int[6]), .QN(n1047) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_18_ ( .D(n1346), .CK(clk), .RN(n1179), .Q(
        DP_coeffs_ff_int[5]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_19_ ( .D(n1347), .CK(clk), .RN(n1179), .Q(
        DP_coeffs_ff_int[4]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_20_ ( .D(n1348), .CK(clk), .RN(n1179), .Q(
        DP_coeffs_ff_int[3]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_21_ ( .D(n1349), .CK(clk), .RN(n1179), .Q(
        DP_coeffs_ff_int[2]), .QN(n1141) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_22_ ( .D(n1350), .CK(clk), .RN(n1179), .Q(
        DP_coeffs_ff_int[1]) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_23_ ( .D(n1351), .CK(clk), .RN(n1179), .Q(
        DP_coeffs_ff_int[0]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_0_ ( .D(n1352), .CK(clk), .RN(n1180), .Q(
        DP_coeffs_ff_int[47]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_1_ ( .D(n1353), .CK(clk), .RN(n1180), .Q(
        DP_coeffs_ff_int[46]), .QN(n1096) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_2_ ( .D(n1354), .CK(clk), .RN(n1180), .Q(
        DP_coeffs_ff_int[45]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_3_ ( .D(n1355), .CK(clk), .RN(n1180), .Q(
        DP_coeffs_ff_int[44]), .QN(n1053) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_4_ ( .D(n1356), .CK(clk), .RN(n1180), .Q(
        DP_coeffs_ff_int[43]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_5_ ( .D(n1357), .CK(clk), .RN(n1180), .Q(
        DP_coeffs_ff_int[42]), .QN(n1057) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_6_ ( .D(n1358), .CK(clk), .RN(n1180), .Q(
        DP_coeffs_ff_int[41]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_7_ ( .D(n1359), .CK(clk), .RN(n1180), .Q(
        DP_coeffs_ff_int[40]), .QN(n1060) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_8_ ( .D(n1360), .CK(clk), .RN(n1180), .Q(
        DP_coeffs_ff_int[39]), .QN(n1017) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_9_ ( .D(n1361), .CK(clk), .RN(n1180), .Q(
        DP_coeffs_ff_int[38]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_10_ ( .D(n1362), .CK(clk), .RN(n1180), .Q(
        DP_coeffs_ff_int[37]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_11_ ( .D(n1363), .CK(clk), .RN(n1180), .Q(
        DP_coeffs_ff_int[36]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_12_ ( .D(n1364), .CK(clk), .RN(n1181), .Q(
        DP_coeffs_ff_int[35]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_13_ ( .D(n1365), .CK(clk), .RN(n1181), .Q(
        DP_coeffs_ff_int[34]), .QN(n1021) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_14_ ( .D(n1366), .CK(clk), .RN(n1181), .Q(
        DP_coeffs_ff_int[33]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_15_ ( .D(n1367), .CK(clk), .RN(n1181), .Q(
        DP_coeffs_ff_int[32]), .QN(n1029) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_16_ ( .D(n1368), .CK(clk), .RN(n1181), .Q(
        DP_coeffs_ff_int[31]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_17_ ( .D(n1369), .CK(clk), .RN(n1181), .Q(
        DP_coeffs_ff_int[30]), .QN(n1025) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_18_ ( .D(n1370), .CK(clk), .RN(n1181), .Q(
        DP_coeffs_ff_int[29]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_19_ ( .D(n1371), .CK(clk), .RN(n1181), .Q(
        DP_coeffs_ff_int[28]), .QN(n1023) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_20_ ( .D(n1372), .CK(clk), .RN(n1181), .Q(
        DP_coeffs_ff_int[27]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_21_ ( .D(n1373), .CK(clk), .RN(n1181), .Q(
        DP_coeffs_ff_int[26]), .QN(n1066) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_22_ ( .D(n1374), .CK(clk), .RN(n1181), .Q(
        DP_coeffs_ff_int[25]) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_23_ ( .D(n1375), .CK(clk), .RN(n1181), .Q(
        DP_coeffs_ff_int[24]), .QN(n1094) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_0_ ( .D(n1376), .CK(clk), .RN(n1182), .Q(
        DP_coeffs_ff_int[71]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_1_ ( .D(n1377), .CK(clk), .RN(n1182), .Q(
        DP_coeffs_ff_int[70]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_2_ ( .D(n1378), .CK(clk), .RN(n1182), .Q(
        DP_coeffs_ff_int[69]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_3_ ( .D(n1379), .CK(clk), .RN(n1182), .Q(
        DP_coeffs_ff_int[68]), .QN(n1070) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_4_ ( .D(n1380), .CK(clk), .RN(n1182), .Q(
        DP_coeffs_ff_int[67]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_5_ ( .D(n1381), .CK(clk), .RN(n1182), .Q(
        DP_coeffs_ff_int[66]), .QN(n1109) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_6_ ( .D(n1382), .CK(clk), .RN(n1182), .Q(
        DP_coeffs_ff_int[65]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_7_ ( .D(n1383), .CK(clk), .RN(n1182), .Q(
        DP_coeffs_ff_int[64]), .QN(n1103) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_8_ ( .D(n1384), .CK(clk), .RN(n1182), .Q(
        DP_coeffs_ff_int[63]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_9_ ( .D(n1385), .CK(clk), .RN(n1182), .Q(
        DP_coeffs_ff_int[62]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_10_ ( .D(n1386), .CK(clk), .RN(n1182), .Q(
        DP_coeffs_ff_int[61]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_11_ ( .D(n1387), .CK(clk), .RN(n1182), .Q(
        DP_coeffs_ff_int[60]), .QN(n1051) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_12_ ( .D(n1388), .CK(clk), .RN(n1183), .Q(
        DP_coeffs_ff_int[59]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_13_ ( .D(n1389), .CK(clk), .RN(n1183), .Q(
        DP_coeffs_ff_int[58]), .QN(n1044) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_14_ ( .D(n1390), .CK(clk), .RN(n1183), .Q(
        DP_coeffs_ff_int[57]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_15_ ( .D(n1391), .CK(clk), .RN(n1183), .Q(
        DP_coeffs_ff_int[56]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_16_ ( .D(n1392), .CK(clk), .RN(n1183), .Q(
        DP_coeffs_ff_int[55]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_17_ ( .D(n1393), .CK(clk), .RN(n1183), .Q(
        DP_coeffs_ff_int[54]), .QN(n1006) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_18_ ( .D(n1394), .CK(clk), .RN(n1183), .Q(
        DP_coeffs_ff_int[53]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_19_ ( .D(n1395), .CK(clk), .RN(n1183), .Q(
        DP_coeffs_ff_int[52]), .QN(n1040) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_20_ ( .D(n1396), .CK(clk), .RN(n1183), .Q(
        DP_coeffs_ff_int[51]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_21_ ( .D(n1397), .CK(clk), .RN(n1183), .Q(
        DP_coeffs_ff_int[50]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_22_ ( .D(n1398), .CK(clk), .RN(n1183), .Q(
        DP_coeffs_ff_int[49]) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_23_ ( .D(n1399), .CK(clk), .RN(n1183), .Q(
        DP_coeffs_ff_int[48]), .QN(n1000) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_0_ ( .D(n1400), .CK(clk), .RN(n1184), .Q(
        DP_coeffs_ff_int[95]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_1_ ( .D(n1401), .CK(clk), .RN(n1184), .Q(
        DP_coeffs_ff_int[94]), .QN(n1101) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_2_ ( .D(n1402), .CK(clk), .RN(n1184), .Q(
        DP_coeffs_ff_int[93]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_3_ ( .D(n1403), .CK(clk), .RN(n1184), .Q(
        DP_coeffs_ff_int[92]), .QN(n1091) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_4_ ( .D(n1404), .CK(clk), .RN(n1184), .Q(
        DP_coeffs_ff_int[91]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_5_ ( .D(n1405), .CK(clk), .RN(n1184), .Q(
        DP_coeffs_ff_int[90]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_6_ ( .D(n1406), .CK(clk), .RN(n1184), .Q(
        DP_coeffs_ff_int[89]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_7_ ( .D(n1407), .CK(clk), .RN(n1184), .Q(
        DP_coeffs_ff_int[88]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_8_ ( .D(n1408), .CK(clk), .RN(n1184), .Q(
        DP_coeffs_ff_int[87]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_9_ ( .D(n1409), .CK(clk), .RN(n1184), .Q(
        DP_coeffs_ff_int[86]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_10_ ( .D(n1410), .CK(clk), .RN(n1184), .Q(
        DP_coeffs_ff_int[85]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_11_ ( .D(n1411), .CK(clk), .RN(n1184), .Q(
        DP_coeffs_ff_int[84]), .QN(n1019) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_12_ ( .D(n1412), .CK(clk), .RN(n1185), .Q(
        DP_coeffs_ff_int[83]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_13_ ( .D(n1413), .CK(clk), .RN(n1185), .Q(
        DP_coeffs_ff_int[82]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_14_ ( .D(n1414), .CK(clk), .RN(n1185), .Q(
        DP_coeffs_ff_int[81]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_15_ ( .D(n1415), .CK(clk), .RN(n1185), .Q(
        DP_coeffs_ff_int[80]), .QN(n1080) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_16_ ( .D(n1416), .CK(clk), .RN(n1185), .Q(
        DP_coeffs_ff_int[79]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_17_ ( .D(n1417), .CK(clk), .RN(n1185), .Q(
        DP_coeffs_ff_int[78]), .QN(n1072) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_18_ ( .D(n1418), .CK(clk), .RN(n1185), .Q(
        DP_coeffs_ff_int[77]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_19_ ( .D(n1419), .CK(clk), .RN(n1185), .Q(
        DP_coeffs_ff_int[76]), .QN(n1074) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_20_ ( .D(n1420), .CK(clk), .RN(n1185), .Q(
        DP_coeffs_ff_int[75]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_21_ ( .D(n1421), .CK(clk), .RN(n1185), .Q(
        DP_coeffs_ff_int[74]), .QN(n1027) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_22_ ( .D(n1422), .CK(clk), .RN(n1185), .Q(
        DP_coeffs_ff_int[73]) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_23_ ( .D(n1423), .CK(clk), .RN(n1185), .Q(
        DP_coeffs_ff_int[72]) );
  DFFR_X1 DP_reg_ret0_Q_reg_0_ ( .D(DP_sw0_coeff_ret0[0]), .CK(clk), .RN(n1186), .Q(DP_ret0[0]) );
  DFFR_X1 DP_reg_ret0_Q_reg_1_ ( .D(DP_sw0_coeff_ret0[1]), .CK(clk), .RN(n1186), .Q(DP_ret0[1]) );
  DFFR_X1 DP_reg_ret0_Q_reg_2_ ( .D(DP_sw0_coeff_ret0[2]), .CK(clk), .RN(n1186), .Q(DP_ret0[2]) );
  DFFR_X1 DP_reg_ret0_Q_reg_3_ ( .D(DP_sw0_coeff_ret0[3]), .CK(clk), .RN(n1186), .Q(DP_ret0[3]) );
  DFFR_X1 DP_reg_ret0_Q_reg_4_ ( .D(DP_sw0_coeff_ret0[4]), .CK(clk), .RN(n1186), .Q(DP_ret0[4]) );
  DFFR_X1 DP_reg_ret0_Q_reg_5_ ( .D(DP_sw0_coeff_ret0[5]), .CK(clk), .RN(n1186), .Q(DP_ret0[5]) );
  DFFR_X1 DP_reg_ret0_Q_reg_6_ ( .D(DP_sw0_coeff_ret0[6]), .CK(clk), .RN(n1186), .Q(DP_ret0[6]) );
  DFFR_X1 DP_reg_ret0_Q_reg_7_ ( .D(DP_sw0_coeff_ret0[7]), .CK(clk), .RN(n1186), .Q(DP_ret0[7]) );
  DFFR_X1 DP_reg_ret0_Q_reg_8_ ( .D(DP_sw0_coeff_ret0[8]), .CK(clk), .RN(n1186), .Q(DP_ret0[8]) );
  DFFR_X1 DP_reg_ret0_Q_reg_9_ ( .D(DP_sw0_coeff_ret0[9]), .CK(clk), .RN(n1186), .Q(DP_ret0[9]) );
  DFFR_X1 DP_reg_ret0_Q_reg_10_ ( .D(DP_sw0_coeff_ret0[10]), .CK(clk), .RN(
        n1186), .Q(DP_ret0[10]) );
  DFFR_X1 DP_reg_ret0_Q_reg_11_ ( .D(DP_sw0_coeff_ret0[11]), .CK(clk), .RN(
        n1186), .Q(DP_ret0[11]) );
  DFFR_X1 DP_reg_ret0_Q_reg_12_ ( .D(DP_sw0_coeff_ret0[12]), .CK(clk), .RN(
        n1187), .Q(DP_ret0[12]) );
  DFFR_X1 DP_reg_ret0_Q_reg_13_ ( .D(DP_sw0_coeff_ret0[13]), .CK(clk), .RN(
        n1187), .Q(DP_ret0[13]) );
  DFFR_X1 DP_reg_ret0_Q_reg_14_ ( .D(DP_sw0_coeff_ret0[14]), .CK(clk), .RN(
        n1187), .Q(DP_ret0[14]) );
  DFFR_X1 DP_reg_ret0_Q_reg_15_ ( .D(DP_sw0_coeff_ret0[15]), .CK(clk), .RN(
        n1187), .Q(DP_ret0[15]) );
  DFFR_X1 DP_reg_ret0_Q_reg_16_ ( .D(DP_sw0_coeff_ret0[16]), .CK(clk), .RN(
        n1187), .Q(DP_ret0[16]) );
  DFFR_X1 DP_reg_ret0_Q_reg_17_ ( .D(DP_sw0_coeff_ret0[17]), .CK(clk), .RN(
        n1187), .Q(DP_ret0[17]) );
  DFFR_X1 DP_reg_ret0_Q_reg_18_ ( .D(DP_sw0_coeff_ret0[18]), .CK(clk), .RN(
        n1187), .Q(DP_ret0[18]) );
  DFFR_X1 DP_reg_ret0_Q_reg_19_ ( .D(DP_sw0_coeff_ret0[19]), .CK(clk), .RN(
        n1187), .Q(DP_ret0[19]) );
  DFFR_X1 DP_reg_ret0_Q_reg_20_ ( .D(DP_sw0_coeff_ret0[20]), .CK(clk), .RN(
        n1187), .Q(DP_ret0[20]) );
  DFFR_X1 DP_reg_ret0_Q_reg_21_ ( .D(DP_sw0_coeff_ret0[21]), .CK(clk), .RN(
        n1187), .Q(DP_ret0[21]) );
  DFFR_X1 DP_reg_ret0_Q_reg_22_ ( .D(DP_sw0_coeff_ret0[22]), .CK(clk), .RN(
        n1187), .Q(DP_ret0[22]) );
  DFFR_X1 DP_reg_ret0_Q_reg_23_ ( .D(DP_sw0_coeff_ret0[23]), .CK(clk), .RN(
        n1187), .Q(DP_ret0[23]) );
  DFFR_X1 DP_reg_ret1_Q_reg_0_ ( .D(DP_sw1_coeff_ret1[0]), .CK(clk), .RN(n1188), .Q(DP_ret1[0]) );
  DFFR_X1 DP_reg_ret1_Q_reg_1_ ( .D(DP_sw1_coeff_ret1[1]), .CK(clk), .RN(n1188), .Q(DP_ret1[1]) );
  DFFR_X1 DP_reg_ret1_Q_reg_2_ ( .D(DP_sw1_coeff_ret1[2]), .CK(clk), .RN(n1188), .Q(DP_ret1[2]) );
  DFFR_X1 DP_reg_ret1_Q_reg_3_ ( .D(DP_sw1_coeff_ret1[3]), .CK(clk), .RN(n1188), .Q(DP_ret1[3]) );
  DFFR_X1 DP_reg_ret1_Q_reg_4_ ( .D(DP_sw1_coeff_ret1[4]), .CK(clk), .RN(n1188), .Q(DP_ret1[4]) );
  DFFR_X1 DP_reg_ret1_Q_reg_5_ ( .D(DP_sw1_coeff_ret1[5]), .CK(clk), .RN(n1188), .Q(DP_ret1[5]) );
  DFFR_X1 DP_reg_ret1_Q_reg_6_ ( .D(DP_sw1_coeff_ret1[6]), .CK(clk), .RN(n1188), .Q(DP_ret1[6]) );
  DFFR_X1 DP_reg_ret1_Q_reg_7_ ( .D(DP_sw1_coeff_ret1[7]), .CK(clk), .RN(n1188), .Q(DP_ret1[7]) );
  DFFR_X1 DP_reg_ret1_Q_reg_8_ ( .D(DP_sw1_coeff_ret1[8]), .CK(clk), .RN(n1188), .Q(DP_ret1[8]) );
  DFFR_X1 DP_reg_ret1_Q_reg_10_ ( .D(DP_sw1_coeff_ret1[10]), .CK(clk), .RN(
        n1188), .Q(DP_ret1[10]) );
  DFFR_X1 DP_reg_ret1_Q_reg_11_ ( .D(DP_sw1_coeff_ret1[11]), .CK(clk), .RN(
        n1188), .Q(DP_ret1[11]) );
  DFFR_X1 DP_reg_ret1_Q_reg_12_ ( .D(DP_sw1_coeff_ret1[12]), .CK(clk), .RN(
        n1189), .Q(DP_ret1[12]) );
  DFFR_X1 DP_reg_ret1_Q_reg_14_ ( .D(DP_sw1_coeff_ret1[14]), .CK(clk), .RN(
        n1189), .Q(DP_ret1[14]) );
  DFFR_X1 DP_reg_ret1_Q_reg_17_ ( .D(DP_sw1_coeff_ret1[17]), .CK(clk), .RN(
        n1189), .Q(DP_ret1[17]) );
  DFFR_X1 DP_reg_ret1_Q_reg_21_ ( .D(DP_sw1_coeff_ret1[21]), .CK(clk), .RN(
        n1189), .Q(DP_ret1[21]) );
  DFFR_X1 DP_reg_ret1_Q_reg_23_ ( .D(DP_sw1_coeff_ret1[23]), .CK(clk), .RN(
        n1189), .Q(DP_ret1[23]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_0_ ( .D(DP_w_0_), .CK(clk), .RN(n1190), .Q(
        DP_pipe00[0]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_1_ ( .D(DP_w_1_), .CK(clk), .RN(n1190), .Q(
        DP_pipe00[1]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_2_ ( .D(DP_w_2_), .CK(clk), .RN(n1190), .Q(
        DP_pipe00[2]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_3_ ( .D(DP_w_3_), .CK(clk), .RN(n1190), .Q(
        DP_pipe00[3]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_4_ ( .D(DP_w_4_), .CK(clk), .RN(n1190), .Q(
        DP_pipe00[4]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_5_ ( .D(DP_w_5_), .CK(clk), .RN(n1190), .Q(
        DP_pipe00[5]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_6_ ( .D(DP_w_6_), .CK(clk), .RN(n1190), .Q(
        DP_pipe00[6]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_7_ ( .D(DP_w_7_), .CK(clk), .RN(n1190), .Q(
        DP_pipe00[7]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_8_ ( .D(DP_w_8_), .CK(clk), .RN(n1190), .Q(
        DP_pipe00[8]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_9_ ( .D(DP_w_9_), .CK(clk), .RN(n1190), .Q(
        DP_pipe00[9]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_10_ ( .D(DP_w_10_), .CK(clk), .RN(n1190), .Q(
        DP_pipe00[10]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_11_ ( .D(DP_w_11_), .CK(clk), .RN(n1190), .Q(
        DP_pipe00[11]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_12_ ( .D(DP_w_12_), .CK(clk), .RN(n1191), .Q(
        DP_pipe00[12]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_13_ ( .D(DP_w_13_), .CK(clk), .RN(n1191), .Q(
        DP_pipe00[13]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_14_ ( .D(DP_w_14_), .CK(clk), .RN(n1191), .Q(
        DP_pipe00[14]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_15_ ( .D(DP_w_15_), .CK(clk), .RN(n1191), .Q(
        DP_pipe00[15]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_16_ ( .D(DP_w_16_), .CK(clk), .RN(n1191), .Q(
        DP_pipe00[16]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_17_ ( .D(DP_w_17_), .CK(clk), .RN(n1191), .Q(
        DP_pipe00[17]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_18_ ( .D(DP_w_18_), .CK(clk), .RN(n1191), .Q(
        DP_pipe00[18]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_19_ ( .D(DP_w_19_), .CK(clk), .RN(n1191), .Q(
        DP_pipe00[19]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_20_ ( .D(DP_w_20_), .CK(clk), .RN(n1191), .Q(
        DP_pipe00[20]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_21_ ( .D(DP_w_21_), .CK(clk), .RN(n1191), .Q(
        DP_pipe00[21]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_22_ ( .D(DP_w_22_), .CK(clk), .RN(n1191), .Q(
        DP_pipe00[22]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_23_ ( .D(DP_w_23_), .CK(clk), .RN(n1191), .Q(
        DP_pipe00[23]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_0_ ( .D(DP_pipe0_coeff_pipe00[0]), .CK(clk), 
        .RN(n1192), .Q(DP_pipe10[0]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_1_ ( .D(DP_pipe0_coeff_pipe00[1]), .CK(clk), 
        .RN(n1192), .Q(DP_pipe10[1]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_2_ ( .D(DP_pipe0_coeff_pipe00[2]), .CK(clk), 
        .RN(n1192), .Q(DP_pipe10[2]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_3_ ( .D(DP_pipe0_coeff_pipe00[3]), .CK(clk), 
        .RN(n1192), .Q(DP_pipe10[3]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_4_ ( .D(DP_pipe0_coeff_pipe00[4]), .CK(clk), 
        .RN(n1192), .Q(DP_pipe10[4]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_5_ ( .D(DP_pipe0_coeff_pipe00[5]), .CK(clk), 
        .RN(n1192), .Q(DP_pipe10[5]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_6_ ( .D(DP_pipe0_coeff_pipe00[6]), .CK(clk), 
        .RN(n1192), .Q(DP_pipe10[6]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_7_ ( .D(DP_pipe0_coeff_pipe00[7]), .CK(clk), 
        .RN(n1192), .Q(DP_pipe10[7]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_8_ ( .D(DP_pipe0_coeff_pipe00[8]), .CK(clk), 
        .RN(n1192), .Q(DP_pipe10[8]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_9_ ( .D(DP_pipe0_coeff_pipe00[9]), .CK(clk), 
        .RN(n1192), .Q(DP_pipe10[9]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_10_ ( .D(DP_pipe0_coeff_pipe00[10]), .CK(clk), 
        .RN(n1192), .Q(DP_pipe10[10]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_11_ ( .D(DP_pipe0_coeff_pipe00[11]), .CK(clk), 
        .RN(n1192), .Q(DP_pipe10[11]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_12_ ( .D(DP_pipe0_coeff_pipe00[12]), .CK(clk), 
        .RN(n1193), .Q(DP_pipe10[12]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_23_ ( .D(DP_pipe0_coeff_pipe00[23]), .CK(clk), 
        .RN(n1193), .Q(DP_pipe10[23]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_0_ ( .D(DP_pipe0_coeff_pipe01[0]), .CK(clk), 
        .RN(n1194), .Q(DP_pipe11[0]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_1_ ( .D(DP_pipe0_coeff_pipe01[1]), .CK(clk), 
        .RN(n1194), .Q(DP_pipe11[1]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_2_ ( .D(DP_pipe0_coeff_pipe01[2]), .CK(clk), 
        .RN(n1194), .Q(DP_pipe11[2]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_3_ ( .D(DP_pipe0_coeff_pipe01[3]), .CK(clk), 
        .RN(n1194), .Q(DP_pipe11[3]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_4_ ( .D(DP_pipe0_coeff_pipe01[4]), .CK(clk), 
        .RN(n1194), .Q(DP_pipe11[4]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_5_ ( .D(DP_pipe0_coeff_pipe01[5]), .CK(clk), 
        .RN(n1194), .Q(DP_pipe11[5]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_6_ ( .D(DP_pipe0_coeff_pipe01[6]), .CK(clk), 
        .RN(n1194), .Q(DP_pipe11[6]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_7_ ( .D(DP_pipe0_coeff_pipe01[7]), .CK(clk), 
        .RN(n1194), .Q(DP_pipe11[7]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_8_ ( .D(DP_pipe0_coeff_pipe01[8]), .CK(clk), 
        .RN(n1194), .Q(DP_pipe11[8]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_9_ ( .D(DP_pipe0_coeff_pipe01[9]), .CK(clk), 
        .RN(n1194), .Q(DP_pipe11[9]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_10_ ( .D(DP_pipe0_coeff_pipe01[10]), .CK(clk), 
        .RN(n1194), .Q(DP_pipe11[10]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_11_ ( .D(DP_pipe0_coeff_pipe01[11]), .CK(clk), 
        .RN(n1194), .Q(DP_pipe11[11]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_23_ ( .D(DP_pipe0_coeff_pipe01[23]), .CK(clk), 
        .RN(n1195), .Q(DP_pipe11[23]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_0_ ( .D(DP_pipe0_coeff_pipe02[0]), .CK(clk), 
        .RN(n1196), .Q(DP_pipe12[0]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_1_ ( .D(DP_pipe0_coeff_pipe02[1]), .CK(clk), 
        .RN(n1196), .Q(DP_pipe12[1]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_2_ ( .D(DP_pipe0_coeff_pipe02[2]), .CK(clk), 
        .RN(n1196), .Q(DP_pipe12[2]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_3_ ( .D(DP_pipe0_coeff_pipe02[3]), .CK(clk), 
        .RN(n1196), .Q(DP_pipe12[3]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_4_ ( .D(DP_pipe0_coeff_pipe02[4]), .CK(clk), 
        .RN(n1196), .Q(DP_pipe12[4]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_5_ ( .D(DP_pipe0_coeff_pipe02[5]), .CK(clk), 
        .RN(n1196), .Q(DP_pipe12[5]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_6_ ( .D(DP_pipe0_coeff_pipe02[6]), .CK(clk), 
        .RN(n1196), .Q(DP_pipe12[6]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_7_ ( .D(DP_pipe0_coeff_pipe02[7]), .CK(clk), 
        .RN(n1196), .Q(DP_pipe12[7]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_8_ ( .D(DP_pipe0_coeff_pipe02[8]), .CK(clk), 
        .RN(n1196), .Q(DP_pipe12[8]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_9_ ( .D(DP_pipe0_coeff_pipe02[9]), .CK(clk), 
        .RN(n1196), .Q(DP_pipe12[9]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_10_ ( .D(DP_pipe0_coeff_pipe02[10]), .CK(clk), 
        .RN(n1196), .Q(DP_pipe12[10]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_11_ ( .D(DP_pipe0_coeff_pipe02[11]), .CK(clk), 
        .RN(n1196), .Q(DP_pipe12[11]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_12_ ( .D(DP_pipe0_coeff_pipe02[12]), .CK(clk), 
        .RN(n1197), .Q(DP_pipe12[12]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_13_ ( .D(DP_pipe0_coeff_pipe02[13]), .CK(clk), 
        .RN(n1197), .Q(DP_pipe12[13]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_14_ ( .D(DP_pipe0_coeff_pipe02[14]), .CK(clk), 
        .RN(n1197), .Q(DP_pipe12[14]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_15_ ( .D(DP_pipe0_coeff_pipe02[15]), .CK(clk), 
        .RN(n1197), .Q(DP_pipe12[15]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_16_ ( .D(DP_pipe0_coeff_pipe02[16]), .CK(clk), 
        .RN(n1197), .Q(DP_pipe12[16]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_17_ ( .D(DP_pipe0_coeff_pipe02[17]), .CK(clk), 
        .RN(n1197), .Q(DP_pipe12[17]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_18_ ( .D(DP_pipe0_coeff_pipe02[18]), .CK(clk), 
        .RN(n1197), .Q(DP_pipe12[18]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_19_ ( .D(DP_pipe0_coeff_pipe02[19]), .CK(clk), 
        .RN(n1197), .Q(DP_pipe12[19]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_21_ ( .D(DP_pipe0_coeff_pipe02[21]), .CK(clk), 
        .RN(n1197), .Q(DP_pipe12[21]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_22_ ( .D(DP_pipe0_coeff_pipe02[22]), .CK(clk), 
        .RN(n1197), .Q(DP_pipe12[22]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_23_ ( .D(DP_pipe0_coeff_pipe02[23]), .CK(clk), 
        .RN(n1197), .Q(DP_pipe12[23]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_0_ ( .D(DP_pipe0_coeff_pipe03[0]), .CK(clk), 
        .RN(n1198), .Q(DP_pipe13[0]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_1_ ( .D(DP_pipe0_coeff_pipe03[1]), .CK(clk), 
        .RN(n1198), .Q(DP_pipe13[1]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_2_ ( .D(DP_pipe0_coeff_pipe03[2]), .CK(clk), 
        .RN(n1198), .Q(DP_pipe13[2]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_3_ ( .D(DP_pipe0_coeff_pipe03[3]), .CK(clk), 
        .RN(n1198), .Q(DP_pipe13[3]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_4_ ( .D(DP_pipe0_coeff_pipe03[4]), .CK(clk), 
        .RN(n1198), .Q(DP_pipe13[4]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_5_ ( .D(DP_pipe0_coeff_pipe03[5]), .CK(clk), 
        .RN(n1198), .Q(DP_pipe13[5]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_6_ ( .D(DP_pipe0_coeff_pipe03[6]), .CK(clk), 
        .RN(n1198), .Q(DP_pipe13[6]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_7_ ( .D(DP_pipe0_coeff_pipe03[7]), .CK(clk), 
        .RN(n1198), .Q(DP_pipe13[7]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_8_ ( .D(DP_pipe0_coeff_pipe03[8]), .CK(clk), 
        .RN(n1198), .Q(DP_pipe13[8]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_9_ ( .D(DP_pipe0_coeff_pipe03[9]), .CK(clk), 
        .RN(n1198), .Q(DP_pipe13[9]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_10_ ( .D(DP_pipe0_coeff_pipe03[10]), .CK(clk), 
        .RN(n1198), .Q(DP_pipe13[10]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_11_ ( .D(DP_pipe0_coeff_pipe03[11]), .CK(clk), 
        .RN(n1198), .Q(DP_pipe13[11]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_12_ ( .D(DP_pipe0_coeff_pipe03[12]), .CK(clk), 
        .RN(n1199), .Q(DP_pipe13[12]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_23_ ( .D(DP_pipe0_coeff_pipe03[23]), .CK(clk), 
        .RN(n1199), .Q(DP_pipe13[23]) );
  DFFR_X1 CU_presentState_reg_1_ ( .D(n1261), .CK(clk), .RN(n1200), .Q(
        delayed_controls_0__1_), .QN(n1124) );
  DFFR_X1 DP_reg_sw0_Q_reg_23_ ( .D(n1424), .CK(clk), .RN(n1200), .Q(
        DP_sw0_23_), .QN(n1055) );
  DFFR_X1 DP_reg_pipe01_Q_reg_23_ ( .D(DP_sw0_23_), .CK(clk), .RN(n1200), .Q(
        DP_pipe01[23]) );
  DFFR_X1 DP_reg_sw0_Q_reg_22_ ( .D(n1425), .CK(clk), .RN(n1200), .Q(
        DP_sw0_22_), .QN(n1064) );
  DFFR_X1 DP_reg_pipe01_Q_reg_22_ ( .D(DP_sw0_22_), .CK(clk), .RN(n1200), .Q(
        DP_pipe01[22]) );
  DFFR_X1 DP_reg_sw0_Q_reg_21_ ( .D(n1426), .CK(clk), .RN(n1200), .Q(
        DP_sw0_21_) );
  DFFR_X1 DP_reg_pipe01_Q_reg_21_ ( .D(DP_sw0_21_), .CK(clk), .RN(n1200), .Q(
        DP_pipe01[21]) );
  DFFR_X1 DP_reg_sw0_Q_reg_20_ ( .D(n1427), .CK(clk), .RN(n1200), .Q(
        DP_sw0_20_) );
  DFFR_X1 DP_reg_pipe01_Q_reg_20_ ( .D(DP_sw0_20_), .CK(clk), .RN(n1200), .Q(
        DP_pipe01[20]) );
  DFFR_X1 DP_reg_sw0_Q_reg_19_ ( .D(n1428), .CK(clk), .RN(n1200), .Q(
        DP_sw0_19_) );
  DFFR_X1 DP_reg_pipe01_Q_reg_19_ ( .D(DP_sw0_19_), .CK(clk), .RN(n1200), .Q(
        DP_pipe01[19]) );
  DFFR_X1 DP_reg_sw0_Q_reg_18_ ( .D(n1429), .CK(clk), .RN(n1200), .Q(
        DP_sw0_18_) );
  DFFR_X1 DP_reg_pipe01_Q_reg_18_ ( .D(DP_sw0_18_), .CK(clk), .RN(n1201), .Q(
        DP_pipe01[18]) );
  DFFR_X1 DP_reg_sw0_Q_reg_17_ ( .D(n1430), .CK(clk), .RN(n1201), .Q(
        DP_sw0_17_) );
  DFFR_X1 DP_reg_pipe01_Q_reg_17_ ( .D(DP_sw0_17_), .CK(clk), .RN(n1201), .Q(
        DP_pipe01[17]) );
  DFFR_X1 DP_reg_sw0_Q_reg_16_ ( .D(n1431), .CK(clk), .RN(n1201), .Q(
        DP_sw0_16_) );
  DFFR_X1 DP_reg_pipe01_Q_reg_16_ ( .D(DP_sw0_16_), .CK(clk), .RN(n1201), .Q(
        DP_pipe01[16]) );
  DFFR_X1 DP_reg_sw0_Q_reg_15_ ( .D(n1432), .CK(clk), .RN(n1201), .Q(
        DP_sw0_15_) );
  DFFR_X1 DP_reg_pipe01_Q_reg_15_ ( .D(DP_sw0_15_), .CK(clk), .RN(n1201), .Q(
        DP_pipe01[15]) );
  DFFR_X1 DP_reg_sw0_Q_reg_14_ ( .D(n1433), .CK(clk), .RN(n1201), .Q(
        DP_sw0_14_) );
  DFFR_X1 DP_reg_sw0_Q_reg_13_ ( .D(n1434), .CK(clk), .RN(n1201), .Q(
        DP_sw0_13_) );
  DFFR_X1 DP_reg_pipe01_Q_reg_13_ ( .D(DP_sw0_13_), .CK(clk), .RN(n1201), .Q(
        DP_pipe01[13]) );
  DFFR_X1 DP_reg_sw0_Q_reg_12_ ( .D(n1435), .CK(clk), .RN(n1201), .Q(
        DP_sw0_12_) );
  DFFR_X1 DP_reg_pipe01_Q_reg_12_ ( .D(DP_sw0_12_), .CK(clk), .RN(n1202), .Q(
        DP_pipe01[12]) );
  DFFR_X1 DP_reg_sw0_Q_reg_11_ ( .D(n1436), .CK(clk), .RN(n1202), .Q(
        DP_sw0_11_) );
  DFFR_X1 DP_reg_pipe01_Q_reg_11_ ( .D(DP_sw0_11_), .CK(clk), .RN(n1202), .Q(
        DP_pipe01[11]) );
  DFFR_X1 DP_reg_sw0_Q_reg_10_ ( .D(n1437), .CK(clk), .RN(n1202), .Q(
        DP_sw0_10_) );
  DFFR_X1 DP_reg_pipe01_Q_reg_10_ ( .D(DP_sw0_10_), .CK(clk), .RN(n1202), .Q(
        DP_pipe01[10]) );
  DFFR_X1 DP_reg_sw0_Q_reg_9_ ( .D(n1438), .CK(clk), .RN(n1202), .Q(DP_sw0_9_)
         );
  DFFR_X1 DP_reg_pipe01_Q_reg_9_ ( .D(DP_sw0_9_), .CK(clk), .RN(n1202), .Q(
        DP_pipe01[9]) );
  DFFR_X1 DP_reg_sw0_Q_reg_8_ ( .D(n1439), .CK(clk), .RN(n1202), .Q(DP_sw0_8_)
         );
  DFFR_X1 DP_reg_pipe01_Q_reg_8_ ( .D(DP_sw0_8_), .CK(clk), .RN(n1202), .Q(
        DP_pipe01[8]) );
  DFFR_X1 DP_reg_sw0_Q_reg_7_ ( .D(n1440), .CK(clk), .RN(n1202), .Q(DP_sw0_7_)
         );
  DFFR_X1 DP_reg_pipe01_Q_reg_7_ ( .D(DP_sw0_7_), .CK(clk), .RN(n1202), .Q(
        DP_pipe01[7]) );
  DFFR_X1 DP_reg_sw0_Q_reg_6_ ( .D(n1441), .CK(clk), .RN(n1202), .Q(DP_sw0_6_)
         );
  DFFR_X1 DP_reg_pipe01_Q_reg_6_ ( .D(DP_sw0_6_), .CK(clk), .RN(n1203), .Q(
        DP_pipe01[6]) );
  DFFR_X1 DP_reg_sw0_Q_reg_5_ ( .D(n1442), .CK(clk), .RN(n1203), .Q(DP_sw0_5_)
         );
  DFFR_X1 DP_reg_pipe01_Q_reg_5_ ( .D(DP_sw0_5_), .CK(clk), .RN(n1203), .Q(
        DP_pipe01[5]) );
  DFFR_X1 DP_reg_sw0_Q_reg_4_ ( .D(n1443), .CK(clk), .RN(n1203), .Q(DP_sw0_4_)
         );
  DFFR_X1 DP_reg_pipe01_Q_reg_4_ ( .D(DP_sw0_4_), .CK(clk), .RN(n1203), .Q(
        DP_pipe01[4]) );
  DFFR_X1 DP_reg_sw0_Q_reg_3_ ( .D(n1444), .CK(clk), .RN(n1203), .Q(DP_sw0_3_)
         );
  DFFR_X1 DP_reg_pipe01_Q_reg_3_ ( .D(DP_sw0_3_), .CK(clk), .RN(n1203), .Q(
        DP_pipe01[3]) );
  DFFR_X1 DP_reg_sw0_Q_reg_2_ ( .D(n1445), .CK(clk), .RN(n1203), .Q(DP_sw0_2_)
         );
  DFFR_X1 DP_reg_pipe01_Q_reg_2_ ( .D(DP_sw0_2_), .CK(clk), .RN(n1203), .Q(
        DP_pipe01[2]) );
  DFFR_X1 DP_reg_sw0_Q_reg_1_ ( .D(n1446), .CK(clk), .RN(n1203), .Q(DP_sw0_1_)
         );
  DFFR_X1 DP_reg_pipe01_Q_reg_1_ ( .D(DP_sw0_1_), .CK(clk), .RN(n1203), .Q(
        DP_pipe01[1]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_0_ ( .D(DP_sw0_0_), .CK(clk), .RN(n1204), .Q(
        DP_pipe01[0]) );
  DFFR_X1 DP_reg_sw1_Q_reg_23_ ( .D(n1448), .CK(clk), .RN(n1204), .Q(
        DP_sw1_23_) );
  DFFR_X1 DP_reg_pipe02_Q_reg_23_ ( .D(DP_sw1_23_), .CK(clk), .RN(n1204), .Q(
        DP_pipe02[23]) );
  DFFR_X1 DP_reg_sw1_Q_reg_22_ ( .D(n1449), .CK(clk), .RN(n1204), .Q(
        DP_sw1_22_) );
  DFFR_X1 DP_reg_pipe02_Q_reg_22_ ( .D(DP_sw1_22_), .CK(clk), .RN(n1204), .Q(
        DP_pipe02[22]) );
  DFFR_X1 DP_reg_sw1_Q_reg_21_ ( .D(n1450), .CK(clk), .RN(n1204), .Q(
        DP_sw1_21_) );
  DFFR_X1 DP_reg_pipe02_Q_reg_21_ ( .D(DP_sw1_21_), .CK(clk), .RN(n1204), .Q(
        DP_pipe02[21]) );
  DFFR_X1 DP_reg_sw1_Q_reg_20_ ( .D(n1451), .CK(clk), .RN(n1204), .Q(
        DP_sw1_20_) );
  DFFR_X1 DP_reg_pipe02_Q_reg_20_ ( .D(DP_sw1_20_), .CK(clk), .RN(n1204), .Q(
        DP_pipe02[20]) );
  DFFR_X1 DP_reg_sw1_Q_reg_19_ ( .D(n1452), .CK(clk), .RN(n1204), .Q(
        DP_sw1_19_) );
  DFFR_X1 DP_reg_pipe02_Q_reg_19_ ( .D(DP_sw1_19_), .CK(clk), .RN(n1204), .Q(
        DP_pipe02[19]) );
  DFFR_X1 DP_reg_sw1_Q_reg_18_ ( .D(n1453), .CK(clk), .RN(n1204), .Q(
        DP_sw1_18_) );
  DFFR_X1 DP_reg_pipe02_Q_reg_18_ ( .D(DP_sw1_18_), .CK(clk), .RN(n1205), .Q(
        DP_pipe02[18]) );
  DFFR_X1 DP_reg_sw1_Q_reg_17_ ( .D(n1454), .CK(clk), .RN(n1205), .Q(
        DP_sw1_17_) );
  DFFR_X1 DP_reg_pipe02_Q_reg_17_ ( .D(DP_sw1_17_), .CK(clk), .RN(n1205), .Q(
        DP_pipe02[17]) );
  DFFR_X1 DP_reg_sw1_Q_reg_16_ ( .D(n1455), .CK(clk), .RN(n1205), .Q(
        DP_sw1_16_) );
  DFFR_X1 DP_reg_pipe02_Q_reg_16_ ( .D(DP_sw1_16_), .CK(clk), .RN(n1205), .Q(
        DP_pipe02[16]) );
  DFFR_X1 DP_reg_sw1_Q_reg_15_ ( .D(n1456), .CK(clk), .RN(n1205), .Q(
        DP_sw1_15_) );
  DFFR_X1 DP_reg_pipe02_Q_reg_15_ ( .D(DP_sw1_15_), .CK(clk), .RN(n1205), .Q(
        DP_pipe02[15]) );
  DFFR_X1 DP_reg_sw1_Q_reg_14_ ( .D(n1457), .CK(clk), .RN(n1205), .Q(
        DP_sw1_14_) );
  DFFR_X1 DP_reg_pipe02_Q_reg_14_ ( .D(DP_sw1_14_), .CK(clk), .RN(n1205), .Q(
        DP_pipe02[14]) );
  DFFR_X1 DP_reg_sw1_Q_reg_13_ ( .D(n1458), .CK(clk), .RN(n1205), .Q(
        DP_sw1_13_) );
  DFFR_X1 DP_reg_pipe02_Q_reg_13_ ( .D(DP_sw1_13_), .CK(clk), .RN(n1205), .Q(
        DP_pipe02[13]) );
  DFFR_X1 DP_reg_sw1_Q_reg_12_ ( .D(n1459), .CK(clk), .RN(n1205), .Q(
        DP_sw1_12_) );
  DFFR_X1 DP_reg_pipe02_Q_reg_12_ ( .D(DP_sw1_12_), .CK(clk), .RN(n1206), .Q(
        DP_pipe02[12]) );
  DFFR_X1 DP_reg_sw1_Q_reg_11_ ( .D(n1460), .CK(clk), .RN(n1206), .Q(
        DP_sw1_11_) );
  DFFR_X1 DP_reg_pipe02_Q_reg_11_ ( .D(DP_sw1_11_), .CK(clk), .RN(n1206), .Q(
        DP_pipe02[11]) );
  DFFR_X1 DP_reg_sw1_Q_reg_10_ ( .D(n1461), .CK(clk), .RN(n1206), .Q(
        DP_sw1_10_) );
  DFFR_X1 DP_reg_pipe02_Q_reg_10_ ( .D(DP_sw1_10_), .CK(clk), .RN(n1206), .Q(
        DP_pipe02[10]) );
  DFFR_X1 DP_reg_sw1_Q_reg_9_ ( .D(n1462), .CK(clk), .RN(n1206), .Q(DP_sw1_9_)
         );
  DFFR_X1 DP_reg_pipe02_Q_reg_9_ ( .D(DP_sw1_9_), .CK(clk), .RN(n1206), .Q(
        DP_pipe02[9]) );
  DFFR_X1 DP_reg_pipe02_Q_reg_8_ ( .D(DP_sw1_8_), .CK(clk), .RN(n1206), .Q(
        DP_pipe02[8]) );
  DFFR_X1 DP_reg_sw1_Q_reg_7_ ( .D(n1464), .CK(clk), .RN(n1206), .Q(DP_sw1_7_)
         );
  DFFR_X1 DP_reg_pipe02_Q_reg_7_ ( .D(DP_sw1_7_), .CK(clk), .RN(n1206), .Q(
        DP_pipe02[7]) );
  DFFR_X1 DP_reg_sw1_Q_reg_6_ ( .D(n1465), .CK(clk), .RN(n1206), .Q(DP_sw1_6_)
         );
  DFFR_X1 DP_reg_pipe02_Q_reg_6_ ( .D(DP_sw1_6_), .CK(clk), .RN(n1207), .Q(
        DP_pipe02[6]) );
  DFFR_X1 DP_reg_sw1_Q_reg_5_ ( .D(n1466), .CK(clk), .RN(n1207), .Q(DP_sw1_5_)
         );
  DFFR_X1 DP_reg_pipe02_Q_reg_5_ ( .D(DP_sw1_5_), .CK(clk), .RN(n1207), .Q(
        DP_pipe02[5]) );
  DFFR_X1 DP_reg_sw1_Q_reg_4_ ( .D(n1467), .CK(clk), .RN(n1207), .Q(DP_sw1_4_)
         );
  DFFR_X1 DP_reg_pipe02_Q_reg_4_ ( .D(DP_sw1_4_), .CK(clk), .RN(n1207), .Q(
        DP_pipe02[4]) );
  DFFR_X1 DP_reg_sw1_Q_reg_3_ ( .D(n1468), .CK(clk), .RN(n1207), .Q(DP_sw1_3_)
         );
  DFFR_X1 DP_reg_pipe02_Q_reg_3_ ( .D(DP_sw1_3_), .CK(clk), .RN(n1207), .Q(
        DP_pipe02[3]) );
  DFFR_X1 DP_reg_sw1_Q_reg_2_ ( .D(n1469), .CK(clk), .RN(n1207), .Q(DP_sw1_2_)
         );
  DFFR_X1 DP_reg_pipe02_Q_reg_2_ ( .D(DP_sw1_2_), .CK(clk), .RN(n1207), .Q(
        DP_pipe02[2]) );
  DFFR_X1 DP_reg_sw1_Q_reg_1_ ( .D(n1470), .CK(clk), .RN(n1207), .Q(DP_sw1_1_)
         );
  DFFR_X1 DP_reg_pipe02_Q_reg_1_ ( .D(DP_sw1_1_), .CK(clk), .RN(n1207), .Q(
        DP_pipe02[1]) );
  DFFR_X1 DP_reg_sw1_Q_reg_0_ ( .D(n1471), .CK(clk), .RN(n1207), .Q(DP_sw1_0_), 
        .QN(n1068) );
  DFFR_X1 DP_reg_sw2_Q_reg_23_ ( .D(n575), .CK(clk), .RN(n1208), .Q(n1259) );
  DFFR_X1 DP_reg_pipe03_Q_reg_23_ ( .D(n1259), .CK(clk), .RN(n1208), .Q(
        DP_pipe03[23]) );
  DFFR_X1 DP_reg_sw2_Q_reg_22_ ( .D(n573), .CK(clk), .RN(n1208), .Q(n1258) );
  DFFR_X1 DP_reg_pipe03_Q_reg_22_ ( .D(n1258), .CK(clk), .RN(n1208), .Q(
        DP_pipe03[22]) );
  DFFR_X1 DP_reg_sw2_Q_reg_21_ ( .D(n571), .CK(clk), .RN(n1208), .Q(n1257) );
  DFFR_X1 DP_reg_pipe03_Q_reg_21_ ( .D(n1257), .CK(clk), .RN(n1208), .Q(
        DP_pipe03[21]) );
  DFFR_X1 DP_reg_sw2_Q_reg_20_ ( .D(n569), .CK(clk), .RN(n1208), .Q(n1256) );
  DFFR_X1 DP_reg_pipe03_Q_reg_20_ ( .D(n1256), .CK(clk), .RN(n1208), .Q(
        DP_pipe03[20]) );
  DFFR_X1 DP_reg_sw2_Q_reg_19_ ( .D(n567), .CK(clk), .RN(n1208), .Q(n1255) );
  DFFR_X1 DP_reg_pipe03_Q_reg_19_ ( .D(n1255), .CK(clk), .RN(n1208), .Q(
        DP_pipe03[19]) );
  DFFR_X1 DP_reg_sw2_Q_reg_18_ ( .D(n565), .CK(clk), .RN(n1208), .Q(n1254) );
  DFFR_X1 DP_reg_pipe03_Q_reg_18_ ( .D(n1254), .CK(clk), .RN(n1209), .Q(
        DP_pipe03[18]) );
  DFFR_X1 DP_reg_sw2_Q_reg_17_ ( .D(n563), .CK(clk), .RN(n1209), .Q(n1253) );
  DFFR_X1 DP_reg_pipe03_Q_reg_17_ ( .D(n1253), .CK(clk), .RN(n1209), .Q(
        DP_pipe03[17]) );
  DFFR_X1 DP_reg_sw2_Q_reg_16_ ( .D(n561), .CK(clk), .RN(n1209), .Q(n1252) );
  DFFR_X1 DP_reg_pipe03_Q_reg_16_ ( .D(n1252), .CK(clk), .RN(n1209), .Q(
        DP_pipe03[16]) );
  DFFR_X1 DP_reg_sw2_Q_reg_15_ ( .D(n559), .CK(clk), .RN(n1209), .Q(n1251) );
  DFFR_X1 DP_reg_pipe03_Q_reg_15_ ( .D(n1251), .CK(clk), .RN(n1209), .Q(
        DP_pipe03[15]) );
  DFFR_X1 DP_reg_sw2_Q_reg_14_ ( .D(n557), .CK(clk), .RN(n1209), .Q(n1250) );
  DFFR_X1 DP_reg_pipe03_Q_reg_14_ ( .D(n1250), .CK(clk), .RN(n1209), .Q(
        DP_pipe03[14]) );
  DFFR_X1 DP_reg_sw2_Q_reg_13_ ( .D(n555), .CK(clk), .RN(n1209), .Q(n1249) );
  DFFR_X1 DP_reg_pipe03_Q_reg_13_ ( .D(n1249), .CK(clk), .RN(n1209), .Q(
        DP_pipe03[13]) );
  DFFR_X1 DP_reg_sw2_Q_reg_12_ ( .D(n553), .CK(clk), .RN(n1209), .Q(n1248) );
  DFFR_X1 DP_reg_pipe03_Q_reg_12_ ( .D(n1248), .CK(clk), .RN(n1210), .Q(
        DP_pipe03[12]) );
  DFFR_X1 DP_reg_sw2_Q_reg_11_ ( .D(n551), .CK(clk), .RN(n1210), .Q(n1247) );
  DFFR_X1 DP_reg_pipe03_Q_reg_11_ ( .D(n1247), .CK(clk), .RN(n1210), .Q(
        DP_pipe03[11]) );
  DFFR_X1 DP_reg_sw2_Q_reg_10_ ( .D(n549), .CK(clk), .RN(n1210), .Q(n1246) );
  DFFR_X1 DP_reg_pipe03_Q_reg_10_ ( .D(n1246), .CK(clk), .RN(n1210), .Q(
        DP_pipe03[10]) );
  DFFR_X1 DP_reg_sw2_Q_reg_9_ ( .D(n547), .CK(clk), .RN(n1210), .Q(n1245) );
  DFFR_X1 DP_reg_pipe03_Q_reg_9_ ( .D(n1245), .CK(clk), .RN(n1210), .Q(
        DP_pipe03[9]) );
  DFFR_X1 DP_reg_sw2_Q_reg_8_ ( .D(n545), .CK(clk), .RN(n1210), .Q(n1244) );
  DFFR_X1 DP_reg_pipe03_Q_reg_8_ ( .D(n1244), .CK(clk), .RN(n1210), .Q(
        DP_pipe03[8]) );
  DFFR_X1 DP_reg_sw2_Q_reg_7_ ( .D(n543), .CK(clk), .RN(n1210), .Q(n1243) );
  DFFR_X1 DP_reg_pipe03_Q_reg_7_ ( .D(n1243), .CK(clk), .RN(n1210), .Q(
        DP_pipe03[7]) );
  DFFR_X1 DP_reg_sw2_Q_reg_6_ ( .D(n541), .CK(clk), .RN(n1210), .Q(n1242) );
  DFFR_X1 DP_reg_pipe03_Q_reg_6_ ( .D(n1242), .CK(clk), .RN(n1211), .Q(
        DP_pipe03[6]) );
  DFFR_X1 DP_reg_sw2_Q_reg_5_ ( .D(n539), .CK(clk), .RN(n1211), .Q(n1241) );
  DFFR_X1 DP_reg_pipe03_Q_reg_5_ ( .D(n1241), .CK(clk), .RN(n1211), .Q(
        DP_pipe03[5]) );
  DFFR_X1 DP_reg_sw2_Q_reg_4_ ( .D(n537), .CK(clk), .RN(n1211), .Q(n1240) );
  DFFR_X1 DP_reg_pipe03_Q_reg_4_ ( .D(n1240), .CK(clk), .RN(n1211), .Q(
        DP_pipe03[4]) );
  DFFR_X1 DP_reg_sw2_Q_reg_3_ ( .D(n535), .CK(clk), .RN(n1211), .Q(n1239) );
  DFFR_X1 DP_reg_pipe03_Q_reg_3_ ( .D(n1239), .CK(clk), .RN(n1211), .Q(
        DP_pipe03[3]) );
  DFFR_X1 DP_reg_sw2_Q_reg_2_ ( .D(n533), .CK(clk), .RN(n1211), .Q(n1238) );
  DFFR_X1 DP_reg_pipe03_Q_reg_2_ ( .D(n1238), .CK(clk), .RN(n1211), .Q(
        DP_pipe03[2]) );
  DFFR_X1 DP_reg_sw2_Q_reg_1_ ( .D(n531), .CK(clk), .RN(n1211), .Q(n1237) );
  DFFR_X1 DP_reg_pipe03_Q_reg_1_ ( .D(n1237), .CK(clk), .RN(n1211), .Q(
        DP_pipe03[1]) );
  DFFR_X1 DP_reg_sw2_Q_reg_0_ ( .D(n529), .CK(clk), .RN(n1211), .Q(n1236) );
  DFFR_X1 CU_presentState_reg_0_ ( .D(CU_nextState_0_), .CK(clk), .RN(n1212), 
        .QN(n1112) );
  DFFR_X1 reg_delay_0_Q_reg_0_ ( .D(delayed_controls_0__1_), .CK(clk), .RN(
        n1212), .Q(delayed_controls_1__1_) );
  DFFR_X1 reg_delay_0_Q_reg_1_ ( .D(n1261), .CK(clk), .RN(n1212), .Q(
        delayed_controls_1__0_) );
  DFFR_X1 reg_delay_1_Q_reg_0_ ( .D(delayed_controls_1__1_), .CK(clk), .RN(
        n1212), .Q(vOut) );
  DFFR_X1 reg_delay_1_Q_reg_1_ ( .D(delayed_controls_1__0_), .CK(clk), .RN(
        n1212), .Q(delayed_controls_2__0_), .QN(n1123) );
  DFFR_X1 DP_reg_out_Q_reg_11_ ( .D(n524), .CK(clk), .RN(n1212), .Q(dOut[11])
         );
  DFFR_X1 DP_reg_out_Q_reg_10_ ( .D(n523), .CK(clk), .RN(n1212), .Q(dOut[10]), 
        .QN(n280) );
  DFFR_X1 DP_reg_out_Q_reg_9_ ( .D(n522), .CK(clk), .RN(n1212), .Q(dOut[9]) );
  DFFR_X1 DP_reg_out_Q_reg_8_ ( .D(n521), .CK(clk), .RN(n1212), .Q(dOut[8]) );
  DFFR_X1 DP_reg_out_Q_reg_7_ ( .D(n520), .CK(clk), .RN(n1212), .Q(dOut[7]) );
  DFFR_X1 DP_reg_out_Q_reg_6_ ( .D(n519), .CK(clk), .RN(n1212), .Q(dOut[6]) );
  DFFR_X1 DP_reg_out_Q_reg_5_ ( .D(n518), .CK(clk), .RN(n1213), .Q(dOut[5]) );
  DFFR_X1 DP_reg_out_Q_reg_4_ ( .D(n517), .CK(clk), .RN(n1213), .Q(dOut[4]) );
  DFFR_X1 DP_reg_out_Q_reg_3_ ( .D(n516), .CK(clk), .RN(n1213), .Q(dOut[3]) );
  DFFR_X1 DP_reg_out_Q_reg_2_ ( .D(n515), .CK(clk), .RN(n1213), .Q(dOut[2]) );
  DFFR_X1 DP_reg_out_Q_reg_1_ ( .D(n514), .CK(clk), .RN(n1213), .Q(dOut[1]) );
  DFFR_X1 DP_reg_out_Q_reg_0_ ( .D(n513), .CK(clk), .RN(n1213), .Q(dOut[0]) );
  iir_filter_DW01_add_6 add_2_root_add_0_root_DP_add_223 ( .A({DP_pipe11[23], 
        DP_pipe11[22], DP_pipe11[21], DP_pipe11[20], DP_pipe11[19], 
        DP_pipe11[18], DP_pipe11[17], DP_pipe11[16], DP_pipe11[15], 
        DP_pipe11[14], DP_pipe11[13], DP_pipe11[12], DP_pipe11[11], 
        DP_pipe11[10], DP_pipe11[9], DP_pipe11[8], DP_pipe11[7], DP_pipe11[6], 
        DP_pipe11[5], DP_pipe11[4], DP_pipe11[3], DP_pipe11[2], DP_pipe11[1], 
        DP_pipe11[0]}), .B({DP_pipe13[23], DP_pipe13[22], DP_pipe13[21], 
        DP_pipe13[20], DP_pipe13[19], DP_pipe13[18], DP_pipe13[17], 
        DP_pipe13[16], DP_pipe13[15], DP_pipe13[14], DP_pipe13[13], 
        DP_pipe13[12], DP_pipe13[11], DP_pipe13[10], DP_pipe13[9], 
        DP_pipe13[8], DP_pipe13[7], DP_pipe13[6], DP_pipe13[5], DP_pipe13[4], 
        DP_pipe13[3], DP_pipe13[2], DP_pipe13[1], DP_pipe13[0]}), .SUM({
        DP_ff_23_, DP_ff_22_, DP_ff_21_, DP_ff_20_, DP_ff_19_, DP_ff_18_, 
        DP_ff_17_, DP_ff_16_, DP_ff_15_, DP_ff_14_, DP_ff_13_, DP_ff_12_, 
        DP_ff_11_, DP_ff_10_, DP_ff_9_, DP_ff_8_, DP_ff_7_, DP_ff_6_, DP_ff_5_, 
        DP_ff_4_, DP_ff_3_, DP_ff_2_, DP_ff_1_, DP_ff_0_}), .CI(1'b0) );
  iir_filter_DW01_add_5 add_1_root_add_0_root_DP_add_223 ( .A({DP_pipe10[23], 
        DP_pipe10[22], DP_pipe10[21], DP_pipe10[20], DP_pipe10[19], 
        DP_pipe10[18], DP_pipe10[17], DP_pipe10[16], DP_pipe10[15], 
        DP_pipe10[14], DP_pipe10[13], DP_pipe10[12], DP_pipe10[11], 
        DP_pipe10[10], DP_pipe10[9], DP_pipe10[8], DP_pipe10[7], DP_pipe10[6], 
        DP_pipe10[5], DP_pipe10[4], DP_pipe10[3], DP_pipe10[2], DP_pipe10[1], 
        DP_pipe10[0]}), .B({DP_pipe12[23], DP_pipe12[22], DP_pipe12[21], 
        DP_pipe12[20], DP_pipe12[19], DP_pipe12[18], DP_pipe12[17], 
        DP_pipe12[16], DP_pipe12[15], DP_pipe12[14], DP_pipe12[13], 
        DP_pipe12[12], DP_pipe12[11], DP_pipe12[10], DP_pipe12[9], 
        DP_pipe12[8], DP_pipe12[7], DP_pipe12[6], DP_pipe12[5], DP_pipe12[4], 
        DP_pipe12[3], DP_pipe12[2], DP_pipe12[1], DP_pipe12[0]}), .SUM({
        DP_ff_part_23_, DP_ff_part_22_, DP_ff_part_21_, DP_ff_part_20_, 
        DP_ff_part_19_, DP_ff_part_18_, DP_ff_part_17_, DP_ff_part_16_, 
        DP_ff_part_15_, DP_ff_part_14_, DP_ff_part_13_, DP_ff_part_12_, 
        DP_ff_part_11_, DP_ff_part_10_, DP_ff_part_9_, DP_ff_part_8_, 
        DP_ff_part_7_, DP_ff_part_6_, DP_ff_part_5_, DP_ff_part_4_, 
        DP_ff_part_3_, DP_ff_part_2_, DP_ff_part_1_, DP_ff_part_0_}), .CI(1'b0) );
  iir_filter_DW01_add_1 add_1_root_sub_0_root_DP_sub_217 ( .A({DP_ret0[23], 
        DP_ret0[22], DP_ret0[21], DP_ret0[20], DP_ret0[19], DP_ret0[18], 
        DP_ret0[17], DP_ret0[16], DP_ret0[15], DP_ret0[14], DP_ret0[13], 
        DP_ret0[12], DP_ret0[11], DP_ret0[10], DP_ret0[9], DP_ret0[8], 
        DP_ret0[7], DP_ret0[6], DP_ret0[5], DP_ret0[4], DP_ret0[3], DP_ret0[2], 
        DP_ret0[1], DP_ret0[0]}), .B({DP_ret1[23], DP_ret1[22], DP_ret1[21], 
        DP_ret1[20], DP_ret1[19], DP_ret1[18], DP_ret1[17], DP_ret1[16], 
        DP_ret1[15], DP_ret1[14], DP_ret1[13], DP_ret1[12], DP_ret1[11], 
        DP_ret1[10], DP_ret1[9], DP_ret1[8], DP_ret1[7], DP_ret1[6], 
        DP_ret1[5], DP_ret1[4], DP_ret1[3], DP_ret1[2], DP_ret1[1], DP_ret1[0]}), .SUM({DP_fb_23_, DP_fb_22_, DP_fb_21_, DP_fb_20_, DP_fb_19_, DP_fb_18_, 
        DP_fb_17_, DP_fb_16_, DP_fb_15_, DP_fb_14_, DP_fb_13_, DP_fb_12_, 
        DP_fb_11_, DP_fb_10_, DP_fb_9_, DP_fb_8_, DP_fb_7_, DP_fb_6_, DP_fb_5_, 
        DP_fb_4_, DP_fb_3_, DP_fb_2_, DP_fb_1_, DP_fb_0_}), .CI(1'b0) );
  iir_filter_DW01_sub_1 sub_0_root_sub_0_root_DP_sub_217 ( .A({DP_x[11], 
        DP_x[11], DP_x[10], DP_x[9], DP_x[8], DP_x[7], DP_x[6], DP_x[5], 
        DP_x[4], DP_x[3], DP_x[2], DP_x[1], DP_x[0], 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({DP_fb_23_, DP_fb_22_, 
        DP_fb_21_, DP_fb_20_, DP_fb_19_, DP_fb_18_, DP_fb_17_, DP_fb_16_, 
        DP_fb_15_, DP_fb_14_, DP_fb_13_, DP_fb_12_, DP_fb_11_, DP_fb_10_, 
        DP_fb_9_, DP_fb_8_, DP_fb_7_, DP_fb_6_, DP_fb_5_, DP_fb_4_, DP_fb_3_, 
        DP_fb_2_, DP_fb_1_, DP_fb_0_}), .DIFF({DP_w_23_, DP_w_22_, DP_w_21_, 
        DP_w_20_, DP_w_19_, DP_w_18_, DP_w_17_, DP_w_16_, DP_w_15_, DP_w_14_, 
        DP_w_13_, DP_w_12_, DP_w_11_, DP_w_10_, DP_w_9_, DP_w_8_, DP_w_7_, 
        DP_w_6_, DP_w_5_, DP_w_4_, DP_w_3_, DP_w_2_, DP_w_1_, DP_w_0_}), .CI(
        1'b0) );
  iir_filter_DW01_add_2 add_0_root_add_0_root_DP_add_223 ( .A({DP_ff_23_, 
        DP_ff_22_, DP_ff_21_, DP_ff_20_, DP_ff_19_, DP_ff_18_, DP_ff_17_, 
        DP_ff_16_, DP_ff_15_, DP_ff_14_, DP_ff_13_, DP_ff_12_, DP_ff_11_, 
        DP_ff_10_, DP_ff_9_, DP_ff_8_, DP_ff_7_, DP_ff_6_, DP_ff_5_, DP_ff_4_, 
        DP_ff_3_, DP_ff_2_, DP_ff_1_, DP_ff_0_}), .B({DP_ff_part_23_, 
        DP_ff_part_22_, DP_ff_part_21_, DP_ff_part_20_, DP_ff_part_19_, 
        DP_ff_part_18_, DP_ff_part_17_, DP_ff_part_16_, DP_ff_part_15_, 
        DP_ff_part_14_, DP_ff_part_13_, DP_ff_part_12_, DP_ff_part_11_, 
        DP_ff_part_10_, DP_ff_part_9_, DP_ff_part_8_, DP_ff_part_7_, 
        DP_ff_part_6_, DP_ff_part_5_, DP_ff_part_4_, DP_ff_part_3_, 
        DP_ff_part_2_, DP_ff_part_1_, DP_ff_part_0_}), .SUM({DP_y_23, DP_y_11_, 
        DP_y_10_, DP_y_9_, DP_y_8_, DP_y_7_, DP_y_6_, DP_y_5_, DP_y_4_, 
        DP_y_3_, DP_y_2_, DP_y_1_, DP_y_0_, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10}), .CI(1'b0) );
  iir_filter_DW_mult_tc_0 DP_mult_206 ( .a({DP_coeffs_ff_int[0], 
        DP_coeffs_ff_int[1], n1142, DP_coeffs_ff_int[3], DP_coeffs_ff_int[4], 
        DP_coeffs_ff_int[5], n1048, DP_coeffs_ff_int[7], n1077, 
        DP_coeffs_ff_int[9], DP_coeffs_ff_int[10], DP_coeffs_ff_int[11], 
        DP_coeffs_ff_int[12], DP_coeffs_ff_int[13], DP_coeffs_ff_int[14], 
        DP_coeffs_ff_int[15], DP_coeffs_ff_int[16], DP_coeffs_ff_int[17], 
        DP_coeffs_ff_int[18], DP_coeffs_ff_int[19], n998, DP_coeffs_ff_int[21], 
        n1138, DP_coeffs_ff_int[23]}), .b({DP_pipe00[23], DP_pipe00[22], 
        DP_pipe00[21], DP_pipe00[20], DP_pipe00[19], DP_pipe00[18], 
        DP_pipe00[17], DP_pipe00[16], DP_pipe00[15], DP_pipe00[14], 
        DP_pipe00[13], DP_pipe00[12], DP_pipe00[11], DP_pipe00[10], 
        DP_pipe00[9], DP_pipe00[8], DP_pipe00[7], DP_pipe00[6], DP_pipe00[5], 
        DP_pipe00[4], DP_pipe00[3], DP_pipe00[2], DP_pipe00[1], DP_pipe00[0]}), 
        .product({DP_pipe0_coeff_pipe00[23], SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, DP_pipe0_coeff_pipe00[22], 
        DP_pipe0_coeff_pipe00[21], DP_pipe0_coeff_pipe00[20], 
        DP_pipe0_coeff_pipe00[19], DP_pipe0_coeff_pipe00[18], 
        DP_pipe0_coeff_pipe00[17], DP_pipe0_coeff_pipe00[16], 
        DP_pipe0_coeff_pipe00[15], DP_pipe0_coeff_pipe00[14], 
        DP_pipe0_coeff_pipe00[13], DP_pipe0_coeff_pipe00[12], 
        DP_pipe0_coeff_pipe00[11], DP_pipe0_coeff_pipe00[10], 
        DP_pipe0_coeff_pipe00[9], DP_pipe0_coeff_pipe00[8], 
        DP_pipe0_coeff_pipe00[7], DP_pipe0_coeff_pipe00[6], 
        DP_pipe0_coeff_pipe00[5], DP_pipe0_coeff_pipe00[4], 
        DP_pipe0_coeff_pipe00[3], DP_pipe0_coeff_pipe00[2], 
        DP_pipe0_coeff_pipe00[1], DP_pipe0_coeff_pipe00[0], 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34}) );
  iir_filter_DW_mult_tc_2 DP_mult_207 ( .a({n1095, DP_coeffs_ff_int[25], n1067, 
        DP_coeffs_ff_int[27], n1024, DP_coeffs_ff_int[29], n1026, 
        DP_coeffs_ff_int[31], n1030, DP_coeffs_ff_int[33], n1022, 
        DP_coeffs_ff_int[35], DP_coeffs_ff_int[36], DP_coeffs_ff_int[37], 
        DP_coeffs_ff_int[38], n1018, n1061, DP_coeffs_ff_int[41], n1058, 
        DP_coeffs_ff_int[43], n1054, DP_coeffs_ff_int[45], n1097, 
        DP_coeffs_ff_int[47]}), .b({DP_pipe01[23], DP_pipe01[22], 
        DP_pipe01[21], DP_pipe01[20], DP_pipe01[19], DP_pipe01[18], 
        DP_pipe01[17], DP_pipe01[16], DP_pipe01[15], DP_pipe01[14], 
        DP_pipe01[13], DP_pipe01[12], DP_pipe01[11], DP_pipe01[10], 
        DP_pipe01[9], DP_pipe01[8], DP_pipe01[7], DP_pipe01[6], DP_pipe01[5], 
        DP_pipe01[4], DP_pipe01[3], DP_pipe01[2], DP_pipe01[1], DP_pipe01[0]}), 
        .product({DP_pipe0_coeff_pipe01[23], SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, DP_pipe0_coeff_pipe01[22], 
        DP_pipe0_coeff_pipe01[21], DP_pipe0_coeff_pipe01[20], 
        DP_pipe0_coeff_pipe01[19], DP_pipe0_coeff_pipe01[18], 
        DP_pipe0_coeff_pipe01[17], DP_pipe0_coeff_pipe01[16], 
        DP_pipe0_coeff_pipe01[15], DP_pipe0_coeff_pipe01[14], 
        DP_pipe0_coeff_pipe01[13], DP_pipe0_coeff_pipe01[12], 
        DP_pipe0_coeff_pipe01[11], DP_pipe0_coeff_pipe01[10], 
        DP_pipe0_coeff_pipe01[9], DP_pipe0_coeff_pipe01[8], 
        DP_pipe0_coeff_pipe01[7], DP_pipe0_coeff_pipe01[6], 
        DP_pipe0_coeff_pipe01[5], DP_pipe0_coeff_pipe01[4], 
        DP_pipe0_coeff_pipe01[3], DP_pipe0_coeff_pipe01[2], 
        DP_pipe0_coeff_pipe01[1], DP_pipe0_coeff_pipe01[0], 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, 
        SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48, 
        SYNOPSYS_UNCONNECTED__49, SYNOPSYS_UNCONNECTED__50, 
        SYNOPSYS_UNCONNECTED__51, SYNOPSYS_UNCONNECTED__52, 
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54, 
        SYNOPSYS_UNCONNECTED__55, SYNOPSYS_UNCONNECTED__56, 
        SYNOPSYS_UNCONNECTED__57, SYNOPSYS_UNCONNECTED__58}) );
  iir_filter_DW_mult_tc_4 DP_mult_208 ( .a({n1001, DP_coeffs_ff_int[49], 
        DP_coeffs_ff_int[50], DP_coeffs_ff_int[51], n1041, 
        DP_coeffs_ff_int[53], n1007, DP_coeffs_ff_int[55], 
        DP_coeffs_ff_int[56], DP_coeffs_ff_int[57], n1045, 
        DP_coeffs_ff_int[59], n1052, DP_coeffs_ff_int[61], 
        DP_coeffs_ff_int[62], DP_coeffs_ff_int[63], n1104, 
        DP_coeffs_ff_int[65], n1110, DP_coeffs_ff_int[67], n1071, 
        DP_coeffs_ff_int[69], DP_coeffs_ff_int[70], DP_coeffs_ff_int[71]}), 
        .b({DP_pipe02[23], DP_pipe02[22], DP_pipe02[21], DP_pipe02[20], 
        DP_pipe02[19], DP_pipe02[18], DP_pipe02[17], DP_pipe02[16], 
        DP_pipe02[15], DP_pipe02[14], DP_pipe02[13], DP_pipe02[12], 
        DP_pipe02[11], DP_pipe02[10], DP_pipe02[9], DP_pipe02[8], DP_pipe02[7], 
        DP_pipe02[6], DP_pipe02[5], DP_pipe02[4], DP_pipe02[3], DP_pipe02[2], 
        DP_pipe02[1], DP_pipe02[0]}), .product({DP_pipe0_coeff_pipe02[23], 
        SYNOPSYS_UNCONNECTED__59, SYNOPSYS_UNCONNECTED__60, 
        DP_pipe0_coeff_pipe02[22], DP_pipe0_coeff_pipe02[21], 
        DP_pipe0_coeff_pipe02[20], DP_pipe0_coeff_pipe02[19], 
        DP_pipe0_coeff_pipe02[18], DP_pipe0_coeff_pipe02[17], 
        DP_pipe0_coeff_pipe02[16], DP_pipe0_coeff_pipe02[15], 
        DP_pipe0_coeff_pipe02[14], DP_pipe0_coeff_pipe02[13], 
        DP_pipe0_coeff_pipe02[12], DP_pipe0_coeff_pipe02[11], 
        DP_pipe0_coeff_pipe02[10], DP_pipe0_coeff_pipe02[9], 
        DP_pipe0_coeff_pipe02[8], DP_pipe0_coeff_pipe02[7], 
        DP_pipe0_coeff_pipe02[6], DP_pipe0_coeff_pipe02[5], 
        DP_pipe0_coeff_pipe02[4], DP_pipe0_coeff_pipe02[3], 
        DP_pipe0_coeff_pipe02[2], DP_pipe0_coeff_pipe02[1], 
        DP_pipe0_coeff_pipe02[0], SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82}) );
  iir_filter_DW_mult_tc_5 DP_mult_209 ( .a({DP_coeffs_ff_int[72], 
        DP_coeffs_ff_int[73], n1028, DP_coeffs_ff_int[75], n1075, 
        DP_coeffs_ff_int[77], n1073, DP_coeffs_ff_int[79], n1081, 
        DP_coeffs_ff_int[81], DP_coeffs_ff_int[82], DP_coeffs_ff_int[83], 
        n1020, DP_coeffs_ff_int[85], DP_coeffs_ff_int[86], 
        DP_coeffs_ff_int[87], DP_coeffs_ff_int[88], DP_coeffs_ff_int[89], 
        DP_coeffs_ff_int[90], DP_coeffs_ff_int[91], n1092, 
        DP_coeffs_ff_int[93], n1102, DP_coeffs_ff_int[95]}), .b({DP_pipe03[23], 
        DP_pipe03[22], DP_pipe03[21], DP_pipe03[20], DP_pipe03[19], 
        DP_pipe03[18], DP_pipe03[17], DP_pipe03[16], DP_pipe03[15], 
        DP_pipe03[14], DP_pipe03[13], DP_pipe03[12], DP_pipe03[11], 
        DP_pipe03[10], DP_pipe03[9], DP_pipe03[8], DP_pipe03[7], DP_pipe03[6], 
        DP_pipe03[5], DP_pipe03[4], DP_pipe03[3], DP_pipe03[2], DP_pipe03[1], 
        DP_pipe03[0]}), .product({DP_pipe0_coeff_pipe03[23], 
        SYNOPSYS_UNCONNECTED__83, SYNOPSYS_UNCONNECTED__84, 
        DP_pipe0_coeff_pipe03[22], DP_pipe0_coeff_pipe03[21], 
        DP_pipe0_coeff_pipe03[20], DP_pipe0_coeff_pipe03[19], 
        DP_pipe0_coeff_pipe03[18], DP_pipe0_coeff_pipe03[17], 
        DP_pipe0_coeff_pipe03[16], DP_pipe0_coeff_pipe03[15], 
        DP_pipe0_coeff_pipe03[14], DP_pipe0_coeff_pipe03[13], 
        DP_pipe0_coeff_pipe03[12], DP_pipe0_coeff_pipe03[11], 
        DP_pipe0_coeff_pipe03[10], DP_pipe0_coeff_pipe03[9], 
        DP_pipe0_coeff_pipe03[8], DP_pipe0_coeff_pipe03[7], 
        DP_pipe0_coeff_pipe03[6], DP_pipe0_coeff_pipe03[5], 
        DP_pipe0_coeff_pipe03[4], DP_pipe0_coeff_pipe03[3], 
        DP_pipe0_coeff_pipe03[2], DP_pipe0_coeff_pipe03[1], 
        DP_pipe0_coeff_pipe03[0], SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106}) );
  iir_filter_DW_mult_tc_1 DP_mult_204 ( .a({DP_coeffs_fb_int[0], 
        DP_coeffs_fb_int[1], n1100, DP_coeffs_fb_int[3], n1090, 
        DP_coeffs_fb_int[5], DP_coeffs_fb_int[6], DP_coeffs_fb_int[7], 
        DP_coeffs_fb_int[8], DP_coeffs_fb_int[9], n1032, n1063, n1087, 
        DP_coeffs_fb_int[13], DP_coeffs_fb_int[14], DP_coeffs_fb_int[15], 
        n1043, DP_coeffs_fb_int[17], n1106, DP_coeffs_fb_int[19], n1079, 
        DP_coeffs_fb_int[21], n1108, DP_coeffs_fb_int[23]}), .b({n1056, n1065, 
        DP_sw0_21_, DP_sw0_20_, DP_sw0_19_, DP_sw0_18_, DP_sw0_17_, DP_sw0_16_, 
        DP_sw0_15_, DP_sw0_14_, DP_sw0_13_, DP_sw0_12_, DP_sw0_11_, DP_sw0_10_, 
        DP_sw0_9_, DP_sw0_8_, DP_sw0_7_, DP_sw0_6_, DP_sw0_5_, DP_sw0_4_, 
        DP_sw0_3_, DP_sw0_2_, DP_sw0_1_, DP_sw0_0_}), .product({
        DP_sw0_coeff_ret0[23], SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, DP_sw0_coeff_ret0[22], 
        DP_sw0_coeff_ret0[21], DP_sw0_coeff_ret0[20], DP_sw0_coeff_ret0[19], 
        DP_sw0_coeff_ret0[18], DP_sw0_coeff_ret0[17], DP_sw0_coeff_ret0[16], 
        DP_sw0_coeff_ret0[15], DP_sw0_coeff_ret0[14], DP_sw0_coeff_ret0[13], 
        DP_sw0_coeff_ret0[12], DP_sw0_coeff_ret0[11], DP_sw0_coeff_ret0[10], 
        DP_sw0_coeff_ret0[9], DP_sw0_coeff_ret0[8], DP_sw0_coeff_ret0[7], 
        DP_sw0_coeff_ret0[6], DP_sw0_coeff_ret0[5], DP_sw0_coeff_ret0[4], 
        DP_sw0_coeff_ret0[3], DP_sw0_coeff_ret0[2], DP_sw0_coeff_ret0[1], 
        DP_sw0_coeff_ret0[0], SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130}) );
  iir_filter_DW_mult_tc_3 DP_mult_205 ( .a({DP_coeffs_fb_int[24], 
        DP_coeffs_fb_int[25], DP_coeffs_fb_int[26], DP_coeffs_fb_int[27], 
        DP_coeffs_fb_int[28], DP_coeffs_fb_int[29], DP_coeffs_fb_int[30], 
        DP_coeffs_fb_int[31], DP_coeffs_fb_int[32], DP_coeffs_fb_int[33], 
        n1009, DP_coeffs_fb_int[35], n1005, DP_coeffs_fb_int[37], n1140, 
        DP_coeffs_fb_int[39], n1085, DP_coeffs_fb_int[41], 
        DP_coeffs_fb_int[42], DP_coeffs_fb_int[43], DP_coeffs_fb_int[44], 
        DP_coeffs_fb_int[45], DP_coeffs_fb_int[46], DP_coeffs_fb_int[47]}), 
        .b({DP_sw1_23_, DP_sw1_22_, DP_sw1_21_, DP_sw1_20_, DP_sw1_19_, 
        DP_sw1_18_, DP_sw1_17_, DP_sw1_16_, DP_sw1_15_, DP_sw1_14_, DP_sw1_13_, 
        DP_sw1_12_, DP_sw1_11_, DP_sw1_10_, DP_sw1_9_, DP_sw1_8_, DP_sw1_7_, 
        DP_sw1_6_, DP_sw1_5_, DP_sw1_4_, DP_sw1_3_, DP_sw1_2_, DP_sw1_1_, 
        n1069}), .product({DP_sw1_coeff_ret1[23], SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, DP_sw1_coeff_ret1[22], 
        DP_sw1_coeff_ret1[21], DP_sw1_coeff_ret1[20], DP_sw1_coeff_ret1[19], 
        DP_sw1_coeff_ret1[18], DP_sw1_coeff_ret1[17], DP_sw1_coeff_ret1[16], 
        DP_sw1_coeff_ret1[15], DP_sw1_coeff_ret1[14], DP_sw1_coeff_ret1[13], 
        DP_sw1_coeff_ret1[12], DP_sw1_coeff_ret1[11], DP_sw1_coeff_ret1[10], 
        DP_sw1_coeff_ret1[9], DP_sw1_coeff_ret1[8], DP_sw1_coeff_ret1[7], 
        DP_sw1_coeff_ret1[6], DP_sw1_coeff_ret1[5], DP_sw1_coeff_ret1[4], 
        DP_sw1_coeff_ret1[3], DP_sw1_coeff_ret1[2], DP_sw1_coeff_ret1[1], 
        DP_sw1_coeff_ret1[0], SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154}) );
  DFFR_X1 DP_reg_ret1_Q_reg_13_ ( .D(DP_sw1_coeff_ret1[13]), .CK(clk), .RN(
        n1189), .Q(DP_ret1[13]) );
  DFFR_X1 DP_reg_ret1_Q_reg_18_ ( .D(DP_sw1_coeff_ret1[18]), .CK(clk), .RN(
        n1189), .Q(DP_ret1[18]) );
  DFFR_X1 DP_reg_ret1_Q_reg_15_ ( .D(DP_sw1_coeff_ret1[15]), .CK(clk), .RN(
        n1189), .Q(DP_ret1[15]) );
  DFFR_X2 DP_reg_sw0_Q_reg_0_ ( .D(n1447), .CK(clk), .RN(n1203), .Q(DP_sw0_0_)
         );
  DFFR_X2 DP_reg_pipe02_Q_reg_0_ ( .D(DP_sw1_0_), .CK(clk), .RN(n1208), .Q(
        DP_pipe02[0]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_15_ ( .D(DP_pipe0_coeff_pipe00[15]), .CK(clk), 
        .RN(n1193), .Q(DP_pipe10[15]) );
  DFFR_X2 DP_reg_pipe03_Q_reg_0_ ( .D(n1236), .CK(clk), .RN(n1212), .Q(
        DP_pipe03[0]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_18_ ( .D(DP_pipe0_coeff_pipe00[18]), .CK(clk), 
        .RN(n1193), .Q(DP_pipe10[18]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_20_ ( .D(DP_pipe0_coeff_pipe03[20]), .CK(clk), 
        .RN(n1199), .Q(DP_pipe13[20]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_21_ ( .D(DP_pipe0_coeff_pipe03[21]), .CK(clk), 
        .RN(n1199), .Q(DP_pipe13[21]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_19_ ( .D(DP_pipe0_coeff_pipe03[19]), .CK(clk), 
        .RN(n1199), .Q(DP_pipe13[19]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_14_ ( .D(DP_pipe0_coeff_pipe03[14]), .CK(clk), 
        .RN(n1199), .Q(DP_pipe13[14]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_16_ ( .D(DP_pipe0_coeff_pipe03[16]), .CK(clk), 
        .RN(n1199), .Q(DP_pipe13[16]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_17_ ( .D(DP_pipe0_coeff_pipe03[17]), .CK(clk), 
        .RN(n1199), .Q(DP_pipe13[17]) );
  DFFR_X2 DP_reg_pipe01_Q_reg_14_ ( .D(DP_sw0_14_), .CK(clk), .RN(n1201), .Q(
        DP_pipe01[14]) );
  DFFR_X1 DP_reg_ret1_Q_reg_19_ ( .D(DP_sw1_coeff_ret1[19]), .CK(clk), .RN(
        n1189), .Q(DP_ret1[19]) );
  DFFR_X1 DP_reg_ret1_Q_reg_20_ ( .D(DP_sw1_coeff_ret1[20]), .CK(clk), .RN(
        n1189), .Q(DP_ret1[20]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_20_ ( .D(DP_pipe0_coeff_pipe02[20]), .CK(clk), 
        .RN(n1197), .Q(DP_pipe12[20]) );
  DFFR_X1 DP_reg_ret1_Q_reg_9_ ( .D(DP_sw1_coeff_ret1[9]), .CK(clk), .RN(n1188), .Q(DP_ret1[9]) );
  DFFR_X1 DP_reg_ret1_Q_reg_16_ ( .D(DP_sw1_coeff_ret1[16]), .CK(clk), .RN(
        n1189), .Q(DP_ret1[16]) );
  DFFR_X2 DP_reg_pipe11_Q_reg_17_ ( .D(DP_pipe0_coeff_pipe01[17]), .CK(clk), 
        .RN(n1195), .Q(DP_pipe11[17]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_13_ ( .D(DP_pipe0_coeff_pipe01[13]), .CK(clk), 
        .RN(n1195), .Q(DP_pipe11[13]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_14_ ( .D(DP_pipe0_coeff_pipe01[14]), .CK(clk), 
        .RN(n1195), .Q(DP_pipe11[14]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_18_ ( .D(DP_pipe0_coeff_pipe01[18]), .CK(clk), 
        .RN(n1195), .Q(DP_pipe11[18]) );
  DFFR_X1 DP_reg_ret1_Q_reg_22_ ( .D(DP_sw1_coeff_ret1[22]), .CK(clk), .RN(
        n1189), .Q(DP_ret1[22]) );
  DFFR_X2 DP_reg_sw1_Q_reg_8_ ( .D(n1463), .CK(clk), .RN(n1206), .Q(DP_sw1_8_)
         );
  DFFR_X1 DP_reg_pipe13_Q_reg_15_ ( .D(DP_pipe0_coeff_pipe03[15]), .CK(clk), 
        .RN(n1199), .Q(DP_pipe13[15]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_18_ ( .D(DP_pipe0_coeff_pipe03[18]), .CK(clk), 
        .RN(n1199), .Q(DP_pipe13[18]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_13_ ( .D(DP_pipe0_coeff_pipe03[13]), .CK(clk), 
        .RN(n1199), .Q(DP_pipe13[13]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_16_ ( .D(DP_pipe0_coeff_pipe01[16]), .CK(clk), 
        .RN(n1195), .Q(DP_pipe11[16]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_22_ ( .D(DP_pipe0_coeff_pipe01[22]), .CK(clk), 
        .RN(n1195), .Q(DP_pipe11[22]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_22_ ( .D(DP_pipe0_coeff_pipe03[22]), .CK(clk), 
        .RN(n1199), .Q(DP_pipe13[22]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_20_ ( .D(DP_pipe0_coeff_pipe01[20]), .CK(clk), 
        .RN(n1195), .Q(DP_pipe11[20]) );
  DFFR_X2 DP_reg_pipe11_Q_reg_19_ ( .D(DP_pipe0_coeff_pipe01[19]), .CK(clk), 
        .RN(n1195), .Q(DP_pipe11[19]) );
  DFFR_X2 DP_reg_pipe10_Q_reg_20_ ( .D(DP_pipe0_coeff_pipe00[20]), .CK(clk), 
        .RN(n1193), .Q(DP_pipe10[20]) );
  DFFR_X2 DP_reg_pipe10_Q_reg_19_ ( .D(DP_pipe0_coeff_pipe00[19]), .CK(clk), 
        .RN(n1193), .Q(DP_pipe10[19]) );
  DFFR_X2 DP_reg_pipe10_Q_reg_22_ ( .D(DP_pipe0_coeff_pipe00[22]), .CK(clk), 
        .RN(n1193), .Q(DP_pipe10[22]) );
  DFFR_X2 DP_reg_pipe10_Q_reg_16_ ( .D(DP_pipe0_coeff_pipe00[16]), .CK(clk), 
        .RN(n1193), .Q(DP_pipe10[16]) );
  DFFR_X2 DP_reg_pipe10_Q_reg_17_ ( .D(DP_pipe0_coeff_pipe00[17]), .CK(clk), 
        .RN(n1193), .Q(DP_pipe10[17]) );
  DFFR_X2 DP_reg_pipe10_Q_reg_14_ ( .D(DP_pipe0_coeff_pipe00[14]), .CK(clk), 
        .RN(n1193), .Q(DP_pipe10[14]) );
  DFFR_X2 DP_reg_pipe10_Q_reg_13_ ( .D(DP_pipe0_coeff_pipe00[13]), .CK(clk), 
        .RN(n1193), .Q(DP_pipe10[13]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_15_ ( .D(DP_pipe0_coeff_pipe01[15]), .CK(clk), 
        .RN(n1195), .Q(DP_pipe11[15]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_21_ ( .D(DP_pipe0_coeff_pipe01[21]), .CK(clk), 
        .RN(n1195), .Q(DP_pipe11[21]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_12_ ( .D(DP_pipe0_coeff_pipe01[12]), .CK(clk), 
        .RN(n1195), .Q(DP_pipe11[12]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_21_ ( .D(DP_pipe0_coeff_pipe00[21]), .CK(clk), 
        .RN(n1193), .Q(DP_pipe10[21]) );
  INV_X1 U494 ( .A(n997), .ZN(n998) );
  INV_X1 U495 ( .A(n1000), .ZN(n1001) );
  INV_X1 U496 ( .A(n1004), .ZN(n1005) );
  INV_X1 U497 ( .A(n1006), .ZN(n1007) );
  INV_X1 U498 ( .A(n1008), .ZN(n1009) );
  INV_X1 U499 ( .A(n1017), .ZN(n1018) );
  INV_X1 U500 ( .A(n1019), .ZN(n1020) );
  INV_X1 U501 ( .A(n1021), .ZN(n1022) );
  INV_X1 U502 ( .A(n1023), .ZN(n1024) );
  INV_X1 U503 ( .A(n1025), .ZN(n1026) );
  INV_X1 U504 ( .A(n1027), .ZN(n1028) );
  INV_X1 U505 ( .A(n1029), .ZN(n1030) );
  INV_X1 U506 ( .A(n1031), .ZN(n1032) );
  INV_X2 U507 ( .A(n1089), .ZN(n1090) );
  CLKBUF_X3 U508 ( .A(n1234), .Z(n1034) );
  OAI21_X1 U509 ( .B1(DP_y_11_), .B2(n1221), .A(delayed_controls_2__0_), .ZN(
        n1234) );
  NAND3_X2 U510 ( .A1(DP_y_11_), .A2(delayed_controls_2__0_), .A3(n1221), .ZN(
        n1232) );
  INV_X1 U511 ( .A(n1037), .ZN(n1038) );
  INV_X1 U512 ( .A(n1040), .ZN(n1041) );
  INV_X1 U513 ( .A(n1042), .ZN(n1043) );
  INV_X1 U514 ( .A(n1044), .ZN(n1045) );
  INV_X1 U515 ( .A(n1047), .ZN(n1048) );
  INV_X1 U516 ( .A(n1051), .ZN(n1052) );
  INV_X2 U517 ( .A(n1080), .ZN(n1081) );
  INV_X1 U518 ( .A(n1053), .ZN(n1054) );
  INV_X2 U519 ( .A(n1055), .ZN(n1056) );
  INV_X1 U520 ( .A(n1057), .ZN(n1058) );
  INV_X1 U521 ( .A(n1060), .ZN(n1061) );
  INV_X1 U522 ( .A(n1062), .ZN(n1063) );
  INV_X2 U523 ( .A(n1064), .ZN(n1065) );
  INV_X1 U524 ( .A(n1066), .ZN(n1067) );
  INV_X2 U525 ( .A(n1068), .ZN(n1069) );
  INV_X1 U526 ( .A(n1070), .ZN(n1071) );
  INV_X2 U527 ( .A(n1072), .ZN(n1073) );
  INV_X1 U528 ( .A(n1074), .ZN(n1075) );
  INV_X1 U529 ( .A(n1076), .ZN(n1077) );
  INV_X1 U530 ( .A(n1078), .ZN(n1079) );
  INV_X1 U531 ( .A(n1084), .ZN(n1085) );
  INV_X1 U532 ( .A(n1086), .ZN(n1087) );
  INV_X1 U533 ( .A(n1091), .ZN(n1092) );
  INV_X1 U534 ( .A(n1094), .ZN(n1095) );
  INV_X1 U535 ( .A(n1096), .ZN(n1097) );
  INV_X1 U536 ( .A(n1099), .ZN(n1100) );
  INV_X1 U537 ( .A(n1101), .ZN(n1102) );
  INV_X1 U538 ( .A(n1103), .ZN(n1104) );
  INV_X1 U539 ( .A(n1105), .ZN(n1106) );
  INV_X1 U540 ( .A(n1107), .ZN(n1108) );
  INV_X1 U541 ( .A(n1109), .ZN(n1110) );
  XOR2_X1 U542 ( .A(n1124), .B(n1112), .Z(n1261) );
  MUX2_X1 U543 ( .A(DP_x[0]), .B(dIn[0]), .S(n1170), .Z(n1268) );
  BUF_X1 U544 ( .A(n1151), .Z(n1154) );
  BUF_X1 U545 ( .A(n1151), .Z(n1155) );
  BUF_X1 U546 ( .A(n1152), .Z(n1156) );
  BUF_X1 U547 ( .A(n1151), .Z(n1153) );
  BUF_X1 U548 ( .A(n1152), .Z(n1157) );
  BUF_X1 U549 ( .A(n1260), .Z(n1151) );
  BUF_X1 U550 ( .A(n1260), .Z(n1152) );
  BUF_X1 U551 ( .A(n1171), .Z(n1161) );
  BUF_X1 U552 ( .A(n1172), .Z(n1158) );
  CLKBUF_X3 U553 ( .A(n1171), .Z(n1165) );
  BUF_X1 U554 ( .A(n1171), .Z(n1162) );
  BUF_X1 U555 ( .A(n1171), .Z(n1163) );
  BUF_X1 U556 ( .A(n1171), .Z(n1164) );
  CLKBUF_X3 U557 ( .A(n1170), .Z(n1168) );
  BUF_X1 U558 ( .A(n1170), .Z(n1169) );
  BUF_X1 U559 ( .A(n1170), .Z(n1166) );
  BUF_X1 U560 ( .A(n1170), .Z(n1167) );
  BUF_X1 U561 ( .A(n1172), .Z(n1159) );
  BUF_X1 U562 ( .A(n1172), .Z(n1160) );
  NAND2_X1 U563 ( .A1(n1123), .A2(dOut[0]), .ZN(n1113) );
  NAND2_X1 U564 ( .A1(n1123), .A2(dOut[1]), .ZN(n1114) );
  NAND2_X1 U565 ( .A1(n1123), .A2(dOut[2]), .ZN(n1115) );
  NAND2_X1 U566 ( .A1(n1123), .A2(dOut[3]), .ZN(n1116) );
  NAND2_X1 U567 ( .A1(n1123), .A2(dOut[4]), .ZN(n1117) );
  NAND2_X1 U568 ( .A1(n1123), .A2(dOut[5]), .ZN(n1118) );
  NAND2_X1 U569 ( .A1(n1123), .A2(dOut[6]), .ZN(n1119) );
  NAND2_X1 U570 ( .A1(n1123), .A2(dOut[7]), .ZN(n1120) );
  NAND2_X1 U571 ( .A1(n1123), .A2(dOut[8]), .ZN(n1121) );
  NAND2_X1 U572 ( .A1(n1123), .A2(dOut[9]), .ZN(n1122) );
  BUF_X1 U573 ( .A(vIn), .Z(n1172) );
  BUF_X1 U574 ( .A(rst_n), .Z(n1214) );
  BUF_X1 U575 ( .A(rst_n), .Z(n1215) );
  BUF_X1 U576 ( .A(rst_n), .Z(n1216) );
  BUF_X1 U577 ( .A(rst_n), .Z(n1217) );
  BUF_X1 U578 ( .A(rst_n), .Z(n1218) );
  BUF_X1 U579 ( .A(rst_n), .Z(n1219) );
  BUF_X1 U580 ( .A(rst_n), .Z(n1220) );
  INV_X1 U581 ( .A(n1137), .ZN(n1138) );
  INV_X1 U582 ( .A(n1139), .ZN(n1140) );
  INV_X1 U583 ( .A(n1141), .ZN(n1142) );
  CLKBUF_X2 U584 ( .A(vIn), .Z(n1170) );
  CLKBUF_X2 U585 ( .A(vIn), .Z(n1171) );
  CLKBUF_X1 U586 ( .A(n1220), .Z(n1173) );
  CLKBUF_X1 U587 ( .A(n1220), .Z(n1174) );
  CLKBUF_X1 U588 ( .A(n1220), .Z(n1175) );
  CLKBUF_X1 U589 ( .A(n1220), .Z(n1176) );
  CLKBUF_X1 U590 ( .A(n1220), .Z(n1177) );
  CLKBUF_X1 U591 ( .A(n1219), .Z(n1178) );
  CLKBUF_X1 U592 ( .A(n1219), .Z(n1179) );
  CLKBUF_X1 U593 ( .A(n1219), .Z(n1180) );
  CLKBUF_X1 U594 ( .A(n1219), .Z(n1181) );
  CLKBUF_X1 U595 ( .A(n1219), .Z(n1182) );
  CLKBUF_X1 U596 ( .A(n1219), .Z(n1183) );
  CLKBUF_X1 U597 ( .A(n1218), .Z(n1184) );
  CLKBUF_X1 U598 ( .A(n1218), .Z(n1185) );
  CLKBUF_X1 U599 ( .A(n1218), .Z(n1186) );
  CLKBUF_X1 U600 ( .A(n1218), .Z(n1187) );
  CLKBUF_X1 U601 ( .A(n1218), .Z(n1188) );
  CLKBUF_X1 U602 ( .A(n1218), .Z(n1189) );
  CLKBUF_X1 U603 ( .A(n1217), .Z(n1190) );
  CLKBUF_X1 U604 ( .A(n1217), .Z(n1191) );
  CLKBUF_X1 U605 ( .A(n1217), .Z(n1192) );
  CLKBUF_X1 U606 ( .A(n1217), .Z(n1193) );
  CLKBUF_X1 U607 ( .A(n1217), .Z(n1194) );
  CLKBUF_X1 U608 ( .A(n1217), .Z(n1195) );
  CLKBUF_X1 U609 ( .A(n1216), .Z(n1196) );
  CLKBUF_X1 U610 ( .A(n1216), .Z(n1197) );
  CLKBUF_X1 U611 ( .A(n1216), .Z(n1198) );
  CLKBUF_X1 U612 ( .A(n1216), .Z(n1199) );
  CLKBUF_X1 U613 ( .A(n1216), .Z(n1200) );
  CLKBUF_X1 U614 ( .A(n1216), .Z(n1201) );
  CLKBUF_X1 U615 ( .A(n1215), .Z(n1202) );
  CLKBUF_X1 U616 ( .A(n1215), .Z(n1203) );
  CLKBUF_X1 U617 ( .A(n1215), .Z(n1204) );
  CLKBUF_X1 U618 ( .A(n1215), .Z(n1205) );
  CLKBUF_X1 U619 ( .A(n1215), .Z(n1206) );
  CLKBUF_X1 U620 ( .A(n1215), .Z(n1207) );
  CLKBUF_X1 U621 ( .A(n1214), .Z(n1208) );
  CLKBUF_X1 U622 ( .A(n1214), .Z(n1209) );
  CLKBUF_X1 U623 ( .A(n1214), .Z(n1210) );
  CLKBUF_X1 U624 ( .A(n1214), .Z(n1211) );
  CLKBUF_X1 U625 ( .A(n1214), .Z(n1212) );
  CLKBUF_X1 U626 ( .A(n1214), .Z(n1213) );
  INV_X1 U627 ( .A(DP_y_23), .ZN(n1221) );
  INV_X1 U628 ( .A(DP_y_0_), .ZN(n1222) );
  OAI211_X1 U629 ( .C1(n1034), .C2(n1222), .A(n1232), .B(n1113), .ZN(n513) );
  INV_X1 U630 ( .A(DP_y_1_), .ZN(n1223) );
  OAI211_X1 U631 ( .C1(n1034), .C2(n1223), .A(n1232), .B(n1114), .ZN(n514) );
  INV_X1 U632 ( .A(DP_y_2_), .ZN(n1224) );
  OAI211_X1 U633 ( .C1(n1034), .C2(n1224), .A(n1232), .B(n1115), .ZN(n515) );
  INV_X1 U634 ( .A(DP_y_3_), .ZN(n1225) );
  OAI211_X1 U635 ( .C1(n1034), .C2(n1225), .A(n1232), .B(n1116), .ZN(n516) );
  INV_X1 U636 ( .A(DP_y_4_), .ZN(n1226) );
  OAI211_X1 U637 ( .C1(n1034), .C2(n1226), .A(n1232), .B(n1117), .ZN(n517) );
  INV_X1 U638 ( .A(DP_y_5_), .ZN(n1227) );
  OAI211_X1 U639 ( .C1(n1034), .C2(n1227), .A(n1232), .B(n1118), .ZN(n518) );
  INV_X1 U640 ( .A(DP_y_6_), .ZN(n1228) );
  OAI211_X1 U641 ( .C1(n1034), .C2(n1228), .A(n1232), .B(n1119), .ZN(n519) );
  INV_X1 U642 ( .A(DP_y_7_), .ZN(n1229) );
  OAI211_X1 U643 ( .C1(n1034), .C2(n1229), .A(n1232), .B(n1120), .ZN(n520) );
  INV_X1 U644 ( .A(DP_y_8_), .ZN(n1230) );
  OAI211_X1 U645 ( .C1(n1034), .C2(n1230), .A(n1232), .B(n1121), .ZN(n521) );
  INV_X1 U646 ( .A(DP_y_9_), .ZN(n1231) );
  OAI211_X1 U647 ( .C1(n1034), .C2(n1231), .A(n1232), .B(n1122), .ZN(n522) );
  INV_X1 U648 ( .A(DP_y_10_), .ZN(n1233) );
  OAI221_X1 U649 ( .B1(delayed_controls_2__0_), .B2(n280), .C1(n1034), .C2(
        n1233), .A(n1232), .ZN(n523) );
  MUX2_X1 U650 ( .A(dOut[11]), .B(DP_y_23), .S(delayed_controls_2__0_), .Z(
        n524) );
  INV_X1 U651 ( .A(n1261), .ZN(n1260) );
  XNOR2_X1 U652 ( .A(n1158), .B(n1153), .ZN(CU_nextState_0_) );
  MUX2_X1 U653 ( .A(DP_sw1_0_), .B(n1236), .S(n1153), .Z(n529) );
  MUX2_X1 U654 ( .A(DP_sw1_1_), .B(n1237), .S(n1153), .Z(n531) );
  MUX2_X1 U655 ( .A(DP_sw1_2_), .B(n1238), .S(n1153), .Z(n533) );
  MUX2_X1 U656 ( .A(DP_sw1_3_), .B(n1239), .S(n1153), .Z(n535) );
  MUX2_X1 U657 ( .A(DP_sw1_4_), .B(n1240), .S(n1153), .Z(n537) );
  MUX2_X1 U658 ( .A(DP_sw1_5_), .B(n1241), .S(n1153), .Z(n539) );
  MUX2_X1 U659 ( .A(DP_sw1_6_), .B(n1242), .S(n1153), .Z(n541) );
  MUX2_X1 U660 ( .A(DP_sw1_7_), .B(n1243), .S(n1153), .Z(n543) );
  MUX2_X1 U661 ( .A(DP_sw1_8_), .B(n1244), .S(n1153), .Z(n545) );
  MUX2_X1 U662 ( .A(DP_sw1_9_), .B(n1245), .S(n1153), .Z(n547) );
  MUX2_X1 U663 ( .A(DP_sw1_10_), .B(n1246), .S(n1153), .Z(n549) );
  MUX2_X1 U664 ( .A(DP_sw1_11_), .B(n1247), .S(n1153), .Z(n551) );
  MUX2_X1 U665 ( .A(DP_sw1_12_), .B(n1248), .S(n1153), .Z(n553) );
  MUX2_X1 U666 ( .A(DP_sw1_13_), .B(n1249), .S(n1154), .Z(n555) );
  MUX2_X1 U667 ( .A(DP_sw1_14_), .B(n1250), .S(n1154), .Z(n557) );
  MUX2_X1 U668 ( .A(DP_sw1_15_), .B(n1251), .S(n1154), .Z(n559) );
  MUX2_X1 U669 ( .A(DP_sw1_16_), .B(n1252), .S(n1154), .Z(n561) );
  MUX2_X1 U670 ( .A(DP_sw1_17_), .B(n1253), .S(n1154), .Z(n563) );
  MUX2_X1 U671 ( .A(DP_sw1_18_), .B(n1254), .S(n1154), .Z(n565) );
  MUX2_X1 U672 ( .A(DP_sw1_19_), .B(n1255), .S(n1154), .Z(n567) );
  MUX2_X1 U673 ( .A(DP_sw1_20_), .B(n1256), .S(n1154), .Z(n569) );
  MUX2_X1 U674 ( .A(DP_sw1_21_), .B(n1257), .S(n1154), .Z(n571) );
  MUX2_X1 U675 ( .A(DP_sw1_22_), .B(n1258), .S(n1154), .Z(n573) );
  MUX2_X1 U676 ( .A(DP_sw1_23_), .B(n1259), .S(n1154), .Z(n575) );
  MUX2_X1 U677 ( .A(DP_sw0_0_), .B(DP_sw1_0_), .S(n1154), .Z(n1471) );
  MUX2_X1 U678 ( .A(DP_sw0_1_), .B(DP_sw1_1_), .S(n1154), .Z(n1470) );
  MUX2_X1 U679 ( .A(DP_sw0_2_), .B(DP_sw1_2_), .S(n1154), .Z(n1469) );
  MUX2_X1 U680 ( .A(DP_sw0_3_), .B(DP_sw1_3_), .S(n1154), .Z(n1468) );
  MUX2_X1 U681 ( .A(DP_sw0_4_), .B(DP_sw1_4_), .S(n1155), .Z(n1467) );
  MUX2_X1 U682 ( .A(DP_sw0_5_), .B(DP_sw1_5_), .S(n1155), .Z(n1466) );
  MUX2_X1 U683 ( .A(DP_sw0_6_), .B(DP_sw1_6_), .S(n1155), .Z(n1465) );
  MUX2_X1 U684 ( .A(DP_sw0_7_), .B(DP_sw1_7_), .S(n1155), .Z(n1464) );
  MUX2_X1 U685 ( .A(DP_sw0_8_), .B(DP_sw1_8_), .S(n1155), .Z(n1463) );
  MUX2_X1 U686 ( .A(DP_sw0_9_), .B(DP_sw1_9_), .S(n1155), .Z(n1462) );
  MUX2_X1 U687 ( .A(DP_sw0_10_), .B(DP_sw1_10_), .S(n1155), .Z(n1461) );
  MUX2_X1 U688 ( .A(DP_sw0_11_), .B(DP_sw1_11_), .S(n1155), .Z(n1460) );
  MUX2_X1 U689 ( .A(DP_sw0_12_), .B(DP_sw1_12_), .S(n1155), .Z(n1459) );
  MUX2_X1 U690 ( .A(DP_sw0_13_), .B(DP_sw1_13_), .S(n1155), .Z(n1458) );
  MUX2_X1 U691 ( .A(DP_sw0_14_), .B(DP_sw1_14_), .S(n1155), .Z(n1457) );
  MUX2_X1 U692 ( .A(DP_sw0_15_), .B(DP_sw1_15_), .S(n1155), .Z(n1456) );
  MUX2_X1 U693 ( .A(DP_sw0_16_), .B(DP_sw1_16_), .S(n1155), .Z(n1455) );
  MUX2_X1 U694 ( .A(DP_sw0_17_), .B(DP_sw1_17_), .S(n1155), .Z(n1454) );
  MUX2_X1 U695 ( .A(DP_sw0_18_), .B(DP_sw1_18_), .S(n1155), .Z(n1453) );
  MUX2_X1 U696 ( .A(DP_sw0_19_), .B(DP_sw1_19_), .S(n1156), .Z(n1452) );
  MUX2_X1 U697 ( .A(DP_sw0_20_), .B(DP_sw1_20_), .S(n1156), .Z(n1451) );
  MUX2_X1 U698 ( .A(DP_sw0_21_), .B(DP_sw1_21_), .S(n1156), .Z(n1450) );
  MUX2_X1 U699 ( .A(DP_sw0_22_), .B(DP_sw1_22_), .S(n1156), .Z(n1449) );
  MUX2_X1 U700 ( .A(DP_sw0_23_), .B(DP_sw1_23_), .S(n1156), .Z(n1448) );
  MUX2_X1 U701 ( .A(DP_w_0_), .B(DP_sw0_0_), .S(n1156), .Z(n1447) );
  MUX2_X1 U702 ( .A(DP_w_1_), .B(DP_sw0_1_), .S(n1156), .Z(n1446) );
  MUX2_X1 U703 ( .A(DP_w_2_), .B(DP_sw0_2_), .S(n1156), .Z(n1445) );
  MUX2_X1 U704 ( .A(DP_w_3_), .B(DP_sw0_3_), .S(n1156), .Z(n1444) );
  MUX2_X1 U705 ( .A(DP_w_4_), .B(DP_sw0_4_), .S(n1156), .Z(n1443) );
  MUX2_X1 U706 ( .A(DP_w_5_), .B(DP_sw0_5_), .S(n1156), .Z(n1442) );
  MUX2_X1 U707 ( .A(DP_w_6_), .B(DP_sw0_6_), .S(n1156), .Z(n1441) );
  MUX2_X1 U708 ( .A(DP_w_7_), .B(DP_sw0_7_), .S(n1156), .Z(n1440) );
  MUX2_X1 U709 ( .A(DP_w_8_), .B(DP_sw0_8_), .S(n1156), .Z(n1439) );
  MUX2_X1 U710 ( .A(DP_w_9_), .B(DP_sw0_9_), .S(n1156), .Z(n1438) );
  MUX2_X1 U711 ( .A(DP_w_10_), .B(DP_sw0_10_), .S(n1157), .Z(n1437) );
  MUX2_X1 U712 ( .A(DP_w_11_), .B(DP_sw0_11_), .S(n1157), .Z(n1436) );
  MUX2_X1 U713 ( .A(DP_w_12_), .B(DP_sw0_12_), .S(n1157), .Z(n1435) );
  MUX2_X1 U714 ( .A(DP_w_13_), .B(DP_sw0_13_), .S(n1157), .Z(n1434) );
  MUX2_X1 U715 ( .A(DP_w_14_), .B(DP_sw0_14_), .S(n1157), .Z(n1433) );
  MUX2_X1 U716 ( .A(DP_w_15_), .B(DP_sw0_15_), .S(n1157), .Z(n1432) );
  MUX2_X1 U717 ( .A(DP_w_16_), .B(DP_sw0_16_), .S(n1157), .Z(n1431) );
  MUX2_X1 U718 ( .A(DP_w_17_), .B(DP_sw0_17_), .S(n1157), .Z(n1430) );
  MUX2_X1 U719 ( .A(DP_w_18_), .B(DP_sw0_18_), .S(n1157), .Z(n1429) );
  MUX2_X1 U720 ( .A(DP_w_19_), .B(DP_sw0_19_), .S(n1157), .Z(n1428) );
  MUX2_X1 U721 ( .A(DP_w_20_), .B(DP_sw0_20_), .S(n1157), .Z(n1427) );
  MUX2_X1 U722 ( .A(DP_w_21_), .B(DP_sw0_21_), .S(n1157), .Z(n1426) );
  MUX2_X1 U723 ( .A(DP_w_22_), .B(DP_sw0_22_), .S(n1157), .Z(n1425) );
  MUX2_X1 U724 ( .A(DP_w_23_), .B(DP_sw0_23_), .S(n1157), .Z(n1424) );
  MUX2_X1 U725 ( .A(DP_coeffs_ff_int[72]), .B(coeffs_ff[23]), .S(n1158), .Z(
        n1423) );
  MUX2_X1 U726 ( .A(DP_coeffs_ff_int[73]), .B(coeffs_ff[22]), .S(n1158), .Z(
        n1422) );
  MUX2_X1 U727 ( .A(DP_coeffs_ff_int[74]), .B(coeffs_ff[21]), .S(n1158), .Z(
        n1421) );
  MUX2_X1 U728 ( .A(DP_coeffs_ff_int[75]), .B(coeffs_ff[20]), .S(n1158), .Z(
        n1420) );
  MUX2_X1 U729 ( .A(DP_coeffs_ff_int[76]), .B(coeffs_ff[19]), .S(n1158), .Z(
        n1419) );
  MUX2_X1 U730 ( .A(DP_coeffs_ff_int[77]), .B(coeffs_ff[18]), .S(n1158), .Z(
        n1418) );
  MUX2_X1 U731 ( .A(DP_coeffs_ff_int[78]), .B(coeffs_ff[17]), .S(n1158), .Z(
        n1417) );
  MUX2_X1 U732 ( .A(DP_coeffs_ff_int[79]), .B(coeffs_ff[16]), .S(n1158), .Z(
        n1416) );
  MUX2_X1 U733 ( .A(DP_coeffs_ff_int[80]), .B(coeffs_ff[15]), .S(n1158), .Z(
        n1415) );
  MUX2_X1 U734 ( .A(DP_coeffs_ff_int[81]), .B(coeffs_ff[14]), .S(n1158), .Z(
        n1414) );
  MUX2_X1 U735 ( .A(DP_coeffs_ff_int[82]), .B(coeffs_ff[13]), .S(n1158), .Z(
        n1413) );
  MUX2_X1 U736 ( .A(DP_coeffs_ff_int[83]), .B(coeffs_ff[12]), .S(n1158), .Z(
        n1412) );
  MUX2_X1 U737 ( .A(DP_coeffs_ff_int[84]), .B(coeffs_ff[11]), .S(n1159), .Z(
        n1411) );
  MUX2_X1 U738 ( .A(DP_coeffs_ff_int[85]), .B(coeffs_ff[10]), .S(n1159), .Z(
        n1410) );
  MUX2_X1 U739 ( .A(DP_coeffs_ff_int[86]), .B(coeffs_ff[9]), .S(n1159), .Z(
        n1409) );
  MUX2_X1 U740 ( .A(DP_coeffs_ff_int[87]), .B(coeffs_ff[8]), .S(n1159), .Z(
        n1408) );
  MUX2_X1 U741 ( .A(DP_coeffs_ff_int[88]), .B(coeffs_ff[7]), .S(n1159), .Z(
        n1407) );
  MUX2_X1 U742 ( .A(DP_coeffs_ff_int[89]), .B(coeffs_ff[6]), .S(n1159), .Z(
        n1406) );
  MUX2_X1 U743 ( .A(DP_coeffs_ff_int[90]), .B(coeffs_ff[5]), .S(n1159), .Z(
        n1405) );
  MUX2_X1 U744 ( .A(DP_coeffs_ff_int[91]), .B(coeffs_ff[4]), .S(n1159), .Z(
        n1404) );
  MUX2_X1 U745 ( .A(DP_coeffs_ff_int[92]), .B(coeffs_ff[3]), .S(n1159), .Z(
        n1403) );
  MUX2_X1 U746 ( .A(DP_coeffs_ff_int[93]), .B(coeffs_ff[2]), .S(n1159), .Z(
        n1402) );
  MUX2_X1 U747 ( .A(DP_coeffs_ff_int[94]), .B(coeffs_ff[1]), .S(n1159), .Z(
        n1401) );
  MUX2_X1 U748 ( .A(DP_coeffs_ff_int[95]), .B(coeffs_ff[0]), .S(n1159), .Z(
        n1400) );
  MUX2_X1 U749 ( .A(DP_coeffs_ff_int[48]), .B(coeffs_ff[47]), .S(n1159), .Z(
        n1399) );
  MUX2_X1 U750 ( .A(DP_coeffs_ff_int[49]), .B(coeffs_ff[46]), .S(n1160), .Z(
        n1398) );
  MUX2_X1 U751 ( .A(DP_coeffs_ff_int[50]), .B(coeffs_ff[45]), .S(n1160), .Z(
        n1397) );
  MUX2_X1 U752 ( .A(DP_coeffs_ff_int[51]), .B(coeffs_ff[44]), .S(n1160), .Z(
        n1396) );
  MUX2_X1 U753 ( .A(DP_coeffs_ff_int[52]), .B(coeffs_ff[43]), .S(n1160), .Z(
        n1395) );
  MUX2_X1 U754 ( .A(DP_coeffs_ff_int[53]), .B(coeffs_ff[42]), .S(n1160), .Z(
        n1394) );
  MUX2_X1 U755 ( .A(DP_coeffs_ff_int[54]), .B(coeffs_ff[41]), .S(n1160), .Z(
        n1393) );
  MUX2_X1 U756 ( .A(DP_coeffs_ff_int[55]), .B(coeffs_ff[40]), .S(n1160), .Z(
        n1392) );
  MUX2_X1 U757 ( .A(DP_coeffs_ff_int[56]), .B(coeffs_ff[39]), .S(n1160), .Z(
        n1391) );
  MUX2_X1 U758 ( .A(DP_coeffs_ff_int[57]), .B(coeffs_ff[38]), .S(n1160), .Z(
        n1390) );
  MUX2_X1 U759 ( .A(DP_coeffs_ff_int[58]), .B(coeffs_ff[37]), .S(n1160), .Z(
        n1389) );
  MUX2_X1 U760 ( .A(DP_coeffs_ff_int[59]), .B(coeffs_ff[36]), .S(n1160), .Z(
        n1388) );
  MUX2_X1 U761 ( .A(DP_coeffs_ff_int[60]), .B(coeffs_ff[35]), .S(n1160), .Z(
        n1387) );
  MUX2_X1 U762 ( .A(DP_coeffs_ff_int[61]), .B(coeffs_ff[34]), .S(n1160), .Z(
        n1386) );
  MUX2_X1 U763 ( .A(DP_coeffs_ff_int[62]), .B(coeffs_ff[33]), .S(n1161), .Z(
        n1385) );
  MUX2_X1 U764 ( .A(DP_coeffs_ff_int[63]), .B(coeffs_ff[32]), .S(n1161), .Z(
        n1384) );
  MUX2_X1 U765 ( .A(DP_coeffs_ff_int[64]), .B(coeffs_ff[31]), .S(n1161), .Z(
        n1383) );
  MUX2_X1 U766 ( .A(DP_coeffs_ff_int[65]), .B(coeffs_ff[30]), .S(n1161), .Z(
        n1382) );
  MUX2_X1 U767 ( .A(DP_coeffs_ff_int[66]), .B(coeffs_ff[29]), .S(n1161), .Z(
        n1381) );
  MUX2_X1 U768 ( .A(DP_coeffs_ff_int[67]), .B(coeffs_ff[28]), .S(n1161), .Z(
        n1380) );
  MUX2_X1 U769 ( .A(DP_coeffs_ff_int[68]), .B(coeffs_ff[27]), .S(n1161), .Z(
        n1379) );
  MUX2_X1 U770 ( .A(DP_coeffs_ff_int[69]), .B(coeffs_ff[26]), .S(n1161), .Z(
        n1378) );
  MUX2_X1 U771 ( .A(DP_coeffs_ff_int[70]), .B(coeffs_ff[25]), .S(n1161), .Z(
        n1377) );
  MUX2_X1 U772 ( .A(DP_coeffs_ff_int[71]), .B(coeffs_ff[24]), .S(n1161), .Z(
        n1376) );
  MUX2_X1 U773 ( .A(DP_coeffs_ff_int[24]), .B(coeffs_ff[71]), .S(n1161), .Z(
        n1375) );
  MUX2_X1 U774 ( .A(DP_coeffs_ff_int[25]), .B(coeffs_ff[70]), .S(n1161), .Z(
        n1374) );
  MUX2_X1 U775 ( .A(DP_coeffs_ff_int[26]), .B(coeffs_ff[69]), .S(n1161), .Z(
        n1373) );
  MUX2_X1 U776 ( .A(DP_coeffs_ff_int[27]), .B(coeffs_ff[68]), .S(n1162), .Z(
        n1372) );
  MUX2_X1 U777 ( .A(DP_coeffs_ff_int[28]), .B(coeffs_ff[67]), .S(n1162), .Z(
        n1371) );
  MUX2_X1 U778 ( .A(DP_coeffs_ff_int[29]), .B(coeffs_ff[66]), .S(n1162), .Z(
        n1370) );
  MUX2_X1 U779 ( .A(DP_coeffs_ff_int[30]), .B(coeffs_ff[65]), .S(n1162), .Z(
        n1369) );
  MUX2_X1 U780 ( .A(DP_coeffs_ff_int[31]), .B(coeffs_ff[64]), .S(n1162), .Z(
        n1368) );
  MUX2_X1 U781 ( .A(DP_coeffs_ff_int[32]), .B(coeffs_ff[63]), .S(n1162), .Z(
        n1367) );
  MUX2_X1 U782 ( .A(DP_coeffs_ff_int[33]), .B(coeffs_ff[62]), .S(n1162), .Z(
        n1366) );
  MUX2_X1 U783 ( .A(DP_coeffs_ff_int[34]), .B(coeffs_ff[61]), .S(n1162), .Z(
        n1365) );
  MUX2_X1 U784 ( .A(DP_coeffs_ff_int[35]), .B(coeffs_ff[60]), .S(n1162), .Z(
        n1364) );
  MUX2_X1 U785 ( .A(DP_coeffs_ff_int[36]), .B(coeffs_ff[59]), .S(n1162), .Z(
        n1363) );
  MUX2_X1 U786 ( .A(DP_coeffs_ff_int[37]), .B(coeffs_ff[58]), .S(n1162), .Z(
        n1362) );
  MUX2_X1 U787 ( .A(DP_coeffs_ff_int[38]), .B(coeffs_ff[57]), .S(n1162), .Z(
        n1361) );
  MUX2_X1 U788 ( .A(DP_coeffs_ff_int[39]), .B(coeffs_ff[56]), .S(n1162), .Z(
        n1360) );
  MUX2_X1 U789 ( .A(DP_coeffs_ff_int[40]), .B(coeffs_ff[55]), .S(n1163), .Z(
        n1359) );
  MUX2_X1 U790 ( .A(DP_coeffs_ff_int[41]), .B(coeffs_ff[54]), .S(n1163), .Z(
        n1358) );
  MUX2_X1 U791 ( .A(DP_coeffs_ff_int[42]), .B(coeffs_ff[53]), .S(n1163), .Z(
        n1357) );
  MUX2_X1 U792 ( .A(DP_coeffs_ff_int[43]), .B(coeffs_ff[52]), .S(n1163), .Z(
        n1356) );
  MUX2_X1 U793 ( .A(DP_coeffs_ff_int[44]), .B(coeffs_ff[51]), .S(n1163), .Z(
        n1355) );
  MUX2_X1 U794 ( .A(DP_coeffs_ff_int[45]), .B(coeffs_ff[50]), .S(n1163), .Z(
        n1354) );
  MUX2_X1 U795 ( .A(DP_coeffs_ff_int[46]), .B(coeffs_ff[49]), .S(n1163), .Z(
        n1353) );
  MUX2_X1 U796 ( .A(DP_coeffs_ff_int[47]), .B(coeffs_ff[48]), .S(n1163), .Z(
        n1352) );
  MUX2_X1 U797 ( .A(DP_coeffs_ff_int[0]), .B(coeffs_ff[95]), .S(n1163), .Z(
        n1351) );
  MUX2_X1 U798 ( .A(DP_coeffs_ff_int[1]), .B(coeffs_ff[94]), .S(n1163), .Z(
        n1350) );
  MUX2_X1 U799 ( .A(DP_coeffs_ff_int[2]), .B(coeffs_ff[93]), .S(n1163), .Z(
        n1349) );
  MUX2_X1 U800 ( .A(DP_coeffs_ff_int[3]), .B(coeffs_ff[92]), .S(n1163), .Z(
        n1348) );
  MUX2_X1 U801 ( .A(DP_coeffs_ff_int[4]), .B(coeffs_ff[91]), .S(n1163), .Z(
        n1347) );
  MUX2_X1 U802 ( .A(DP_coeffs_ff_int[5]), .B(coeffs_ff[90]), .S(n1164), .Z(
        n1346) );
  MUX2_X1 U803 ( .A(DP_coeffs_ff_int[6]), .B(coeffs_ff[89]), .S(n1164), .Z(
        n1345) );
  MUX2_X1 U804 ( .A(DP_coeffs_ff_int[7]), .B(coeffs_ff[88]), .S(n1164), .Z(
        n1344) );
  MUX2_X1 U805 ( .A(DP_coeffs_ff_int[8]), .B(coeffs_ff[87]), .S(n1164), .Z(
        n1343) );
  MUX2_X1 U806 ( .A(DP_coeffs_ff_int[9]), .B(coeffs_ff[86]), .S(n1164), .Z(
        n1342) );
  MUX2_X1 U807 ( .A(DP_coeffs_ff_int[10]), .B(coeffs_ff[85]), .S(n1164), .Z(
        n1341) );
  MUX2_X1 U808 ( .A(DP_coeffs_ff_int[11]), .B(coeffs_ff[84]), .S(n1164), .Z(
        n1340) );
  MUX2_X1 U809 ( .A(DP_coeffs_ff_int[12]), .B(coeffs_ff[83]), .S(n1164), .Z(
        n1339) );
  MUX2_X1 U810 ( .A(DP_coeffs_ff_int[13]), .B(coeffs_ff[82]), .S(n1164), .Z(
        n1338) );
  MUX2_X1 U811 ( .A(DP_coeffs_ff_int[14]), .B(coeffs_ff[81]), .S(n1164), .Z(
        n1337) );
  MUX2_X1 U812 ( .A(DP_coeffs_ff_int[15]), .B(coeffs_ff[80]), .S(n1164), .Z(
        n1336) );
  MUX2_X1 U813 ( .A(DP_coeffs_ff_int[16]), .B(coeffs_ff[79]), .S(n1164), .Z(
        n1335) );
  MUX2_X1 U814 ( .A(DP_coeffs_ff_int[17]), .B(coeffs_ff[78]), .S(n1164), .Z(
        n1334) );
  MUX2_X1 U815 ( .A(DP_coeffs_ff_int[18]), .B(coeffs_ff[77]), .S(n1165), .Z(
        n1333) );
  MUX2_X1 U816 ( .A(DP_coeffs_ff_int[19]), .B(coeffs_ff[76]), .S(n1165), .Z(
        n1332) );
  MUX2_X1 U817 ( .A(DP_coeffs_ff_int[20]), .B(coeffs_ff[75]), .S(n1165), .Z(
        n1331) );
  MUX2_X1 U818 ( .A(DP_coeffs_ff_int[21]), .B(coeffs_ff[74]), .S(n1165), .Z(
        n1330) );
  MUX2_X1 U819 ( .A(DP_coeffs_ff_int[22]), .B(coeffs_ff[73]), .S(n1165), .Z(
        n1329) );
  MUX2_X1 U820 ( .A(DP_coeffs_ff_int[23]), .B(coeffs_ff[72]), .S(n1165), .Z(
        n1328) );
  MUX2_X1 U821 ( .A(DP_coeffs_fb_int[24]), .B(coeffs_fb[23]), .S(n1165), .Z(
        n1327) );
  MUX2_X1 U822 ( .A(DP_coeffs_fb_int[25]), .B(coeffs_fb[22]), .S(n1165), .Z(
        n1326) );
  MUX2_X1 U823 ( .A(DP_coeffs_fb_int[26]), .B(coeffs_fb[21]), .S(n1165), .Z(
        n1325) );
  MUX2_X1 U824 ( .A(DP_coeffs_fb_int[27]), .B(coeffs_fb[20]), .S(n1165), .Z(
        n1324) );
  MUX2_X1 U825 ( .A(DP_coeffs_fb_int[28]), .B(coeffs_fb[19]), .S(n1165), .Z(
        n1323) );
  MUX2_X1 U826 ( .A(DP_coeffs_fb_int[29]), .B(coeffs_fb[18]), .S(n1165), .Z(
        n1322) );
  MUX2_X1 U827 ( .A(DP_coeffs_fb_int[30]), .B(coeffs_fb[17]), .S(n1165), .Z(
        n1321) );
  MUX2_X1 U828 ( .A(DP_coeffs_fb_int[31]), .B(coeffs_fb[16]), .S(n1166), .Z(
        n1320) );
  MUX2_X1 U829 ( .A(DP_coeffs_fb_int[32]), .B(coeffs_fb[15]), .S(n1166), .Z(
        n1319) );
  MUX2_X1 U830 ( .A(DP_coeffs_fb_int[33]), .B(coeffs_fb[14]), .S(n1166), .Z(
        n1318) );
  MUX2_X1 U831 ( .A(DP_coeffs_fb_int[34]), .B(coeffs_fb[13]), .S(n1166), .Z(
        n1317) );
  MUX2_X1 U832 ( .A(DP_coeffs_fb_int[35]), .B(coeffs_fb[12]), .S(n1166), .Z(
        n1316) );
  MUX2_X1 U833 ( .A(DP_coeffs_fb_int[36]), .B(coeffs_fb[11]), .S(n1166), .Z(
        n1315) );
  MUX2_X1 U834 ( .A(DP_coeffs_fb_int[37]), .B(coeffs_fb[10]), .S(n1166), .Z(
        n1314) );
  MUX2_X1 U835 ( .A(DP_coeffs_fb_int[38]), .B(coeffs_fb[9]), .S(n1166), .Z(
        n1313) );
  MUX2_X1 U836 ( .A(DP_coeffs_fb_int[39]), .B(coeffs_fb[8]), .S(n1166), .Z(
        n1312) );
  MUX2_X1 U837 ( .A(DP_coeffs_fb_int[40]), .B(coeffs_fb[7]), .S(n1166), .Z(
        n1311) );
  MUX2_X1 U838 ( .A(DP_coeffs_fb_int[41]), .B(coeffs_fb[6]), .S(n1166), .Z(
        n1310) );
  MUX2_X1 U839 ( .A(DP_coeffs_fb_int[42]), .B(coeffs_fb[5]), .S(n1166), .Z(
        n1309) );
  MUX2_X1 U840 ( .A(DP_coeffs_fb_int[43]), .B(coeffs_fb[4]), .S(n1166), .Z(
        n1308) );
  MUX2_X1 U841 ( .A(n1038), .B(coeffs_fb[3]), .S(n1167), .Z(n1307) );
  MUX2_X1 U842 ( .A(DP_coeffs_fb_int[45]), .B(coeffs_fb[2]), .S(n1167), .Z(
        n1306) );
  MUX2_X1 U843 ( .A(DP_coeffs_fb_int[46]), .B(coeffs_fb[1]), .S(n1167), .Z(
        n1305) );
  MUX2_X1 U844 ( .A(DP_coeffs_fb_int[47]), .B(coeffs_fb[0]), .S(n1167), .Z(
        n1304) );
  MUX2_X1 U845 ( .A(DP_coeffs_fb_int[0]), .B(coeffs_fb[47]), .S(n1167), .Z(
        n1303) );
  MUX2_X1 U846 ( .A(DP_coeffs_fb_int[1]), .B(coeffs_fb[46]), .S(n1167), .Z(
        n1302) );
  MUX2_X1 U847 ( .A(DP_coeffs_fb_int[2]), .B(coeffs_fb[45]), .S(n1167), .Z(
        n1301) );
  MUX2_X1 U848 ( .A(DP_coeffs_fb_int[3]), .B(coeffs_fb[44]), .S(n1167), .Z(
        n1300) );
  MUX2_X1 U849 ( .A(DP_coeffs_fb_int[4]), .B(coeffs_fb[43]), .S(n1167), .Z(
        n1299) );
  MUX2_X1 U850 ( .A(DP_coeffs_fb_int[5]), .B(coeffs_fb[42]), .S(n1167), .Z(
        n1298) );
  MUX2_X1 U851 ( .A(DP_coeffs_fb_int[6]), .B(coeffs_fb[41]), .S(n1167), .Z(
        n1297) );
  MUX2_X1 U852 ( .A(DP_coeffs_fb_int[7]), .B(coeffs_fb[40]), .S(n1167), .Z(
        n1296) );
  MUX2_X1 U853 ( .A(DP_coeffs_fb_int[8]), .B(coeffs_fb[39]), .S(n1167), .Z(
        n1295) );
  MUX2_X1 U854 ( .A(DP_coeffs_fb_int[9]), .B(coeffs_fb[38]), .S(n1168), .Z(
        n1294) );
  MUX2_X1 U855 ( .A(DP_coeffs_fb_int[10]), .B(coeffs_fb[37]), .S(n1168), .Z(
        n1293) );
  MUX2_X1 U856 ( .A(DP_coeffs_fb_int[11]), .B(coeffs_fb[36]), .S(n1168), .Z(
        n1292) );
  MUX2_X1 U857 ( .A(DP_coeffs_fb_int[12]), .B(coeffs_fb[35]), .S(n1168), .Z(
        n1291) );
  MUX2_X1 U858 ( .A(DP_coeffs_fb_int[13]), .B(coeffs_fb[34]), .S(n1168), .Z(
        n1290) );
  MUX2_X1 U859 ( .A(DP_coeffs_fb_int[14]), .B(coeffs_fb[33]), .S(n1168), .Z(
        n1289) );
  MUX2_X1 U860 ( .A(DP_coeffs_fb_int[15]), .B(coeffs_fb[32]), .S(n1168), .Z(
        n1288) );
  MUX2_X1 U861 ( .A(DP_coeffs_fb_int[16]), .B(coeffs_fb[31]), .S(n1168), .Z(
        n1287) );
  MUX2_X1 U862 ( .A(DP_coeffs_fb_int[17]), .B(coeffs_fb[30]), .S(n1168), .Z(
        n1286) );
  MUX2_X1 U863 ( .A(DP_coeffs_fb_int[18]), .B(coeffs_fb[29]), .S(n1168), .Z(
        n1285) );
  MUX2_X1 U864 ( .A(DP_coeffs_fb_int[19]), .B(coeffs_fb[28]), .S(n1168), .Z(
        n1284) );
  MUX2_X1 U865 ( .A(DP_coeffs_fb_int[20]), .B(coeffs_fb[27]), .S(n1168), .Z(
        n1283) );
  MUX2_X1 U866 ( .A(DP_coeffs_fb_int[21]), .B(coeffs_fb[26]), .S(n1168), .Z(
        n1282) );
  MUX2_X1 U867 ( .A(DP_coeffs_fb_int[22]), .B(coeffs_fb[25]), .S(n1169), .Z(
        n1281) );
  MUX2_X1 U868 ( .A(DP_coeffs_fb_int[23]), .B(coeffs_fb[24]), .S(n1169), .Z(
        n1280) );
  MUX2_X1 U869 ( .A(DP_x[11]), .B(dIn[11]), .S(n1169), .Z(n1279) );
  MUX2_X1 U870 ( .A(DP_x[10]), .B(dIn[10]), .S(n1169), .Z(n1278) );
  MUX2_X1 U871 ( .A(DP_x[9]), .B(dIn[9]), .S(n1169), .Z(n1277) );
  MUX2_X1 U872 ( .A(DP_x[8]), .B(dIn[8]), .S(n1169), .Z(n1276) );
  MUX2_X1 U873 ( .A(DP_x[7]), .B(dIn[7]), .S(n1169), .Z(n1275) );
  MUX2_X1 U874 ( .A(DP_x[6]), .B(dIn[6]), .S(n1169), .Z(n1274) );
  MUX2_X1 U875 ( .A(DP_x[5]), .B(dIn[5]), .S(n1169), .Z(n1273) );
  MUX2_X1 U876 ( .A(DP_x[4]), .B(dIn[4]), .S(n1169), .Z(n1272) );
  MUX2_X1 U877 ( .A(DP_x[3]), .B(dIn[3]), .S(n1169), .Z(n1271) );
  MUX2_X1 U878 ( .A(DP_x[2]), .B(dIn[2]), .S(n1169), .Z(n1270) );
  MUX2_X1 U879 ( .A(DP_x[1]), .B(dIn[1]), .S(n1169), .Z(n1269) );
endmodule

