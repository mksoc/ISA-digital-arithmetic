
module iir_filter_DW02_mult_5 ( A, B, PRODUCT, TC );
  input [23:0] A;
  input [23:0] B;
  output [47:0] PRODUCT;
  input TC;
  wire   n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n351, n352, n353, n354, n355, n356, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n906, n907, n908, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134;

  FA_X1 U182 ( .A(n351), .B(n352), .CI(n304), .CO(n303), .S(PRODUCT[44]) );
  FA_X1 U183 ( .A(n353), .B(n354), .CI(n305), .CO(n304), .S(PRODUCT[43]) );
  FA_X1 U184 ( .A(n355), .B(n358), .CI(n306), .CO(n305), .S(PRODUCT[42]) );
  FA_X1 U185 ( .A(n359), .B(n361), .CI(n307), .CO(n306), .S(PRODUCT[41]) );
  FA_X1 U186 ( .A(n362), .B(n364), .CI(n308), .CO(n307), .S(PRODUCT[40]) );
  FA_X1 U187 ( .A(n365), .B(n370), .CI(n309), .CO(n308), .S(PRODUCT[39]) );
  FA_X1 U188 ( .A(n371), .B(n375), .CI(n310), .CO(n309), .S(PRODUCT[38]) );
  FA_X1 U189 ( .A(n376), .B(n381), .CI(n311), .CO(n310), .S(PRODUCT[37]) );
  FA_X1 U190 ( .A(n382), .B(n389), .CI(n312), .CO(n311), .S(PRODUCT[36]) );
  FA_X1 U191 ( .A(n390), .B(n396), .CI(n313), .CO(n312), .S(PRODUCT[35]) );
  FA_X1 U192 ( .A(n397), .B(n403), .CI(n314), .CO(n313), .S(PRODUCT[34]) );
  FA_X1 U193 ( .A(n404), .B(n413), .CI(n315), .CO(n314), .S(PRODUCT[33]) );
  FA_X1 U194 ( .A(n414), .B(n422), .CI(n316), .CO(n315), .S(PRODUCT[32]) );
  FA_X1 U195 ( .A(n423), .B(n432), .CI(n317), .CO(n316), .S(PRODUCT[31]) );
  FA_X1 U196 ( .A(n433), .B(n444), .CI(n318), .CO(n317), .S(PRODUCT[30]) );
  FA_X1 U197 ( .A(n445), .B(n455), .CI(n319), .CO(n318), .S(PRODUCT[29]) );
  FA_X1 U198 ( .A(n456), .B(n467), .CI(n320), .CO(n319), .S(PRODUCT[28]) );
  FA_X1 U199 ( .A(n468), .B(n481), .CI(n321), .CO(n320), .S(PRODUCT[27]) );
  FA_X1 U200 ( .A(n482), .B(n494), .CI(n322), .CO(n321), .S(PRODUCT[26]) );
  FA_X1 U201 ( .A(n495), .B(n507), .CI(n323), .CO(n322), .S(PRODUCT[25]) );
  FA_X1 U202 ( .A(n508), .B(n906), .CI(n324), .CO(n323), .S(PRODUCT[24]) );
  FA_X1 U203 ( .A(n907), .B(n522), .CI(n325), .CO(n324), .S(PRODUCT[23]) );
  FA_X1 U204 ( .A(n908), .B(n536), .CI(n326), .CO(n325), .S(PRODUCT[22]) );
  FA_X1 U235 ( .A(n356), .B(n749), .CI(n729), .CO(n352), .S(n353) );
  FA_X1 U236 ( .A(n730), .B(n360), .CI(n750), .CO(n354), .S(n355) );
  FA_X1 U238 ( .A(n360), .B(n731), .CI(n751), .CO(n358), .S(n359) );
  FA_X1 U240 ( .A(n752), .B(n363), .CI(n366), .CO(n361), .S(n362) );
  FA_X1 U241 ( .A(n368), .B(n775), .CI(n732), .CO(n356), .S(n363) );
  FA_X1 U242 ( .A(n776), .B(n753), .CI(n367), .CO(n364), .S(n365) );
  FA_X1 U243 ( .A(n733), .B(n374), .CI(n372), .CO(n366), .S(n367) );
  FA_X1 U245 ( .A(n373), .B(n377), .CI(n777), .CO(n370), .S(n371) );
  FA_X1 U246 ( .A(n374), .B(n379), .CI(n754), .CO(n372), .S(n373) );
  FA_X1 U248 ( .A(n778), .B(n378), .CI(n383), .CO(n375), .S(n376) );
  FA_X1 U249 ( .A(n385), .B(n380), .CI(n755), .CO(n377), .S(n378) );
  FA_X1 U250 ( .A(n387), .B(n801), .CI(n734), .CO(n379), .S(n380) );
  FA_X1 U251 ( .A(n802), .B(n779), .CI(n384), .CO(n381), .S(n382) );
  FA_X1 U252 ( .A(n386), .B(n393), .CI(n391), .CO(n383), .S(n384) );
  FA_X1 U253 ( .A(n735), .B(n395), .CI(n756), .CO(n385), .S(n386) );
  FA_X1 U255 ( .A(n392), .B(n398), .CI(n803), .CO(n389), .S(n390) );
  FA_X1 U256 ( .A(n394), .B(n400), .CI(n780), .CO(n391), .S(n392) );
  FA_X1 U257 ( .A(n395), .B(n736), .CI(n757), .CO(n393), .S(n394) );
  FA_X1 U259 ( .A(n804), .B(n399), .CI(n405), .CO(n396), .S(n397) );
  FA_X1 U260 ( .A(n407), .B(n401), .CI(n781), .CO(n398), .S(n399) );
  FA_X1 U261 ( .A(n758), .B(n402), .CI(n409), .CO(n400), .S(n401) );
  FA_X1 U262 ( .A(n411), .B(n827), .CI(n737), .CO(n387), .S(n402) );
  FA_X1 U263 ( .A(n828), .B(n805), .CI(n406), .CO(n403), .S(n404) );
  FA_X1 U264 ( .A(n408), .B(n417), .CI(n415), .CO(n405), .S(n406) );
  FA_X1 U265 ( .A(n410), .B(n759), .CI(n782), .CO(n407), .S(n408) );
  FA_X1 U266 ( .A(n738), .B(n421), .CI(n419), .CO(n409), .S(n410) );
  FA_X1 U268 ( .A(n416), .B(n424), .CI(n829), .CO(n413), .S(n414) );
  FA_X1 U269 ( .A(n418), .B(n426), .CI(n806), .CO(n415), .S(n416) );
  FA_X1 U270 ( .A(n420), .B(n428), .CI(n783), .CO(n417), .S(n418) );
  FA_X1 U271 ( .A(n421), .B(n430), .CI(n760), .CO(n419), .S(n420) );
  FA_X1 U273 ( .A(n830), .B(n425), .CI(n434), .CO(n422), .S(n423) );
  FA_X1 U274 ( .A(n436), .B(n427), .CI(n807), .CO(n424), .S(n425) );
  FA_X1 U275 ( .A(n784), .B(n429), .CI(n438), .CO(n426), .S(n427) );
  FA_X1 U276 ( .A(n440), .B(n431), .CI(n761), .CO(n428), .S(n429) );
  FA_X1 U277 ( .A(n442), .B(n853), .CI(n739), .CO(n430), .S(n431) );
  FA_X1 U278 ( .A(n854), .B(n831), .CI(n435), .CO(n432), .S(n433) );
  FA_X1 U279 ( .A(n437), .B(n448), .CI(n446), .CO(n434), .S(n435) );
  FA_X1 U280 ( .A(n439), .B(n785), .CI(n808), .CO(n436), .S(n437) );
  FA_X1 U281 ( .A(n441), .B(n452), .CI(n450), .CO(n438), .S(n439) );
  FA_X1 U282 ( .A(n740), .B(n454), .CI(n762), .CO(n440), .S(n441) );
  FA_X1 U284 ( .A(n447), .B(n457), .CI(n855), .CO(n444), .S(n445) );
  FA_X1 U285 ( .A(n449), .B(n459), .CI(n832), .CO(n446), .S(n447) );
  FA_X1 U286 ( .A(n451), .B(n461), .CI(n809), .CO(n448), .S(n449) );
  FA_X1 U287 ( .A(n453), .B(n463), .CI(n786), .CO(n450), .S(n451) );
  FA_X1 U288 ( .A(n454), .B(n465), .CI(n763), .CO(n452), .S(n453) );
  FA_X1 U290 ( .A(n856), .B(n458), .CI(n469), .CO(n455), .S(n456) );
  FA_X1 U291 ( .A(n471), .B(n460), .CI(n833), .CO(n457), .S(n458) );
  FA_X1 U292 ( .A(n810), .B(n462), .CI(n473), .CO(n459), .S(n460) );
  FA_X1 U293 ( .A(n475), .B(n464), .CI(n787), .CO(n461), .S(n462) );
  FA_X1 U294 ( .A(n764), .B(n466), .CI(n477), .CO(n463), .S(n464) );
  FA_X1 U295 ( .A(n479), .B(n879), .CI(n741), .CO(n465), .S(n466) );
  FA_X1 U296 ( .A(n880), .B(n857), .CI(n470), .CO(n467), .S(n468) );
  FA_X1 U297 ( .A(n472), .B(n485), .CI(n483), .CO(n469), .S(n470) );
  FA_X1 U298 ( .A(n474), .B(n811), .CI(n834), .CO(n471), .S(n472) );
  FA_X1 U299 ( .A(n476), .B(n489), .CI(n487), .CO(n473), .S(n474) );
  FA_X1 U300 ( .A(n478), .B(n765), .CI(n788), .CO(n475), .S(n476) );
  FA_X1 U301 ( .A(n742), .B(n493), .CI(n491), .CO(n477), .S(n478) );
  FA_X1 U303 ( .A(n484), .B(n858), .CI(n881), .CO(n481), .S(n482) );
  FA_X1 U304 ( .A(n486), .B(n498), .CI(n496), .CO(n483), .S(n484) );
  FA_X1 U305 ( .A(n488), .B(n812), .CI(n835), .CO(n485), .S(n486) );
  FA_X1 U306 ( .A(n490), .B(n502), .CI(n500), .CO(n487), .S(n488) );
  FA_X1 U307 ( .A(n492), .B(n504), .CI(n789), .CO(n489), .S(n490) );
  FA_X1 U308 ( .A(n743), .B(n493), .CI(n766), .CO(n491), .S(n492) );
  FA_X1 U310 ( .A(n497), .B(n509), .CI(n882), .CO(n494), .S(n495) );
  FA_X1 U311 ( .A(n499), .B(n511), .CI(n859), .CO(n496), .S(n497) );
  FA_X1 U312 ( .A(n501), .B(n513), .CI(n836), .CO(n498), .S(n499) );
  FA_X1 U313 ( .A(n503), .B(n515), .CI(n813), .CO(n500), .S(n501) );
  FA_X1 U314 ( .A(n505), .B(n517), .CI(n790), .CO(n502), .S(n503) );
  FA_X1 U315 ( .A(n506), .B(n744), .CI(n767), .CO(n504), .S(n505) );
  FA_X1 U318 ( .A(n883), .B(n510), .CI(n521), .CO(n507), .S(n508) );
  FA_X1 U319 ( .A(n860), .B(n512), .CI(n523), .CO(n509), .S(n510) );
  FA_X1 U320 ( .A(n837), .B(n514), .CI(n525), .CO(n511), .S(n512) );
  FA_X1 U321 ( .A(n814), .B(n516), .CI(n527), .CO(n513), .S(n514) );
  FA_X1 U322 ( .A(n791), .B(n518), .CI(n529), .CO(n515), .S(n516) );
  FA_X1 U323 ( .A(n768), .B(n520), .CI(n531), .CO(n517), .S(n518) );
  HA_X1 U324 ( .A(n533), .B(n745), .CO(n519), .S(n520) );
  FA_X1 U325 ( .A(n884), .B(n524), .CI(n535), .CO(n521), .S(n522) );
  FA_X1 U326 ( .A(n861), .B(n526), .CI(n537), .CO(n523), .S(n524) );
  FA_X1 U327 ( .A(n838), .B(n528), .CI(n539), .CO(n525), .S(n526) );
  FA_X1 U328 ( .A(n815), .B(n530), .CI(n541), .CO(n527), .S(n528) );
  FA_X1 U329 ( .A(n792), .B(n532), .CI(n543), .CO(n529), .S(n530) );
  FA_X1 U330 ( .A(n769), .B(n534), .CI(n545), .CO(n531), .S(n532) );
  HA_X1 U331 ( .A(n547), .B(n746), .CO(n533), .S(n534) );
  FA_X1 U332 ( .A(n885), .B(n538), .CI(n549), .CO(n535), .S(n536) );
  FA_X1 U333 ( .A(n862), .B(n540), .CI(n551), .CO(n537), .S(n538) );
  FA_X1 U334 ( .A(n839), .B(n542), .CI(n553), .CO(n539), .S(n540) );
  FA_X1 U335 ( .A(n816), .B(n544), .CI(n555), .CO(n541), .S(n542) );
  FA_X1 U336 ( .A(n793), .B(n546), .CI(n557), .CO(n543), .S(n544) );
  FA_X1 U337 ( .A(n770), .B(n548), .CI(n559), .CO(n545), .S(n546) );
  HA_X1 U338 ( .A(n561), .B(n747), .CO(n547), .S(n548) );
  FA_X1 U339 ( .A(n886), .B(n552), .CI(n563), .CO(n549), .S(n550) );
  FA_X1 U340 ( .A(n863), .B(n554), .CI(n565), .CO(n551), .S(n552) );
  FA_X1 U341 ( .A(n840), .B(n556), .CI(n567), .CO(n553), .S(n554) );
  FA_X1 U342 ( .A(n817), .B(n558), .CI(n569), .CO(n555), .S(n556) );
  FA_X1 U343 ( .A(n794), .B(n560), .CI(n571), .CO(n557), .S(n558) );
  FA_X1 U344 ( .A(n771), .B(n562), .CI(n573), .CO(n559), .S(n560) );
  HA_X1 U345 ( .A(n748), .B(n1540), .CO(n561), .S(n562) );
  FA_X1 U346 ( .A(n887), .B(n566), .CI(n575), .CO(n563), .S(n564) );
  FA_X1 U347 ( .A(n864), .B(n568), .CI(n577), .CO(n565), .S(n566) );
  FA_X1 U348 ( .A(n841), .B(n570), .CI(n579), .CO(n567), .S(n568) );
  FA_X1 U349 ( .A(n818), .B(n572), .CI(n581), .CO(n569), .S(n570) );
  FA_X1 U350 ( .A(n795), .B(n574), .CI(n583), .CO(n571), .S(n572) );
  HA_X1 U351 ( .A(n585), .B(n772), .CO(n573), .S(n574) );
  FA_X1 U352 ( .A(n888), .B(n578), .CI(n587), .CO(n575), .S(n576) );
  FA_X1 U353 ( .A(n865), .B(n580), .CI(n589), .CO(n577), .S(n578) );
  FA_X1 U354 ( .A(n842), .B(n582), .CI(n591), .CO(n579), .S(n580) );
  FA_X1 U355 ( .A(n819), .B(n584), .CI(n593), .CO(n581), .S(n582) );
  FA_X1 U356 ( .A(n796), .B(n586), .CI(n595), .CO(n583), .S(n584) );
  HA_X1 U357 ( .A(n597), .B(n773), .CO(n585), .S(n586) );
  FA_X1 U358 ( .A(n889), .B(n590), .CI(n599), .CO(n587), .S(n588) );
  FA_X1 U359 ( .A(n866), .B(n592), .CI(n601), .CO(n589), .S(n590) );
  FA_X1 U360 ( .A(n843), .B(n594), .CI(n603), .CO(n591), .S(n592) );
  FA_X1 U361 ( .A(n820), .B(n596), .CI(n605), .CO(n593), .S(n594) );
  FA_X1 U362 ( .A(n797), .B(n598), .CI(n607), .CO(n595), .S(n596) );
  HA_X1 U363 ( .A(n774), .B(n1542), .CO(n597), .S(n598) );
  FA_X1 U364 ( .A(n890), .B(n602), .CI(n609), .CO(n599), .S(n600) );
  FA_X1 U365 ( .A(n867), .B(n604), .CI(n611), .CO(n601), .S(n602) );
  FA_X1 U366 ( .A(n844), .B(n606), .CI(n613), .CO(n603), .S(n604) );
  FA_X1 U367 ( .A(n821), .B(n608), .CI(n615), .CO(n605), .S(n606) );
  HA_X1 U368 ( .A(n617), .B(n798), .CO(n607), .S(n608) );
  FA_X1 U369 ( .A(n891), .B(n612), .CI(n619), .CO(n609), .S(n610) );
  FA_X1 U370 ( .A(n868), .B(n614), .CI(n621), .CO(n611), .S(n612) );
  FA_X1 U371 ( .A(n845), .B(n616), .CI(n623), .CO(n613), .S(n614) );
  FA_X1 U372 ( .A(n822), .B(n618), .CI(n625), .CO(n615), .S(n616) );
  HA_X1 U373 ( .A(n627), .B(n799), .CO(n617), .S(n618) );
  FA_X1 U374 ( .A(n892), .B(n622), .CI(n629), .CO(n619), .S(n620) );
  FA_X1 U375 ( .A(n869), .B(n624), .CI(n631), .CO(n621), .S(n622) );
  FA_X1 U376 ( .A(n846), .B(n626), .CI(n633), .CO(n623), .S(n624) );
  FA_X1 U377 ( .A(n823), .B(n628), .CI(n635), .CO(n625), .S(n626) );
  HA_X1 U378 ( .A(n800), .B(n1544), .CO(n627), .S(n628) );
  FA_X1 U379 ( .A(n893), .B(n632), .CI(n637), .CO(n629), .S(n630) );
  FA_X1 U380 ( .A(n870), .B(n634), .CI(n639), .CO(n631), .S(n632) );
  FA_X1 U381 ( .A(n847), .B(n636), .CI(n641), .CO(n633), .S(n634) );
  HA_X1 U382 ( .A(n643), .B(n824), .CO(n635), .S(n636) );
  FA_X1 U383 ( .A(n894), .B(n640), .CI(n645), .CO(n637), .S(n638) );
  FA_X1 U384 ( .A(n871), .B(n642), .CI(n647), .CO(n639), .S(n640) );
  FA_X1 U385 ( .A(n848), .B(n644), .CI(n649), .CO(n641), .S(n642) );
  HA_X1 U386 ( .A(n651), .B(n825), .CO(n643), .S(n644) );
  FA_X1 U387 ( .A(n895), .B(n648), .CI(n653), .CO(n645), .S(n646) );
  FA_X1 U388 ( .A(n872), .B(n650), .CI(n655), .CO(n647), .S(n648) );
  FA_X1 U389 ( .A(n849), .B(n652), .CI(n657), .CO(n649), .S(n650) );
  HA_X1 U390 ( .A(n826), .B(n1546), .CO(n651), .S(n652) );
  FA_X1 U391 ( .A(n896), .B(n656), .CI(n659), .CO(n653), .S(n654) );
  FA_X1 U392 ( .A(n873), .B(n658), .CI(n661), .CO(n655), .S(n656) );
  HA_X1 U393 ( .A(n663), .B(n850), .CO(n657), .S(n658) );
  FA_X1 U394 ( .A(n897), .B(n662), .CI(n665), .CO(n659), .S(n660) );
  FA_X1 U395 ( .A(n874), .B(n664), .CI(n667), .CO(n661), .S(n662) );
  HA_X1 U396 ( .A(n669), .B(n851), .CO(n663), .S(n664) );
  FA_X1 U397 ( .A(n898), .B(n668), .CI(n671), .CO(n665), .S(n666) );
  FA_X1 U398 ( .A(n875), .B(n670), .CI(n673), .CO(n667), .S(n668) );
  HA_X1 U399 ( .A(n852), .B(n1548), .CO(n669), .S(n670) );
  FA_X1 U400 ( .A(n899), .B(n674), .CI(n675), .CO(n671), .S(n672) );
  HA_X1 U401 ( .A(n677), .B(n876), .CO(n673), .S(n674) );
  FA_X1 U402 ( .A(n900), .B(n678), .CI(n679), .CO(n675), .S(n676) );
  HA_X1 U403 ( .A(n681), .B(n877), .CO(n677), .S(n678) );
  FA_X1 U404 ( .A(n901), .B(n682), .CI(n683), .CO(n679), .S(n680) );
  HA_X1 U405 ( .A(n878), .B(n1550), .CO(n681), .S(n682) );
  HA_X1 U406 ( .A(n685), .B(n902), .CO(n683), .S(n684) );
  HA_X1 U407 ( .A(n687), .B(n903), .CO(n685), .S(n686) );
  HA_X1 U408 ( .A(n904), .B(n1552), .CO(n687), .S(n688) );
  FA_X1 U1112 ( .A(B[22]), .B(n1554), .CI(n706), .CO(n1374), .S(n1375) );
  FA_X1 U1113 ( .A(B[21]), .B(B[22]), .CI(n707), .CO(n706), .S(n1376) );
  FA_X1 U1114 ( .A(B[20]), .B(B[21]), .CI(n708), .CO(n707), .S(n1377) );
  FA_X1 U1115 ( .A(B[19]), .B(B[20]), .CI(n709), .CO(n708), .S(n1378) );
  FA_X1 U1116 ( .A(B[18]), .B(B[19]), .CI(n710), .CO(n709), .S(n1379) );
  FA_X1 U1117 ( .A(B[17]), .B(B[18]), .CI(n711), .CO(n710), .S(n1380) );
  FA_X1 U1118 ( .A(B[16]), .B(B[17]), .CI(n712), .CO(n711), .S(n1381) );
  FA_X1 U1119 ( .A(B[15]), .B(B[16]), .CI(n713), .CO(n712), .S(n1382) );
  FA_X1 U1120 ( .A(B[14]), .B(B[15]), .CI(n714), .CO(n713), .S(n1383) );
  FA_X1 U1121 ( .A(B[13]), .B(B[14]), .CI(n715), .CO(n714), .S(n1384) );
  FA_X1 U1122 ( .A(B[12]), .B(B[13]), .CI(n716), .CO(n715), .S(n1385) );
  FA_X1 U1123 ( .A(B[11]), .B(B[12]), .CI(n717), .CO(n716), .S(n1386) );
  FA_X1 U1124 ( .A(B[10]), .B(B[11]), .CI(n718), .CO(n717), .S(n1387) );
  FA_X1 U1125 ( .A(B[9]), .B(B[10]), .CI(n719), .CO(n718), .S(n1388) );
  FA_X1 U1126 ( .A(B[8]), .B(B[9]), .CI(n720), .CO(n719), .S(n1389) );
  FA_X1 U1127 ( .A(B[7]), .B(B[8]), .CI(n721), .CO(n720), .S(n1390) );
  FA_X1 U1128 ( .A(B[6]), .B(B[7]), .CI(n722), .CO(n721), .S(n1391) );
  FA_X1 U1129 ( .A(B[5]), .B(B[6]), .CI(n723), .CO(n722), .S(n1392) );
  FA_X1 U1130 ( .A(B[4]), .B(B[5]), .CI(n724), .CO(n723), .S(n1393) );
  FA_X1 U1131 ( .A(B[3]), .B(B[4]), .CI(n725), .CO(n724), .S(n1394) );
  FA_X1 U1132 ( .A(B[2]), .B(B[3]), .CI(n726), .CO(n725), .S(n1395) );
  FA_X1 U1133 ( .A(B[1]), .B(B[2]), .CI(n727), .CO(n726), .S(n1396) );
  HA_X1 U1134 ( .A(B[0]), .B(B[1]), .CO(n727), .S(n1397) );
  OR2_X1 U1138 ( .A1(n2134), .A2(n2133), .ZN(n1534) );
  INV_X1 U1139 ( .A(n1534), .ZN(n1536) );
  INV_X1 U1140 ( .A(n1535), .ZN(n1537) );
  BUF_X1 U1141 ( .A(n1980), .Z(n1538) );
  BUF_X1 U1142 ( .A(n1980), .Z(n1539) );
  NAND3_X1 U1143 ( .A1(n1673), .A2(n1672), .A3(n1671), .ZN(n1586) );
  NAND3_X1 U1144 ( .A1(n1854), .A2(n1853), .A3(n1852), .ZN(n1804) );
  NAND3_X1 U1145 ( .A1(n1794), .A2(n1793), .A3(n1792), .ZN(n1744) );
  NAND3_X1 U1146 ( .A1(n1734), .A2(n1733), .A3(n1732), .ZN(n1684) );
  NAND3_X1 U1147 ( .A1(n2111), .A2(n2112), .A3(n2113), .ZN(n1563) );
  NAND2_X1 U1148 ( .A1(n1911), .A2(n1913), .ZN(n1857) );
  NAND2_X1 U1149 ( .A1(n1851), .A2(n1853), .ZN(n1797) );
  NAND2_X1 U1150 ( .A1(n1791), .A2(n1793), .ZN(n1737) );
  NAND2_X1 U1151 ( .A1(n1731), .A2(n1733), .ZN(n1677) );
  INV_X1 U1152 ( .A(n1553), .ZN(n1552) );
  INV_X1 U1153 ( .A(n1549), .ZN(n1548) );
  INV_X1 U1154 ( .A(n1551), .ZN(n1550) );
  NAND3_X1 U1155 ( .A1(n1914), .A2(n1913), .A3(n1912), .ZN(n1864) );
  NAND3_X1 U1156 ( .A1(n1974), .A2(n1973), .A3(n1972), .ZN(n1924) );
  NAND2_X1 U1157 ( .A1(n2134), .A2(n2132), .ZN(n1976) );
  NAND2_X1 U1158 ( .A1(n1971), .A2(n1973), .ZN(n1917) );
  INV_X1 U1159 ( .A(n1547), .ZN(n1546) );
  INV_X1 U1160 ( .A(n1541), .ZN(n1540) );
  INV_X1 U1161 ( .A(n1543), .ZN(n1542) );
  INV_X1 U1162 ( .A(n1545), .ZN(n1544) );
  INV_X1 U1163 ( .A(n1555), .ZN(n1554) );
  OR2_X1 U1164 ( .A1(n2132), .A2(n2131), .ZN(n1535) );
  NAND2_X1 U1165 ( .A1(A[0]), .A2(n2111), .ZN(n1561) );
  INV_X1 U1166 ( .A(A[5]), .ZN(n1553) );
  INV_X1 U1167 ( .A(A[11]), .ZN(n1549) );
  INV_X1 U1168 ( .A(A[8]), .ZN(n1551) );
  INV_X1 U1169 ( .A(A[14]), .ZN(n1547) );
  INV_X1 U1170 ( .A(A[17]), .ZN(n1545) );
  INV_X1 U1171 ( .A(A[23]), .ZN(n1541) );
  INV_X1 U1172 ( .A(A[20]), .ZN(n1543) );
  NOR2_X4 U1173 ( .A1(n1670), .A2(n1671), .ZN(n1581) );
  NOR2_X4 U1174 ( .A1(n1672), .A2(n1673), .ZN(n1582) );
  NAND2_X2 U1175 ( .A1(n1670), .A2(n1672), .ZN(n1576) );
  NOR2_X4 U1176 ( .A1(n1731), .A2(n1732), .ZN(n1680) );
  NOR2_X4 U1177 ( .A1(n1733), .A2(n1734), .ZN(n1681) );
  NOR2_X4 U1178 ( .A1(n1791), .A2(n1792), .ZN(n1740) );
  NOR2_X4 U1179 ( .A1(n1793), .A2(n1794), .ZN(n1741) );
  NOR2_X4 U1180 ( .A1(n1851), .A2(n1852), .ZN(n1800) );
  NOR2_X4 U1181 ( .A1(n1853), .A2(n1854), .ZN(n1801) );
  NOR2_X4 U1182 ( .A1(n1911), .A2(n1912), .ZN(n1860) );
  NOR2_X4 U1183 ( .A1(n1913), .A2(n1914), .ZN(n1861) );
  NOR2_X4 U1184 ( .A1(n1971), .A2(n1972), .ZN(n1920) );
  NOR2_X4 U1185 ( .A1(n1973), .A2(n1974), .ZN(n1921) );
  INV_X2 U1186 ( .A(B[0]), .ZN(n1574) );
  NOR2_X4 U1187 ( .A1(n2112), .A2(n2111), .ZN(n1558) );
  NOR2_X4 U1188 ( .A1(n2113), .A2(A[0]), .ZN(n1559) );
  INV_X1 U1189 ( .A(B[23]), .ZN(n1555) );
  INV_X1 U1190 ( .A(B[23]), .ZN(n1556) );
  XNOR2_X1 U1191 ( .A(A[2]), .B(n1557), .ZN(n908) );
  AOI221_X1 U1192 ( .B1(B[22]), .B2(n1558), .C1(B[21]), .C2(n1559), .A(n1560), 
        .ZN(n1557) );
  OAI22_X1 U1193 ( .A1(n1561), .A2(n1562), .B1(n1563), .B2(n1564), .ZN(n1560)
         );
  XNOR2_X1 U1194 ( .A(A[2]), .B(n1565), .ZN(n907) );
  AOI221_X1 U1195 ( .B1(B[23]), .B2(n1558), .C1(n1559), .C2(B[22]), .A(n1566), 
        .ZN(n1565) );
  OAI22_X1 U1196 ( .A1(n1561), .A2(n1567), .B1(n1568), .B2(n1563), .ZN(n1566)
         );
  XNOR2_X1 U1197 ( .A(A[2]), .B(n1569), .ZN(n906) );
  AOI221_X1 U1198 ( .B1(B[23]), .B2(n1558), .C1(n1554), .C2(n1559), .A(n1570), 
        .ZN(n1569) );
  OAI22_X1 U1199 ( .A1(n1561), .A2(n1571), .B1(n1572), .B2(n1563), .ZN(n1570)
         );
  XNOR2_X1 U1200 ( .A(n1573), .B(n1553), .ZN(n904) );
  OAI22_X1 U1201 ( .A1(n1574), .A2(n1575), .B1(n1576), .B2(n1574), .ZN(n1573)
         );
  XNOR2_X1 U1202 ( .A(n1577), .B(n1553), .ZN(n903) );
  OAI222_X1 U1203 ( .A1(n1575), .A2(n1578), .B1(n1574), .B2(n1579), .C1(n1576), 
        .C2(n1580), .ZN(n1577) );
  INV_X1 U1204 ( .A(n1581), .ZN(n1579) );
  INV_X1 U1205 ( .A(n1582), .ZN(n1575) );
  XNOR2_X1 U1206 ( .A(n1552), .B(n1583), .ZN(n902) );
  AOI221_X1 U1207 ( .B1(B[2]), .B2(n1582), .C1(B[1]), .C2(n1581), .A(n1584), 
        .ZN(n1583) );
  OAI22_X1 U1208 ( .A1(n1576), .A2(n1585), .B1(n1574), .B2(n1586), .ZN(n1584)
         );
  XNOR2_X1 U1209 ( .A(n1552), .B(n1587), .ZN(n901) );
  AOI221_X1 U1210 ( .B1(B[3]), .B2(n1582), .C1(B[2]), .C2(n1581), .A(n1588), 
        .ZN(n1587) );
  OAI22_X1 U1211 ( .A1(n1576), .A2(n1589), .B1(n1578), .B2(n1586), .ZN(n1588)
         );
  XNOR2_X1 U1212 ( .A(n1552), .B(n1590), .ZN(n900) );
  AOI221_X1 U1213 ( .B1(B[4]), .B2(n1582), .C1(B[3]), .C2(n1581), .A(n1591), 
        .ZN(n1590) );
  OAI22_X1 U1214 ( .A1(n1576), .A2(n1592), .B1(n1593), .B2(n1586), .ZN(n1591)
         );
  XNOR2_X1 U1215 ( .A(n1552), .B(n1594), .ZN(n899) );
  AOI221_X1 U1216 ( .B1(B[5]), .B2(n1582), .C1(B[4]), .C2(n1581), .A(n1595), 
        .ZN(n1594) );
  OAI22_X1 U1217 ( .A1(n1576), .A2(n1596), .B1(n1586), .B2(n1597), .ZN(n1595)
         );
  XNOR2_X1 U1218 ( .A(n1552), .B(n1598), .ZN(n898) );
  AOI221_X1 U1219 ( .B1(B[6]), .B2(n1582), .C1(B[5]), .C2(n1581), .A(n1599), 
        .ZN(n1598) );
  OAI22_X1 U1220 ( .A1(n1576), .A2(n1600), .B1(n1586), .B2(n1601), .ZN(n1599)
         );
  XNOR2_X1 U1221 ( .A(n1552), .B(n1602), .ZN(n897) );
  AOI221_X1 U1222 ( .B1(B[7]), .B2(n1582), .C1(B[6]), .C2(n1581), .A(n1603), 
        .ZN(n1602) );
  OAI22_X1 U1223 ( .A1(n1576), .A2(n1604), .B1(n1586), .B2(n1605), .ZN(n1603)
         );
  XNOR2_X1 U1224 ( .A(n1552), .B(n1606), .ZN(n896) );
  AOI221_X1 U1225 ( .B1(B[8]), .B2(n1582), .C1(B[7]), .C2(n1581), .A(n1607), 
        .ZN(n1606) );
  OAI22_X1 U1226 ( .A1(n1576), .A2(n1608), .B1(n1586), .B2(n1609), .ZN(n1607)
         );
  XNOR2_X1 U1227 ( .A(n1552), .B(n1610), .ZN(n895) );
  AOI221_X1 U1228 ( .B1(B[9]), .B2(n1582), .C1(B[8]), .C2(n1581), .A(n1611), 
        .ZN(n1610) );
  OAI22_X1 U1229 ( .A1(n1576), .A2(n1612), .B1(n1586), .B2(n1613), .ZN(n1611)
         );
  XNOR2_X1 U1230 ( .A(n1552), .B(n1614), .ZN(n894) );
  AOI221_X1 U1231 ( .B1(B[10]), .B2(n1582), .C1(B[9]), .C2(n1581), .A(n1615), 
        .ZN(n1614) );
  OAI22_X1 U1232 ( .A1(n1576), .A2(n1616), .B1(n1586), .B2(n1617), .ZN(n1615)
         );
  XNOR2_X1 U1233 ( .A(n1552), .B(n1618), .ZN(n893) );
  AOI221_X1 U1234 ( .B1(B[11]), .B2(n1582), .C1(B[10]), .C2(n1581), .A(n1619), 
        .ZN(n1618) );
  OAI22_X1 U1235 ( .A1(n1576), .A2(n1620), .B1(n1586), .B2(n1621), .ZN(n1619)
         );
  XNOR2_X1 U1236 ( .A(n1552), .B(n1622), .ZN(n892) );
  AOI221_X1 U1237 ( .B1(B[12]), .B2(n1582), .C1(B[11]), .C2(n1581), .A(n1623), 
        .ZN(n1622) );
  OAI22_X1 U1238 ( .A1(n1576), .A2(n1624), .B1(n1586), .B2(n1625), .ZN(n1623)
         );
  XNOR2_X1 U1239 ( .A(n1552), .B(n1626), .ZN(n891) );
  AOI221_X1 U1240 ( .B1(B[13]), .B2(n1582), .C1(B[12]), .C2(n1581), .A(n1627), 
        .ZN(n1626) );
  OAI22_X1 U1241 ( .A1(n1576), .A2(n1628), .B1(n1586), .B2(n1629), .ZN(n1627)
         );
  XNOR2_X1 U1242 ( .A(n1552), .B(n1630), .ZN(n890) );
  AOI221_X1 U1243 ( .B1(B[14]), .B2(n1582), .C1(B[13]), .C2(n1581), .A(n1631), 
        .ZN(n1630) );
  OAI22_X1 U1244 ( .A1(n1576), .A2(n1632), .B1(n1586), .B2(n1633), .ZN(n1631)
         );
  XNOR2_X1 U1245 ( .A(n1552), .B(n1634), .ZN(n889) );
  AOI221_X1 U1246 ( .B1(B[15]), .B2(n1582), .C1(B[14]), .C2(n1581), .A(n1635), 
        .ZN(n1634) );
  OAI22_X1 U1247 ( .A1(n1576), .A2(n1636), .B1(n1586), .B2(n1637), .ZN(n1635)
         );
  XNOR2_X1 U1248 ( .A(n1552), .B(n1638), .ZN(n888) );
  AOI221_X1 U1249 ( .B1(B[16]), .B2(n1582), .C1(B[15]), .C2(n1581), .A(n1639), 
        .ZN(n1638) );
  OAI22_X1 U1250 ( .A1(n1576), .A2(n1640), .B1(n1586), .B2(n1641), .ZN(n1639)
         );
  XNOR2_X1 U1251 ( .A(n1552), .B(n1642), .ZN(n887) );
  AOI221_X1 U1252 ( .B1(B[17]), .B2(n1582), .C1(B[16]), .C2(n1581), .A(n1643), 
        .ZN(n1642) );
  OAI22_X1 U1253 ( .A1(n1576), .A2(n1644), .B1(n1586), .B2(n1645), .ZN(n1643)
         );
  XNOR2_X1 U1254 ( .A(n1552), .B(n1646), .ZN(n886) );
  AOI221_X1 U1255 ( .B1(B[18]), .B2(n1582), .C1(B[17]), .C2(n1581), .A(n1647), 
        .ZN(n1646) );
  OAI22_X1 U1256 ( .A1(n1576), .A2(n1648), .B1(n1586), .B2(n1649), .ZN(n1647)
         );
  XNOR2_X1 U1257 ( .A(n1552), .B(n1650), .ZN(n885) );
  AOI221_X1 U1258 ( .B1(B[19]), .B2(n1582), .C1(B[18]), .C2(n1581), .A(n1651), 
        .ZN(n1650) );
  OAI22_X1 U1259 ( .A1(n1576), .A2(n1652), .B1(n1586), .B2(n1653), .ZN(n1651)
         );
  XNOR2_X1 U1260 ( .A(A[5]), .B(n1654), .ZN(n884) );
  AOI221_X1 U1261 ( .B1(n1582), .B2(B[20]), .C1(B[19]), .C2(n1581), .A(n1655), 
        .ZN(n1654) );
  OAI22_X1 U1262 ( .A1(n1576), .A2(n1656), .B1(n1586), .B2(n1657), .ZN(n1655)
         );
  XNOR2_X1 U1263 ( .A(A[5]), .B(n1658), .ZN(n883) );
  AOI221_X1 U1264 ( .B1(n1582), .B2(B[21]), .C1(n1581), .C2(B[20]), .A(n1659), 
        .ZN(n1658) );
  OAI22_X1 U1265 ( .A1(n1576), .A2(n1660), .B1(n1586), .B2(n1661), .ZN(n1659)
         );
  XNOR2_X1 U1266 ( .A(A[5]), .B(n1662), .ZN(n882) );
  AOI221_X1 U1267 ( .B1(n1582), .B2(B[22]), .C1(n1581), .C2(B[21]), .A(n1663), 
        .ZN(n1662) );
  OAI22_X1 U1268 ( .A1(n1562), .A2(n1576), .B1(n1564), .B2(n1586), .ZN(n1663)
         );
  XNOR2_X1 U1269 ( .A(A[5]), .B(n1664), .ZN(n881) );
  AOI221_X1 U1270 ( .B1(n1582), .B2(B[23]), .C1(n1581), .C2(B[22]), .A(n1665), 
        .ZN(n1664) );
  OAI22_X1 U1271 ( .A1(n1567), .A2(n1576), .B1(n1568), .B2(n1586), .ZN(n1665)
         );
  XNOR2_X1 U1272 ( .A(A[5]), .B(n1666), .ZN(n880) );
  AOI221_X1 U1273 ( .B1(n1582), .B2(B[23]), .C1(n1581), .C2(n1554), .A(n1667), 
        .ZN(n1666) );
  OAI22_X1 U1274 ( .A1(n1571), .A2(n1576), .B1(n1572), .B2(n1586), .ZN(n1667)
         );
  XNOR2_X1 U1275 ( .A(n1552), .B(n1668), .ZN(n879) );
  OAI221_X1 U1276 ( .B1(n1556), .B2(n1586), .C1(n1556), .C2(n1576), .A(n1669), 
        .ZN(n1668) );
  OAI21_X1 U1277 ( .B1(n1582), .B2(n1581), .A(n1554), .ZN(n1669) );
  INV_X1 U1278 ( .A(n1673), .ZN(n1670) );
  XNOR2_X1 U1279 ( .A(A[3]), .B(A[4]), .ZN(n1671) );
  XNOR2_X1 U1280 ( .A(A[4]), .B(n1553), .ZN(n1672) );
  XOR2_X1 U1281 ( .A(A[3]), .B(n1674), .Z(n1673) );
  XNOR2_X1 U1282 ( .A(n1675), .B(n1551), .ZN(n878) );
  OAI22_X1 U1283 ( .A1(n1574), .A2(n1676), .B1(n1574), .B2(n1677), .ZN(n1675)
         );
  XNOR2_X1 U1284 ( .A(n1678), .B(n1551), .ZN(n877) );
  OAI222_X1 U1285 ( .A1(n1578), .A2(n1676), .B1(n1574), .B2(n1679), .C1(n1580), 
        .C2(n1677), .ZN(n1678) );
  INV_X1 U1286 ( .A(n1680), .ZN(n1679) );
  INV_X1 U1287 ( .A(n1681), .ZN(n1676) );
  XNOR2_X1 U1288 ( .A(n1550), .B(n1682), .ZN(n876) );
  AOI221_X1 U1289 ( .B1(n1681), .B2(B[2]), .C1(n1680), .C2(B[1]), .A(n1683), 
        .ZN(n1682) );
  OAI22_X1 U1290 ( .A1(n1585), .A2(n1677), .B1(n1574), .B2(n1684), .ZN(n1683)
         );
  XNOR2_X1 U1291 ( .A(n1550), .B(n1685), .ZN(n875) );
  AOI221_X1 U1292 ( .B1(n1681), .B2(B[3]), .C1(n1680), .C2(B[2]), .A(n1686), 
        .ZN(n1685) );
  OAI22_X1 U1293 ( .A1(n1589), .A2(n1677), .B1(n1578), .B2(n1684), .ZN(n1686)
         );
  XNOR2_X1 U1294 ( .A(n1550), .B(n1687), .ZN(n874) );
  AOI221_X1 U1295 ( .B1(n1681), .B2(B[4]), .C1(n1680), .C2(B[3]), .A(n1688), 
        .ZN(n1687) );
  OAI22_X1 U1296 ( .A1(n1592), .A2(n1677), .B1(n1593), .B2(n1684), .ZN(n1688)
         );
  XNOR2_X1 U1297 ( .A(n1550), .B(n1689), .ZN(n873) );
  AOI221_X1 U1298 ( .B1(n1681), .B2(B[5]), .C1(n1680), .C2(B[4]), .A(n1690), 
        .ZN(n1689) );
  OAI22_X1 U1299 ( .A1(n1596), .A2(n1677), .B1(n1597), .B2(n1684), .ZN(n1690)
         );
  XNOR2_X1 U1300 ( .A(n1550), .B(n1691), .ZN(n872) );
  AOI221_X1 U1301 ( .B1(n1681), .B2(B[6]), .C1(n1680), .C2(B[5]), .A(n1692), 
        .ZN(n1691) );
  OAI22_X1 U1302 ( .A1(n1600), .A2(n1677), .B1(n1601), .B2(n1684), .ZN(n1692)
         );
  XNOR2_X1 U1303 ( .A(n1550), .B(n1693), .ZN(n871) );
  AOI221_X1 U1304 ( .B1(n1681), .B2(B[7]), .C1(n1680), .C2(B[6]), .A(n1694), 
        .ZN(n1693) );
  OAI22_X1 U1305 ( .A1(n1604), .A2(n1677), .B1(n1605), .B2(n1684), .ZN(n1694)
         );
  XNOR2_X1 U1306 ( .A(n1550), .B(n1695), .ZN(n870) );
  AOI221_X1 U1307 ( .B1(n1681), .B2(B[8]), .C1(n1680), .C2(B[7]), .A(n1696), 
        .ZN(n1695) );
  OAI22_X1 U1308 ( .A1(n1608), .A2(n1677), .B1(n1609), .B2(n1684), .ZN(n1696)
         );
  XNOR2_X1 U1309 ( .A(n1550), .B(n1697), .ZN(n869) );
  AOI221_X1 U1310 ( .B1(n1681), .B2(B[9]), .C1(n1680), .C2(B[8]), .A(n1698), 
        .ZN(n1697) );
  OAI22_X1 U1311 ( .A1(n1612), .A2(n1677), .B1(n1613), .B2(n1684), .ZN(n1698)
         );
  XNOR2_X1 U1312 ( .A(n1550), .B(n1699), .ZN(n868) );
  AOI221_X1 U1313 ( .B1(n1681), .B2(B[10]), .C1(n1680), .C2(B[9]), .A(n1700), 
        .ZN(n1699) );
  OAI22_X1 U1314 ( .A1(n1616), .A2(n1677), .B1(n1617), .B2(n1684), .ZN(n1700)
         );
  XNOR2_X1 U1315 ( .A(n1550), .B(n1701), .ZN(n867) );
  AOI221_X1 U1316 ( .B1(n1681), .B2(B[11]), .C1(n1680), .C2(B[10]), .A(n1702), 
        .ZN(n1701) );
  OAI22_X1 U1317 ( .A1(n1620), .A2(n1677), .B1(n1621), .B2(n1684), .ZN(n1702)
         );
  XNOR2_X1 U1318 ( .A(n1550), .B(n1703), .ZN(n866) );
  AOI221_X1 U1319 ( .B1(n1681), .B2(B[12]), .C1(n1680), .C2(B[11]), .A(n1704), 
        .ZN(n1703) );
  OAI22_X1 U1320 ( .A1(n1624), .A2(n1677), .B1(n1625), .B2(n1684), .ZN(n1704)
         );
  XNOR2_X1 U1321 ( .A(n1550), .B(n1705), .ZN(n865) );
  AOI221_X1 U1322 ( .B1(n1681), .B2(B[13]), .C1(n1680), .C2(B[12]), .A(n1706), 
        .ZN(n1705) );
  OAI22_X1 U1323 ( .A1(n1628), .A2(n1677), .B1(n1629), .B2(n1684), .ZN(n1706)
         );
  XNOR2_X1 U1324 ( .A(n1550), .B(n1707), .ZN(n864) );
  AOI221_X1 U1325 ( .B1(n1681), .B2(B[14]), .C1(n1680), .C2(B[13]), .A(n1708), 
        .ZN(n1707) );
  OAI22_X1 U1326 ( .A1(n1632), .A2(n1677), .B1(n1633), .B2(n1684), .ZN(n1708)
         );
  XNOR2_X1 U1327 ( .A(n1550), .B(n1709), .ZN(n863) );
  AOI221_X1 U1328 ( .B1(n1681), .B2(B[15]), .C1(n1680), .C2(B[14]), .A(n1710), 
        .ZN(n1709) );
  OAI22_X1 U1329 ( .A1(n1636), .A2(n1677), .B1(n1637), .B2(n1684), .ZN(n1710)
         );
  XNOR2_X1 U1330 ( .A(n1550), .B(n1711), .ZN(n862) );
  AOI221_X1 U1331 ( .B1(n1681), .B2(B[16]), .C1(n1680), .C2(B[15]), .A(n1712), 
        .ZN(n1711) );
  OAI22_X1 U1332 ( .A1(n1640), .A2(n1677), .B1(n1641), .B2(n1684), .ZN(n1712)
         );
  XNOR2_X1 U1333 ( .A(n1550), .B(n1713), .ZN(n861) );
  AOI221_X1 U1334 ( .B1(n1681), .B2(B[17]), .C1(n1680), .C2(B[16]), .A(n1714), 
        .ZN(n1713) );
  OAI22_X1 U1335 ( .A1(n1644), .A2(n1677), .B1(n1645), .B2(n1684), .ZN(n1714)
         );
  XNOR2_X1 U1336 ( .A(n1550), .B(n1715), .ZN(n860) );
  AOI221_X1 U1337 ( .B1(n1681), .B2(B[18]), .C1(n1680), .C2(B[17]), .A(n1716), 
        .ZN(n1715) );
  OAI22_X1 U1338 ( .A1(n1648), .A2(n1677), .B1(n1649), .B2(n1684), .ZN(n1716)
         );
  XNOR2_X1 U1339 ( .A(n1550), .B(n1717), .ZN(n859) );
  AOI221_X1 U1340 ( .B1(n1681), .B2(B[19]), .C1(n1680), .C2(B[18]), .A(n1718), 
        .ZN(n1717) );
  OAI22_X1 U1341 ( .A1(n1652), .A2(n1677), .B1(n1653), .B2(n1684), .ZN(n1718)
         );
  XNOR2_X1 U1342 ( .A(A[8]), .B(n1719), .ZN(n858) );
  AOI221_X1 U1343 ( .B1(n1681), .B2(B[20]), .C1(n1680), .C2(B[19]), .A(n1720), 
        .ZN(n1719) );
  OAI22_X1 U1344 ( .A1(n1656), .A2(n1677), .B1(n1657), .B2(n1684), .ZN(n1720)
         );
  XNOR2_X1 U1345 ( .A(A[8]), .B(n1721), .ZN(n857) );
  AOI221_X1 U1346 ( .B1(n1681), .B2(B[21]), .C1(n1680), .C2(B[20]), .A(n1722), 
        .ZN(n1721) );
  OAI22_X1 U1347 ( .A1(n1660), .A2(n1677), .B1(n1661), .B2(n1684), .ZN(n1722)
         );
  XNOR2_X1 U1348 ( .A(A[8]), .B(n1723), .ZN(n856) );
  AOI221_X1 U1349 ( .B1(n1681), .B2(B[22]), .C1(n1680), .C2(B[21]), .A(n1724), 
        .ZN(n1723) );
  OAI22_X1 U1350 ( .A1(n1562), .A2(n1677), .B1(n1564), .B2(n1684), .ZN(n1724)
         );
  XNOR2_X1 U1351 ( .A(A[8]), .B(n1725), .ZN(n855) );
  AOI221_X1 U1352 ( .B1(n1681), .B2(B[23]), .C1(n1680), .C2(B[22]), .A(n1726), 
        .ZN(n1725) );
  OAI22_X1 U1353 ( .A1(n1567), .A2(n1677), .B1(n1568), .B2(n1684), .ZN(n1726)
         );
  XNOR2_X1 U1354 ( .A(A[8]), .B(n1727), .ZN(n854) );
  AOI221_X1 U1355 ( .B1(n1681), .B2(B[23]), .C1(n1680), .C2(n1554), .A(n1728), 
        .ZN(n1727) );
  OAI22_X1 U1356 ( .A1(n1571), .A2(n1677), .B1(n1572), .B2(n1684), .ZN(n1728)
         );
  XNOR2_X1 U1357 ( .A(n1550), .B(n1729), .ZN(n853) );
  OAI221_X1 U1358 ( .B1(n1555), .B2(n1684), .C1(n1556), .C2(n1677), .A(n1730), 
        .ZN(n1729) );
  OAI21_X1 U1359 ( .B1(n1681), .B2(n1680), .A(n1554), .ZN(n1730) );
  INV_X1 U1360 ( .A(n1734), .ZN(n1731) );
  XNOR2_X1 U1361 ( .A(A[6]), .B(A[7]), .ZN(n1732) );
  XNOR2_X1 U1362 ( .A(A[7]), .B(n1551), .ZN(n1733) );
  XOR2_X1 U1363 ( .A(A[6]), .B(n1553), .Z(n1734) );
  XNOR2_X1 U1364 ( .A(n1735), .B(n1549), .ZN(n852) );
  OAI22_X1 U1365 ( .A1(n1574), .A2(n1736), .B1(n1574), .B2(n1737), .ZN(n1735)
         );
  XNOR2_X1 U1366 ( .A(n1738), .B(n1549), .ZN(n851) );
  OAI222_X1 U1367 ( .A1(n1578), .A2(n1736), .B1(n1574), .B2(n1739), .C1(n1580), 
        .C2(n1737), .ZN(n1738) );
  INV_X1 U1368 ( .A(n1740), .ZN(n1739) );
  INV_X1 U1369 ( .A(n1741), .ZN(n1736) );
  XNOR2_X1 U1370 ( .A(n1548), .B(n1742), .ZN(n850) );
  AOI221_X1 U1371 ( .B1(n1741), .B2(B[2]), .C1(n1740), .C2(B[1]), .A(n1743), 
        .ZN(n1742) );
  OAI22_X1 U1372 ( .A1(n1585), .A2(n1737), .B1(n1574), .B2(n1744), .ZN(n1743)
         );
  XNOR2_X1 U1373 ( .A(n1548), .B(n1745), .ZN(n849) );
  AOI221_X1 U1374 ( .B1(n1741), .B2(B[3]), .C1(n1740), .C2(B[2]), .A(n1746), 
        .ZN(n1745) );
  OAI22_X1 U1375 ( .A1(n1589), .A2(n1737), .B1(n1578), .B2(n1744), .ZN(n1746)
         );
  XNOR2_X1 U1376 ( .A(n1548), .B(n1747), .ZN(n848) );
  AOI221_X1 U1377 ( .B1(n1741), .B2(B[4]), .C1(n1740), .C2(B[3]), .A(n1748), 
        .ZN(n1747) );
  OAI22_X1 U1378 ( .A1(n1592), .A2(n1737), .B1(n1593), .B2(n1744), .ZN(n1748)
         );
  XNOR2_X1 U1379 ( .A(n1548), .B(n1749), .ZN(n847) );
  AOI221_X1 U1380 ( .B1(n1741), .B2(B[5]), .C1(n1740), .C2(B[4]), .A(n1750), 
        .ZN(n1749) );
  OAI22_X1 U1381 ( .A1(n1596), .A2(n1737), .B1(n1597), .B2(n1744), .ZN(n1750)
         );
  XNOR2_X1 U1382 ( .A(n1548), .B(n1751), .ZN(n846) );
  AOI221_X1 U1383 ( .B1(n1741), .B2(B[6]), .C1(n1740), .C2(B[5]), .A(n1752), 
        .ZN(n1751) );
  OAI22_X1 U1384 ( .A1(n1600), .A2(n1737), .B1(n1601), .B2(n1744), .ZN(n1752)
         );
  XNOR2_X1 U1385 ( .A(n1548), .B(n1753), .ZN(n845) );
  AOI221_X1 U1386 ( .B1(n1741), .B2(B[7]), .C1(n1740), .C2(B[6]), .A(n1754), 
        .ZN(n1753) );
  OAI22_X1 U1387 ( .A1(n1604), .A2(n1737), .B1(n1605), .B2(n1744), .ZN(n1754)
         );
  XNOR2_X1 U1388 ( .A(n1548), .B(n1755), .ZN(n844) );
  AOI221_X1 U1389 ( .B1(n1741), .B2(B[8]), .C1(n1740), .C2(B[7]), .A(n1756), 
        .ZN(n1755) );
  OAI22_X1 U1390 ( .A1(n1608), .A2(n1737), .B1(n1609), .B2(n1744), .ZN(n1756)
         );
  XNOR2_X1 U1391 ( .A(n1548), .B(n1757), .ZN(n843) );
  AOI221_X1 U1392 ( .B1(n1741), .B2(B[9]), .C1(n1740), .C2(B[8]), .A(n1758), 
        .ZN(n1757) );
  OAI22_X1 U1393 ( .A1(n1612), .A2(n1737), .B1(n1613), .B2(n1744), .ZN(n1758)
         );
  XNOR2_X1 U1394 ( .A(n1548), .B(n1759), .ZN(n842) );
  AOI221_X1 U1395 ( .B1(n1741), .B2(B[10]), .C1(n1740), .C2(B[9]), .A(n1760), 
        .ZN(n1759) );
  OAI22_X1 U1396 ( .A1(n1616), .A2(n1737), .B1(n1617), .B2(n1744), .ZN(n1760)
         );
  XNOR2_X1 U1397 ( .A(n1548), .B(n1761), .ZN(n841) );
  AOI221_X1 U1398 ( .B1(n1741), .B2(B[11]), .C1(n1740), .C2(B[10]), .A(n1762), 
        .ZN(n1761) );
  OAI22_X1 U1399 ( .A1(n1620), .A2(n1737), .B1(n1621), .B2(n1744), .ZN(n1762)
         );
  XNOR2_X1 U1400 ( .A(n1548), .B(n1763), .ZN(n840) );
  AOI221_X1 U1401 ( .B1(n1741), .B2(B[12]), .C1(n1740), .C2(B[11]), .A(n1764), 
        .ZN(n1763) );
  OAI22_X1 U1402 ( .A1(n1624), .A2(n1737), .B1(n1625), .B2(n1744), .ZN(n1764)
         );
  XNOR2_X1 U1403 ( .A(n1548), .B(n1765), .ZN(n839) );
  AOI221_X1 U1404 ( .B1(n1741), .B2(B[13]), .C1(n1740), .C2(B[12]), .A(n1766), 
        .ZN(n1765) );
  OAI22_X1 U1405 ( .A1(n1628), .A2(n1737), .B1(n1629), .B2(n1744), .ZN(n1766)
         );
  XNOR2_X1 U1406 ( .A(n1548), .B(n1767), .ZN(n838) );
  AOI221_X1 U1407 ( .B1(n1741), .B2(B[14]), .C1(n1740), .C2(B[13]), .A(n1768), 
        .ZN(n1767) );
  OAI22_X1 U1408 ( .A1(n1632), .A2(n1737), .B1(n1633), .B2(n1744), .ZN(n1768)
         );
  XNOR2_X1 U1409 ( .A(n1548), .B(n1769), .ZN(n837) );
  AOI221_X1 U1410 ( .B1(n1741), .B2(B[15]), .C1(n1740), .C2(B[14]), .A(n1770), 
        .ZN(n1769) );
  OAI22_X1 U1411 ( .A1(n1636), .A2(n1737), .B1(n1637), .B2(n1744), .ZN(n1770)
         );
  XNOR2_X1 U1412 ( .A(n1548), .B(n1771), .ZN(n836) );
  AOI221_X1 U1413 ( .B1(n1741), .B2(B[16]), .C1(n1740), .C2(B[15]), .A(n1772), 
        .ZN(n1771) );
  OAI22_X1 U1414 ( .A1(n1640), .A2(n1737), .B1(n1641), .B2(n1744), .ZN(n1772)
         );
  XNOR2_X1 U1415 ( .A(n1548), .B(n1773), .ZN(n835) );
  AOI221_X1 U1416 ( .B1(n1741), .B2(B[17]), .C1(n1740), .C2(B[16]), .A(n1774), 
        .ZN(n1773) );
  OAI22_X1 U1417 ( .A1(n1644), .A2(n1737), .B1(n1645), .B2(n1744), .ZN(n1774)
         );
  XNOR2_X1 U1418 ( .A(n1548), .B(n1775), .ZN(n834) );
  AOI221_X1 U1419 ( .B1(n1741), .B2(B[18]), .C1(n1740), .C2(B[17]), .A(n1776), 
        .ZN(n1775) );
  OAI22_X1 U1420 ( .A1(n1648), .A2(n1737), .B1(n1649), .B2(n1744), .ZN(n1776)
         );
  XNOR2_X1 U1421 ( .A(n1548), .B(n1777), .ZN(n833) );
  AOI221_X1 U1422 ( .B1(n1741), .B2(B[19]), .C1(n1740), .C2(B[18]), .A(n1778), 
        .ZN(n1777) );
  OAI22_X1 U1423 ( .A1(n1652), .A2(n1737), .B1(n1653), .B2(n1744), .ZN(n1778)
         );
  XNOR2_X1 U1424 ( .A(n1548), .B(n1779), .ZN(n832) );
  AOI221_X1 U1425 ( .B1(n1741), .B2(B[20]), .C1(n1740), .C2(B[19]), .A(n1780), 
        .ZN(n1779) );
  OAI22_X1 U1426 ( .A1(n1656), .A2(n1737), .B1(n1657), .B2(n1744), .ZN(n1780)
         );
  XNOR2_X1 U1427 ( .A(A[11]), .B(n1781), .ZN(n831) );
  AOI221_X1 U1428 ( .B1(n1741), .B2(B[21]), .C1(n1740), .C2(B[20]), .A(n1782), 
        .ZN(n1781) );
  OAI22_X1 U1429 ( .A1(n1660), .A2(n1737), .B1(n1661), .B2(n1744), .ZN(n1782)
         );
  XNOR2_X1 U1430 ( .A(A[11]), .B(n1783), .ZN(n830) );
  AOI221_X1 U1431 ( .B1(n1741), .B2(B[22]), .C1(n1740), .C2(B[21]), .A(n1784), 
        .ZN(n1783) );
  OAI22_X1 U1432 ( .A1(n1562), .A2(n1737), .B1(n1564), .B2(n1744), .ZN(n1784)
         );
  XNOR2_X1 U1433 ( .A(A[11]), .B(n1785), .ZN(n829) );
  AOI221_X1 U1434 ( .B1(n1741), .B2(B[23]), .C1(n1740), .C2(B[22]), .A(n1786), 
        .ZN(n1785) );
  OAI22_X1 U1435 ( .A1(n1567), .A2(n1737), .B1(n1568), .B2(n1744), .ZN(n1786)
         );
  XNOR2_X1 U1436 ( .A(A[11]), .B(n1787), .ZN(n828) );
  AOI221_X1 U1437 ( .B1(n1741), .B2(B[23]), .C1(n1740), .C2(n1554), .A(n1788), 
        .ZN(n1787) );
  OAI22_X1 U1438 ( .A1(n1571), .A2(n1737), .B1(n1572), .B2(n1744), .ZN(n1788)
         );
  XNOR2_X1 U1439 ( .A(A[11]), .B(n1789), .ZN(n827) );
  OAI221_X1 U1440 ( .B1(n1556), .B2(n1744), .C1(n1556), .C2(n1737), .A(n1790), 
        .ZN(n1789) );
  OAI21_X1 U1441 ( .B1(n1741), .B2(n1740), .A(n1554), .ZN(n1790) );
  INV_X1 U1442 ( .A(n1794), .ZN(n1791) );
  XNOR2_X1 U1443 ( .A(A[10]), .B(A[9]), .ZN(n1792) );
  XNOR2_X1 U1444 ( .A(A[10]), .B(n1549), .ZN(n1793) );
  XOR2_X1 U1445 ( .A(A[9]), .B(n1551), .Z(n1794) );
  XNOR2_X1 U1446 ( .A(n1795), .B(n1547), .ZN(n826) );
  OAI22_X1 U1447 ( .A1(n1574), .A2(n1796), .B1(n1574), .B2(n1797), .ZN(n1795)
         );
  XNOR2_X1 U1448 ( .A(n1798), .B(n1547), .ZN(n825) );
  OAI222_X1 U1449 ( .A1(n1578), .A2(n1796), .B1(n1574), .B2(n1799), .C1(n1580), 
        .C2(n1797), .ZN(n1798) );
  INV_X1 U1450 ( .A(n1800), .ZN(n1799) );
  INV_X1 U1451 ( .A(n1801), .ZN(n1796) );
  XNOR2_X1 U1452 ( .A(n1546), .B(n1802), .ZN(n824) );
  AOI221_X1 U1453 ( .B1(n1801), .B2(B[2]), .C1(n1800), .C2(B[1]), .A(n1803), 
        .ZN(n1802) );
  OAI22_X1 U1454 ( .A1(n1585), .A2(n1797), .B1(n1574), .B2(n1804), .ZN(n1803)
         );
  XNOR2_X1 U1455 ( .A(n1546), .B(n1805), .ZN(n823) );
  AOI221_X1 U1456 ( .B1(n1801), .B2(B[3]), .C1(n1800), .C2(B[2]), .A(n1806), 
        .ZN(n1805) );
  OAI22_X1 U1457 ( .A1(n1589), .A2(n1797), .B1(n1578), .B2(n1804), .ZN(n1806)
         );
  XNOR2_X1 U1458 ( .A(n1546), .B(n1807), .ZN(n822) );
  AOI221_X1 U1459 ( .B1(n1801), .B2(B[4]), .C1(n1800), .C2(B[3]), .A(n1808), 
        .ZN(n1807) );
  OAI22_X1 U1460 ( .A1(n1592), .A2(n1797), .B1(n1593), .B2(n1804), .ZN(n1808)
         );
  XNOR2_X1 U1461 ( .A(n1546), .B(n1809), .ZN(n821) );
  AOI221_X1 U1462 ( .B1(n1801), .B2(B[5]), .C1(n1800), .C2(B[4]), .A(n1810), 
        .ZN(n1809) );
  OAI22_X1 U1463 ( .A1(n1596), .A2(n1797), .B1(n1597), .B2(n1804), .ZN(n1810)
         );
  XNOR2_X1 U1464 ( .A(n1546), .B(n1811), .ZN(n820) );
  AOI221_X1 U1465 ( .B1(n1801), .B2(B[6]), .C1(n1800), .C2(B[5]), .A(n1812), 
        .ZN(n1811) );
  OAI22_X1 U1466 ( .A1(n1600), .A2(n1797), .B1(n1601), .B2(n1804), .ZN(n1812)
         );
  XNOR2_X1 U1467 ( .A(n1546), .B(n1813), .ZN(n819) );
  AOI221_X1 U1468 ( .B1(n1801), .B2(B[7]), .C1(n1800), .C2(B[6]), .A(n1814), 
        .ZN(n1813) );
  OAI22_X1 U1469 ( .A1(n1604), .A2(n1797), .B1(n1605), .B2(n1804), .ZN(n1814)
         );
  XNOR2_X1 U1470 ( .A(n1546), .B(n1815), .ZN(n818) );
  AOI221_X1 U1471 ( .B1(n1801), .B2(B[8]), .C1(n1800), .C2(B[7]), .A(n1816), 
        .ZN(n1815) );
  OAI22_X1 U1472 ( .A1(n1608), .A2(n1797), .B1(n1609), .B2(n1804), .ZN(n1816)
         );
  XNOR2_X1 U1473 ( .A(n1546), .B(n1817), .ZN(n817) );
  AOI221_X1 U1474 ( .B1(n1801), .B2(B[9]), .C1(n1800), .C2(B[8]), .A(n1818), 
        .ZN(n1817) );
  OAI22_X1 U1475 ( .A1(n1612), .A2(n1797), .B1(n1613), .B2(n1804), .ZN(n1818)
         );
  XNOR2_X1 U1476 ( .A(n1546), .B(n1819), .ZN(n816) );
  AOI221_X1 U1477 ( .B1(n1801), .B2(B[10]), .C1(n1800), .C2(B[9]), .A(n1820), 
        .ZN(n1819) );
  OAI22_X1 U1478 ( .A1(n1616), .A2(n1797), .B1(n1617), .B2(n1804), .ZN(n1820)
         );
  XNOR2_X1 U1479 ( .A(n1546), .B(n1821), .ZN(n815) );
  AOI221_X1 U1480 ( .B1(n1801), .B2(B[11]), .C1(n1800), .C2(B[10]), .A(n1822), 
        .ZN(n1821) );
  OAI22_X1 U1481 ( .A1(n1620), .A2(n1797), .B1(n1621), .B2(n1804), .ZN(n1822)
         );
  XNOR2_X1 U1482 ( .A(n1546), .B(n1823), .ZN(n814) );
  AOI221_X1 U1483 ( .B1(n1801), .B2(B[12]), .C1(n1800), .C2(B[11]), .A(n1824), 
        .ZN(n1823) );
  OAI22_X1 U1484 ( .A1(n1624), .A2(n1797), .B1(n1625), .B2(n1804), .ZN(n1824)
         );
  XNOR2_X1 U1485 ( .A(n1546), .B(n1825), .ZN(n813) );
  AOI221_X1 U1486 ( .B1(n1801), .B2(B[13]), .C1(n1800), .C2(B[12]), .A(n1826), 
        .ZN(n1825) );
  OAI22_X1 U1487 ( .A1(n1628), .A2(n1797), .B1(n1629), .B2(n1804), .ZN(n1826)
         );
  XNOR2_X1 U1488 ( .A(n1546), .B(n1827), .ZN(n812) );
  AOI221_X1 U1489 ( .B1(n1801), .B2(B[14]), .C1(n1800), .C2(B[13]), .A(n1828), 
        .ZN(n1827) );
  OAI22_X1 U1490 ( .A1(n1632), .A2(n1797), .B1(n1633), .B2(n1804), .ZN(n1828)
         );
  XNOR2_X1 U1491 ( .A(n1546), .B(n1829), .ZN(n811) );
  AOI221_X1 U1492 ( .B1(n1801), .B2(B[15]), .C1(n1800), .C2(B[14]), .A(n1830), 
        .ZN(n1829) );
  OAI22_X1 U1493 ( .A1(n1636), .A2(n1797), .B1(n1637), .B2(n1804), .ZN(n1830)
         );
  XNOR2_X1 U1494 ( .A(n1546), .B(n1831), .ZN(n810) );
  AOI221_X1 U1495 ( .B1(n1801), .B2(B[16]), .C1(n1800), .C2(B[15]), .A(n1832), 
        .ZN(n1831) );
  OAI22_X1 U1496 ( .A1(n1640), .A2(n1797), .B1(n1641), .B2(n1804), .ZN(n1832)
         );
  XNOR2_X1 U1497 ( .A(n1546), .B(n1833), .ZN(n809) );
  AOI221_X1 U1498 ( .B1(n1801), .B2(B[17]), .C1(n1800), .C2(B[16]), .A(n1834), 
        .ZN(n1833) );
  OAI22_X1 U1499 ( .A1(n1644), .A2(n1797), .B1(n1645), .B2(n1804), .ZN(n1834)
         );
  XNOR2_X1 U1500 ( .A(n1546), .B(n1835), .ZN(n808) );
  AOI221_X1 U1501 ( .B1(n1801), .B2(B[18]), .C1(n1800), .C2(B[17]), .A(n1836), 
        .ZN(n1835) );
  OAI22_X1 U1502 ( .A1(n1648), .A2(n1797), .B1(n1649), .B2(n1804), .ZN(n1836)
         );
  XNOR2_X1 U1503 ( .A(n1546), .B(n1837), .ZN(n807) );
  AOI221_X1 U1504 ( .B1(n1801), .B2(B[19]), .C1(n1800), .C2(B[18]), .A(n1838), 
        .ZN(n1837) );
  OAI22_X1 U1505 ( .A1(n1652), .A2(n1797), .B1(n1653), .B2(n1804), .ZN(n1838)
         );
  XNOR2_X1 U1506 ( .A(n1546), .B(n1839), .ZN(n806) );
  AOI221_X1 U1507 ( .B1(n1801), .B2(B[20]), .C1(n1800), .C2(B[19]), .A(n1840), 
        .ZN(n1839) );
  OAI22_X1 U1508 ( .A1(n1656), .A2(n1797), .B1(n1657), .B2(n1804), .ZN(n1840)
         );
  XNOR2_X1 U1509 ( .A(A[14]), .B(n1841), .ZN(n805) );
  AOI221_X1 U1510 ( .B1(n1801), .B2(B[21]), .C1(n1800), .C2(B[20]), .A(n1842), 
        .ZN(n1841) );
  OAI22_X1 U1511 ( .A1(n1660), .A2(n1797), .B1(n1661), .B2(n1804), .ZN(n1842)
         );
  XNOR2_X1 U1512 ( .A(A[14]), .B(n1843), .ZN(n804) );
  AOI221_X1 U1513 ( .B1(n1801), .B2(B[22]), .C1(n1800), .C2(B[21]), .A(n1844), 
        .ZN(n1843) );
  OAI22_X1 U1514 ( .A1(n1562), .A2(n1797), .B1(n1564), .B2(n1804), .ZN(n1844)
         );
  XNOR2_X1 U1515 ( .A(A[14]), .B(n1845), .ZN(n803) );
  AOI221_X1 U1516 ( .B1(n1801), .B2(B[23]), .C1(n1800), .C2(B[22]), .A(n1846), 
        .ZN(n1845) );
  OAI22_X1 U1517 ( .A1(n1567), .A2(n1797), .B1(n1568), .B2(n1804), .ZN(n1846)
         );
  XNOR2_X1 U1518 ( .A(A[14]), .B(n1847), .ZN(n802) );
  AOI221_X1 U1519 ( .B1(n1801), .B2(B[23]), .C1(n1800), .C2(n1554), .A(n1848), 
        .ZN(n1847) );
  OAI22_X1 U1520 ( .A1(n1571), .A2(n1797), .B1(n1572), .B2(n1804), .ZN(n1848)
         );
  XNOR2_X1 U1521 ( .A(A[14]), .B(n1849), .ZN(n801) );
  OAI221_X1 U1522 ( .B1(n1556), .B2(n1804), .C1(n1556), .C2(n1797), .A(n1850), 
        .ZN(n1849) );
  OAI21_X1 U1523 ( .B1(n1801), .B2(n1800), .A(n1554), .ZN(n1850) );
  INV_X1 U1524 ( .A(n1854), .ZN(n1851) );
  XNOR2_X1 U1525 ( .A(A[12]), .B(A[13]), .ZN(n1852) );
  XNOR2_X1 U1526 ( .A(A[13]), .B(n1547), .ZN(n1853) );
  XOR2_X1 U1527 ( .A(A[12]), .B(n1549), .Z(n1854) );
  XNOR2_X1 U1528 ( .A(n1855), .B(n1545), .ZN(n800) );
  OAI22_X1 U1529 ( .A1(n1574), .A2(n1856), .B1(n1574), .B2(n1857), .ZN(n1855)
         );
  XNOR2_X1 U1530 ( .A(n1858), .B(n1545), .ZN(n799) );
  OAI222_X1 U1531 ( .A1(n1578), .A2(n1856), .B1(n1574), .B2(n1859), .C1(n1580), 
        .C2(n1857), .ZN(n1858) );
  INV_X1 U1532 ( .A(n1860), .ZN(n1859) );
  INV_X1 U1533 ( .A(n1861), .ZN(n1856) );
  XNOR2_X1 U1534 ( .A(n1544), .B(n1862), .ZN(n798) );
  AOI221_X1 U1535 ( .B1(n1861), .B2(B[2]), .C1(n1860), .C2(B[1]), .A(n1863), 
        .ZN(n1862) );
  OAI22_X1 U1536 ( .A1(n1585), .A2(n1857), .B1(n1574), .B2(n1864), .ZN(n1863)
         );
  XNOR2_X1 U1537 ( .A(n1544), .B(n1865), .ZN(n797) );
  AOI221_X1 U1538 ( .B1(n1861), .B2(B[3]), .C1(n1860), .C2(B[2]), .A(n1866), 
        .ZN(n1865) );
  OAI22_X1 U1539 ( .A1(n1589), .A2(n1857), .B1(n1578), .B2(n1864), .ZN(n1866)
         );
  XNOR2_X1 U1540 ( .A(n1544), .B(n1867), .ZN(n796) );
  AOI221_X1 U1541 ( .B1(n1861), .B2(B[4]), .C1(n1860), .C2(B[3]), .A(n1868), 
        .ZN(n1867) );
  OAI22_X1 U1542 ( .A1(n1592), .A2(n1857), .B1(n1593), .B2(n1864), .ZN(n1868)
         );
  XNOR2_X1 U1543 ( .A(n1544), .B(n1869), .ZN(n795) );
  AOI221_X1 U1544 ( .B1(n1861), .B2(B[5]), .C1(n1860), .C2(B[4]), .A(n1870), 
        .ZN(n1869) );
  OAI22_X1 U1545 ( .A1(n1596), .A2(n1857), .B1(n1597), .B2(n1864), .ZN(n1870)
         );
  XNOR2_X1 U1546 ( .A(n1544), .B(n1871), .ZN(n794) );
  AOI221_X1 U1547 ( .B1(n1861), .B2(B[6]), .C1(n1860), .C2(B[5]), .A(n1872), 
        .ZN(n1871) );
  OAI22_X1 U1548 ( .A1(n1600), .A2(n1857), .B1(n1601), .B2(n1864), .ZN(n1872)
         );
  XNOR2_X1 U1549 ( .A(n1544), .B(n1873), .ZN(n793) );
  AOI221_X1 U1550 ( .B1(n1861), .B2(B[7]), .C1(n1860), .C2(B[6]), .A(n1874), 
        .ZN(n1873) );
  OAI22_X1 U1551 ( .A1(n1604), .A2(n1857), .B1(n1605), .B2(n1864), .ZN(n1874)
         );
  XNOR2_X1 U1552 ( .A(n1544), .B(n1875), .ZN(n792) );
  AOI221_X1 U1553 ( .B1(n1861), .B2(B[8]), .C1(n1860), .C2(B[7]), .A(n1876), 
        .ZN(n1875) );
  OAI22_X1 U1554 ( .A1(n1608), .A2(n1857), .B1(n1609), .B2(n1864), .ZN(n1876)
         );
  XNOR2_X1 U1555 ( .A(n1544), .B(n1877), .ZN(n791) );
  AOI221_X1 U1556 ( .B1(n1861), .B2(B[9]), .C1(n1860), .C2(B[8]), .A(n1878), 
        .ZN(n1877) );
  OAI22_X1 U1557 ( .A1(n1612), .A2(n1857), .B1(n1613), .B2(n1864), .ZN(n1878)
         );
  XNOR2_X1 U1558 ( .A(n1544), .B(n1879), .ZN(n790) );
  AOI221_X1 U1559 ( .B1(n1861), .B2(B[10]), .C1(n1860), .C2(B[9]), .A(n1880), 
        .ZN(n1879) );
  OAI22_X1 U1560 ( .A1(n1616), .A2(n1857), .B1(n1617), .B2(n1864), .ZN(n1880)
         );
  XNOR2_X1 U1561 ( .A(n1544), .B(n1881), .ZN(n789) );
  AOI221_X1 U1562 ( .B1(n1861), .B2(B[11]), .C1(n1860), .C2(B[10]), .A(n1882), 
        .ZN(n1881) );
  OAI22_X1 U1563 ( .A1(n1620), .A2(n1857), .B1(n1621), .B2(n1864), .ZN(n1882)
         );
  XNOR2_X1 U1564 ( .A(n1544), .B(n1883), .ZN(n788) );
  AOI221_X1 U1565 ( .B1(n1861), .B2(B[12]), .C1(n1860), .C2(B[11]), .A(n1884), 
        .ZN(n1883) );
  OAI22_X1 U1566 ( .A1(n1624), .A2(n1857), .B1(n1625), .B2(n1864), .ZN(n1884)
         );
  XNOR2_X1 U1567 ( .A(n1544), .B(n1885), .ZN(n787) );
  AOI221_X1 U1568 ( .B1(n1861), .B2(B[13]), .C1(n1860), .C2(B[12]), .A(n1886), 
        .ZN(n1885) );
  OAI22_X1 U1569 ( .A1(n1628), .A2(n1857), .B1(n1629), .B2(n1864), .ZN(n1886)
         );
  XNOR2_X1 U1570 ( .A(n1544), .B(n1887), .ZN(n786) );
  AOI221_X1 U1571 ( .B1(n1861), .B2(B[14]), .C1(n1860), .C2(B[13]), .A(n1888), 
        .ZN(n1887) );
  OAI22_X1 U1572 ( .A1(n1632), .A2(n1857), .B1(n1633), .B2(n1864), .ZN(n1888)
         );
  XNOR2_X1 U1573 ( .A(n1544), .B(n1889), .ZN(n785) );
  AOI221_X1 U1574 ( .B1(n1861), .B2(B[15]), .C1(n1860), .C2(B[14]), .A(n1890), 
        .ZN(n1889) );
  OAI22_X1 U1575 ( .A1(n1636), .A2(n1857), .B1(n1637), .B2(n1864), .ZN(n1890)
         );
  XNOR2_X1 U1576 ( .A(n1544), .B(n1891), .ZN(n784) );
  AOI221_X1 U1577 ( .B1(n1861), .B2(B[16]), .C1(n1860), .C2(B[15]), .A(n1892), 
        .ZN(n1891) );
  OAI22_X1 U1578 ( .A1(n1640), .A2(n1857), .B1(n1641), .B2(n1864), .ZN(n1892)
         );
  XNOR2_X1 U1579 ( .A(n1544), .B(n1893), .ZN(n783) );
  AOI221_X1 U1580 ( .B1(n1861), .B2(B[17]), .C1(n1860), .C2(B[16]), .A(n1894), 
        .ZN(n1893) );
  OAI22_X1 U1581 ( .A1(n1644), .A2(n1857), .B1(n1645), .B2(n1864), .ZN(n1894)
         );
  XNOR2_X1 U1582 ( .A(n1544), .B(n1895), .ZN(n782) );
  AOI221_X1 U1583 ( .B1(n1861), .B2(B[18]), .C1(n1860), .C2(B[17]), .A(n1896), 
        .ZN(n1895) );
  OAI22_X1 U1584 ( .A1(n1648), .A2(n1857), .B1(n1649), .B2(n1864), .ZN(n1896)
         );
  XNOR2_X1 U1585 ( .A(n1544), .B(n1897), .ZN(n781) );
  AOI221_X1 U1586 ( .B1(n1861), .B2(B[19]), .C1(n1860), .C2(B[18]), .A(n1898), 
        .ZN(n1897) );
  OAI22_X1 U1587 ( .A1(n1652), .A2(n1857), .B1(n1653), .B2(n1864), .ZN(n1898)
         );
  XNOR2_X1 U1588 ( .A(n1544), .B(n1899), .ZN(n780) );
  AOI221_X1 U1589 ( .B1(n1861), .B2(B[20]), .C1(n1860), .C2(B[19]), .A(n1900), 
        .ZN(n1899) );
  OAI22_X1 U1590 ( .A1(n1656), .A2(n1857), .B1(n1657), .B2(n1864), .ZN(n1900)
         );
  XNOR2_X1 U1591 ( .A(A[17]), .B(n1901), .ZN(n779) );
  AOI221_X1 U1592 ( .B1(n1861), .B2(B[21]), .C1(n1860), .C2(B[20]), .A(n1902), 
        .ZN(n1901) );
  OAI22_X1 U1593 ( .A1(n1660), .A2(n1857), .B1(n1661), .B2(n1864), .ZN(n1902)
         );
  XNOR2_X1 U1594 ( .A(A[17]), .B(n1903), .ZN(n778) );
  AOI221_X1 U1595 ( .B1(n1861), .B2(B[22]), .C1(n1860), .C2(B[21]), .A(n1904), 
        .ZN(n1903) );
  OAI22_X1 U1596 ( .A1(n1562), .A2(n1857), .B1(n1564), .B2(n1864), .ZN(n1904)
         );
  XNOR2_X1 U1597 ( .A(A[17]), .B(n1905), .ZN(n777) );
  AOI221_X1 U1598 ( .B1(n1861), .B2(B[23]), .C1(n1860), .C2(B[22]), .A(n1906), 
        .ZN(n1905) );
  OAI22_X1 U1599 ( .A1(n1567), .A2(n1857), .B1(n1568), .B2(n1864), .ZN(n1906)
         );
  XNOR2_X1 U1600 ( .A(A[17]), .B(n1907), .ZN(n776) );
  AOI221_X1 U1601 ( .B1(n1861), .B2(B[23]), .C1(n1860), .C2(n1554), .A(n1908), 
        .ZN(n1907) );
  OAI22_X1 U1602 ( .A1(n1571), .A2(n1857), .B1(n1572), .B2(n1864), .ZN(n1908)
         );
  XNOR2_X1 U1603 ( .A(A[17]), .B(n1909), .ZN(n775) );
  OAI221_X1 U1604 ( .B1(n1556), .B2(n1864), .C1(n1556), .C2(n1857), .A(n1910), 
        .ZN(n1909) );
  OAI21_X1 U1605 ( .B1(n1861), .B2(n1860), .A(n1554), .ZN(n1910) );
  INV_X1 U1606 ( .A(n1914), .ZN(n1911) );
  XNOR2_X1 U1607 ( .A(A[15]), .B(A[16]), .ZN(n1912) );
  XNOR2_X1 U1608 ( .A(A[16]), .B(n1545), .ZN(n1913) );
  XOR2_X1 U1609 ( .A(A[15]), .B(n1547), .Z(n1914) );
  XNOR2_X1 U1610 ( .A(n1915), .B(n1543), .ZN(n774) );
  OAI22_X1 U1611 ( .A1(n1574), .A2(n1916), .B1(n1574), .B2(n1917), .ZN(n1915)
         );
  XNOR2_X1 U1612 ( .A(n1918), .B(n1543), .ZN(n773) );
  OAI222_X1 U1613 ( .A1(n1578), .A2(n1916), .B1(n1574), .B2(n1919), .C1(n1580), 
        .C2(n1917), .ZN(n1918) );
  INV_X1 U1614 ( .A(n1920), .ZN(n1919) );
  INV_X1 U1615 ( .A(n1921), .ZN(n1916) );
  XNOR2_X1 U1616 ( .A(n1542), .B(n1922), .ZN(n772) );
  AOI221_X1 U1617 ( .B1(n1921), .B2(B[2]), .C1(n1920), .C2(B[1]), .A(n1923), 
        .ZN(n1922) );
  OAI22_X1 U1618 ( .A1(n1585), .A2(n1917), .B1(n1574), .B2(n1924), .ZN(n1923)
         );
  XNOR2_X1 U1619 ( .A(n1542), .B(n1925), .ZN(n771) );
  AOI221_X1 U1620 ( .B1(n1921), .B2(B[3]), .C1(n1920), .C2(B[2]), .A(n1926), 
        .ZN(n1925) );
  OAI22_X1 U1621 ( .A1(n1589), .A2(n1917), .B1(n1578), .B2(n1924), .ZN(n1926)
         );
  XNOR2_X1 U1622 ( .A(n1542), .B(n1927), .ZN(n770) );
  AOI221_X1 U1623 ( .B1(n1921), .B2(B[4]), .C1(n1920), .C2(B[3]), .A(n1928), 
        .ZN(n1927) );
  OAI22_X1 U1624 ( .A1(n1592), .A2(n1917), .B1(n1593), .B2(n1924), .ZN(n1928)
         );
  XNOR2_X1 U1625 ( .A(n1542), .B(n1929), .ZN(n769) );
  AOI221_X1 U1626 ( .B1(n1921), .B2(B[5]), .C1(n1920), .C2(B[4]), .A(n1930), 
        .ZN(n1929) );
  OAI22_X1 U1627 ( .A1(n1596), .A2(n1917), .B1(n1597), .B2(n1924), .ZN(n1930)
         );
  XNOR2_X1 U1628 ( .A(n1542), .B(n1931), .ZN(n768) );
  AOI221_X1 U1629 ( .B1(n1921), .B2(B[6]), .C1(n1920), .C2(B[5]), .A(n1932), 
        .ZN(n1931) );
  OAI22_X1 U1630 ( .A1(n1600), .A2(n1917), .B1(n1601), .B2(n1924), .ZN(n1932)
         );
  XNOR2_X1 U1631 ( .A(n1542), .B(n1933), .ZN(n767) );
  AOI221_X1 U1632 ( .B1(n1921), .B2(B[7]), .C1(n1920), .C2(B[6]), .A(n1934), 
        .ZN(n1933) );
  OAI22_X1 U1633 ( .A1(n1604), .A2(n1917), .B1(n1605), .B2(n1924), .ZN(n1934)
         );
  XNOR2_X1 U1634 ( .A(n1542), .B(n1935), .ZN(n766) );
  AOI221_X1 U1635 ( .B1(n1921), .B2(B[8]), .C1(n1920), .C2(B[7]), .A(n1936), 
        .ZN(n1935) );
  OAI22_X1 U1636 ( .A1(n1608), .A2(n1917), .B1(n1609), .B2(n1924), .ZN(n1936)
         );
  XNOR2_X1 U1637 ( .A(n1542), .B(n1937), .ZN(n765) );
  AOI221_X1 U1638 ( .B1(n1921), .B2(B[9]), .C1(n1920), .C2(B[8]), .A(n1938), 
        .ZN(n1937) );
  OAI22_X1 U1639 ( .A1(n1612), .A2(n1917), .B1(n1613), .B2(n1924), .ZN(n1938)
         );
  XNOR2_X1 U1640 ( .A(n1542), .B(n1939), .ZN(n764) );
  AOI221_X1 U1641 ( .B1(n1921), .B2(B[10]), .C1(n1920), .C2(B[9]), .A(n1940), 
        .ZN(n1939) );
  OAI22_X1 U1642 ( .A1(n1616), .A2(n1917), .B1(n1617), .B2(n1924), .ZN(n1940)
         );
  XNOR2_X1 U1643 ( .A(n1542), .B(n1941), .ZN(n763) );
  AOI221_X1 U1644 ( .B1(n1921), .B2(B[11]), .C1(n1920), .C2(B[10]), .A(n1942), 
        .ZN(n1941) );
  OAI22_X1 U1645 ( .A1(n1620), .A2(n1917), .B1(n1621), .B2(n1924), .ZN(n1942)
         );
  XNOR2_X1 U1646 ( .A(n1542), .B(n1943), .ZN(n762) );
  AOI221_X1 U1647 ( .B1(n1921), .B2(B[12]), .C1(n1920), .C2(B[11]), .A(n1944), 
        .ZN(n1943) );
  OAI22_X1 U1648 ( .A1(n1624), .A2(n1917), .B1(n1625), .B2(n1924), .ZN(n1944)
         );
  XNOR2_X1 U1649 ( .A(n1542), .B(n1945), .ZN(n761) );
  AOI221_X1 U1650 ( .B1(n1921), .B2(B[13]), .C1(n1920), .C2(B[12]), .A(n1946), 
        .ZN(n1945) );
  OAI22_X1 U1651 ( .A1(n1628), .A2(n1917), .B1(n1629), .B2(n1924), .ZN(n1946)
         );
  XNOR2_X1 U1652 ( .A(n1542), .B(n1947), .ZN(n760) );
  AOI221_X1 U1653 ( .B1(n1921), .B2(B[14]), .C1(n1920), .C2(B[13]), .A(n1948), 
        .ZN(n1947) );
  OAI22_X1 U1654 ( .A1(n1632), .A2(n1917), .B1(n1633), .B2(n1924), .ZN(n1948)
         );
  XNOR2_X1 U1655 ( .A(n1542), .B(n1949), .ZN(n759) );
  AOI221_X1 U1656 ( .B1(n1921), .B2(B[15]), .C1(n1920), .C2(B[14]), .A(n1950), 
        .ZN(n1949) );
  OAI22_X1 U1657 ( .A1(n1636), .A2(n1917), .B1(n1637), .B2(n1924), .ZN(n1950)
         );
  XNOR2_X1 U1658 ( .A(n1542), .B(n1951), .ZN(n758) );
  AOI221_X1 U1659 ( .B1(n1921), .B2(B[16]), .C1(n1920), .C2(B[15]), .A(n1952), 
        .ZN(n1951) );
  OAI22_X1 U1660 ( .A1(n1640), .A2(n1917), .B1(n1641), .B2(n1924), .ZN(n1952)
         );
  XNOR2_X1 U1661 ( .A(n1542), .B(n1953), .ZN(n757) );
  AOI221_X1 U1662 ( .B1(n1921), .B2(B[17]), .C1(n1920), .C2(B[16]), .A(n1954), 
        .ZN(n1953) );
  OAI22_X1 U1663 ( .A1(n1644), .A2(n1917), .B1(n1645), .B2(n1924), .ZN(n1954)
         );
  XNOR2_X1 U1664 ( .A(n1542), .B(n1955), .ZN(n756) );
  AOI221_X1 U1665 ( .B1(n1921), .B2(B[18]), .C1(n1920), .C2(B[17]), .A(n1956), 
        .ZN(n1955) );
  OAI22_X1 U1666 ( .A1(n1648), .A2(n1917), .B1(n1649), .B2(n1924), .ZN(n1956)
         );
  XNOR2_X1 U1667 ( .A(n1542), .B(n1957), .ZN(n755) );
  AOI221_X1 U1668 ( .B1(n1921), .B2(B[19]), .C1(n1920), .C2(B[18]), .A(n1958), 
        .ZN(n1957) );
  OAI22_X1 U1669 ( .A1(n1652), .A2(n1917), .B1(n1653), .B2(n1924), .ZN(n1958)
         );
  XNOR2_X1 U1670 ( .A(n1542), .B(n1959), .ZN(n754) );
  AOI221_X1 U1671 ( .B1(n1921), .B2(B[20]), .C1(n1920), .C2(B[19]), .A(n1960), 
        .ZN(n1959) );
  OAI22_X1 U1672 ( .A1(n1656), .A2(n1917), .B1(n1657), .B2(n1924), .ZN(n1960)
         );
  XNOR2_X1 U1673 ( .A(A[20]), .B(n1961), .ZN(n753) );
  AOI221_X1 U1674 ( .B1(n1921), .B2(B[21]), .C1(n1920), .C2(B[20]), .A(n1962), 
        .ZN(n1961) );
  OAI22_X1 U1675 ( .A1(n1660), .A2(n1917), .B1(n1661), .B2(n1924), .ZN(n1962)
         );
  XNOR2_X1 U1676 ( .A(A[20]), .B(n1963), .ZN(n752) );
  AOI221_X1 U1677 ( .B1(n1921), .B2(B[22]), .C1(n1920), .C2(B[21]), .A(n1964), 
        .ZN(n1963) );
  OAI22_X1 U1678 ( .A1(n1562), .A2(n1917), .B1(n1564), .B2(n1924), .ZN(n1964)
         );
  XNOR2_X1 U1679 ( .A(A[20]), .B(n1965), .ZN(n751) );
  AOI221_X1 U1680 ( .B1(n1921), .B2(n1554), .C1(n1920), .C2(B[22]), .A(n1966), 
        .ZN(n1965) );
  OAI22_X1 U1681 ( .A1(n1567), .A2(n1917), .B1(n1568), .B2(n1924), .ZN(n1966)
         );
  XNOR2_X1 U1682 ( .A(A[20]), .B(n1967), .ZN(n750) );
  AOI221_X1 U1683 ( .B1(n1921), .B2(B[23]), .C1(n1920), .C2(n1554), .A(n1968), 
        .ZN(n1967) );
  OAI22_X1 U1684 ( .A1(n1571), .A2(n1917), .B1(n1572), .B2(n1924), .ZN(n1968)
         );
  XNOR2_X1 U1685 ( .A(A[20]), .B(n1969), .ZN(n749) );
  OAI221_X1 U1686 ( .B1(n1556), .B2(n1924), .C1(n1556), .C2(n1917), .A(n1970), 
        .ZN(n1969) );
  OAI21_X1 U1687 ( .B1(n1921), .B2(n1920), .A(n1554), .ZN(n1970) );
  INV_X1 U1688 ( .A(n1974), .ZN(n1971) );
  XNOR2_X1 U1689 ( .A(A[18]), .B(A[19]), .ZN(n1972) );
  XNOR2_X1 U1690 ( .A(A[19]), .B(n1543), .ZN(n1973) );
  XOR2_X1 U1691 ( .A(A[18]), .B(n1545), .Z(n1974) );
  XNOR2_X1 U1692 ( .A(n1975), .B(n1541), .ZN(n748) );
  OAI22_X1 U1693 ( .A1(n1574), .A2(n1535), .B1(n1574), .B2(n1976), .ZN(n1975)
         );
  XNOR2_X1 U1694 ( .A(n1977), .B(n1541), .ZN(n747) );
  OAI222_X1 U1695 ( .A1(n1578), .A2(n1535), .B1(n1574), .B2(n1534), .C1(n1580), 
        .C2(n1976), .ZN(n1977) );
  INV_X1 U1696 ( .A(n1397), .ZN(n1580) );
  XNOR2_X1 U1697 ( .A(n1540), .B(n1978), .ZN(n746) );
  AOI221_X1 U1698 ( .B1(n1537), .B2(B[2]), .C1(n1536), .C2(B[1]), .A(n1979), 
        .ZN(n1978) );
  OAI22_X1 U1699 ( .A1(n1585), .A2(n1976), .B1(n1574), .B2(n1538), .ZN(n1979)
         );
  INV_X1 U1700 ( .A(n1396), .ZN(n1585) );
  XNOR2_X1 U1701 ( .A(n1540), .B(n1981), .ZN(n745) );
  AOI221_X1 U1702 ( .B1(n1537), .B2(B[3]), .C1(n1536), .C2(B[2]), .A(n1982), 
        .ZN(n1981) );
  OAI22_X1 U1703 ( .A1(n1589), .A2(n1976), .B1(n1578), .B2(n1539), .ZN(n1982)
         );
  XNOR2_X1 U1704 ( .A(n1540), .B(n1983), .ZN(n744) );
  AOI221_X1 U1705 ( .B1(n1537), .B2(B[4]), .C1(n1536), .C2(B[3]), .A(n1984), 
        .ZN(n1983) );
  OAI22_X1 U1706 ( .A1(n1592), .A2(n1976), .B1(n1593), .B2(n1539), .ZN(n1984)
         );
  XNOR2_X1 U1707 ( .A(n1540), .B(n1985), .ZN(n743) );
  AOI221_X1 U1708 ( .B1(n1537), .B2(B[5]), .C1(n1536), .C2(B[4]), .A(n1986), 
        .ZN(n1985) );
  OAI22_X1 U1709 ( .A1(n1596), .A2(n1976), .B1(n1597), .B2(n1539), .ZN(n1986)
         );
  XNOR2_X1 U1710 ( .A(n1540), .B(n1987), .ZN(n742) );
  AOI221_X1 U1711 ( .B1(n1537), .B2(B[6]), .C1(n1536), .C2(B[5]), .A(n1988), 
        .ZN(n1987) );
  OAI22_X1 U1712 ( .A1(n1600), .A2(n1976), .B1(n1601), .B2(n1539), .ZN(n1988)
         );
  XNOR2_X1 U1713 ( .A(n1540), .B(n1989), .ZN(n741) );
  AOI221_X1 U1714 ( .B1(n1537), .B2(B[7]), .C1(n1536), .C2(B[6]), .A(n1990), 
        .ZN(n1989) );
  OAI22_X1 U1715 ( .A1(n1604), .A2(n1976), .B1(n1605), .B2(n1539), .ZN(n1990)
         );
  XNOR2_X1 U1716 ( .A(n1540), .B(n1991), .ZN(n740) );
  AOI221_X1 U1717 ( .B1(n1537), .B2(B[9]), .C1(n1536), .C2(B[8]), .A(n1992), 
        .ZN(n1991) );
  OAI22_X1 U1718 ( .A1(n1612), .A2(n1976), .B1(n1613), .B2(n1539), .ZN(n1992)
         );
  XNOR2_X1 U1719 ( .A(n1540), .B(n1993), .ZN(n739) );
  AOI221_X1 U1720 ( .B1(n1537), .B2(B[10]), .C1(n1536), .C2(B[9]), .A(n1994), 
        .ZN(n1993) );
  OAI22_X1 U1721 ( .A1(n1616), .A2(n1976), .B1(n1617), .B2(n1539), .ZN(n1994)
         );
  XNOR2_X1 U1722 ( .A(n1540), .B(n1995), .ZN(n738) );
  AOI221_X1 U1723 ( .B1(n1537), .B2(B[12]), .C1(n1536), .C2(B[11]), .A(n1996), 
        .ZN(n1995) );
  OAI22_X1 U1724 ( .A1(n1624), .A2(n1976), .B1(n1625), .B2(n1539), .ZN(n1996)
         );
  XNOR2_X1 U1725 ( .A(n1540), .B(n1997), .ZN(n737) );
  AOI221_X1 U1726 ( .B1(n1537), .B2(B[13]), .C1(n1536), .C2(B[12]), .A(n1998), 
        .ZN(n1997) );
  OAI22_X1 U1727 ( .A1(n1628), .A2(n1976), .B1(n1629), .B2(n1539), .ZN(n1998)
         );
  XNOR2_X1 U1728 ( .A(n1540), .B(n1999), .ZN(n736) );
  AOI221_X1 U1729 ( .B1(n1537), .B2(B[14]), .C1(n1536), .C2(B[13]), .A(n2000), 
        .ZN(n1999) );
  OAI22_X1 U1730 ( .A1(n1632), .A2(n1976), .B1(n1633), .B2(n1539), .ZN(n2000)
         );
  XNOR2_X1 U1731 ( .A(n1540), .B(n2001), .ZN(n735) );
  AOI221_X1 U1732 ( .B1(n1537), .B2(B[15]), .C1(n1536), .C2(B[14]), .A(n2002), 
        .ZN(n2001) );
  OAI22_X1 U1733 ( .A1(n1636), .A2(n1976), .B1(n1637), .B2(n1539), .ZN(n2002)
         );
  XNOR2_X1 U1734 ( .A(n1540), .B(n2003), .ZN(n734) );
  AOI221_X1 U1735 ( .B1(n1537), .B2(B[16]), .C1(n1536), .C2(B[15]), .A(n2004), 
        .ZN(n2003) );
  OAI22_X1 U1736 ( .A1(n1640), .A2(n1976), .B1(n1641), .B2(n1538), .ZN(n2004)
         );
  XNOR2_X1 U1737 ( .A(n1540), .B(n2005), .ZN(n733) );
  AOI221_X1 U1738 ( .B1(n1537), .B2(B[18]), .C1(n1536), .C2(B[17]), .A(n2006), 
        .ZN(n2005) );
  OAI22_X1 U1739 ( .A1(n1648), .A2(n1976), .B1(n1649), .B2(n1538), .ZN(n2006)
         );
  XNOR2_X1 U1740 ( .A(n1540), .B(n2007), .ZN(n732) );
  AOI221_X1 U1741 ( .B1(n1537), .B2(B[19]), .C1(n1536), .C2(B[18]), .A(n2008), 
        .ZN(n2007) );
  OAI22_X1 U1742 ( .A1(n1652), .A2(n1976), .B1(n1653), .B2(n1538), .ZN(n2008)
         );
  XNOR2_X1 U1743 ( .A(n1540), .B(n2009), .ZN(n731) );
  AOI221_X1 U1744 ( .B1(n1537), .B2(B[20]), .C1(n1536), .C2(B[19]), .A(n2010), 
        .ZN(n2009) );
  OAI22_X1 U1745 ( .A1(n1656), .A2(n1976), .B1(n1657), .B2(n1538), .ZN(n2010)
         );
  XNOR2_X1 U1746 ( .A(A[23]), .B(n2011), .ZN(n730) );
  AOI221_X1 U1747 ( .B1(n1537), .B2(B[21]), .C1(n1536), .C2(B[20]), .A(n2012), 
        .ZN(n2011) );
  OAI22_X1 U1748 ( .A1(n1660), .A2(n1976), .B1(n1661), .B2(n1538), .ZN(n2012)
         );
  XNOR2_X1 U1749 ( .A(A[23]), .B(n2013), .ZN(n729) );
  AOI221_X1 U1750 ( .B1(n1537), .B2(B[22]), .C1(n1536), .C2(B[21]), .A(n2014), 
        .ZN(n2013) );
  OAI22_X1 U1751 ( .A1(n1562), .A2(n1976), .B1(n1564), .B2(n1538), .ZN(n2014)
         );
  INV_X1 U1752 ( .A(B[20]), .ZN(n1564) );
  INV_X1 U1753 ( .A(n1376), .ZN(n1562) );
  XNOR2_X1 U1754 ( .A(n519), .B(n2015), .ZN(n506) );
  INV_X1 U1755 ( .A(n493), .ZN(n479) );
  NOR2_X1 U1756 ( .A1(n2015), .A2(n519), .ZN(n493) );
  XOR2_X1 U1757 ( .A(n2016), .B(n1674), .Z(n2015) );
  OAI221_X1 U1758 ( .B1(n1563), .B2(n1556), .C1(n1561), .C2(n1556), .A(n2017), 
        .ZN(n2016) );
  OAI21_X1 U1759 ( .B1(n1558), .B2(n1559), .A(n1554), .ZN(n2017) );
  INV_X1 U1760 ( .A(n454), .ZN(n442) );
  XOR2_X1 U1761 ( .A(n1540), .B(n2018), .Z(n454) );
  AOI221_X1 U1762 ( .B1(n1537), .B2(B[8]), .C1(n1536), .C2(B[7]), .A(n2019), 
        .ZN(n2018) );
  OAI22_X1 U1763 ( .A1(n1608), .A2(n1976), .B1(n1609), .B2(n1538), .ZN(n2019)
         );
  INV_X1 U1764 ( .A(n421), .ZN(n411) );
  XOR2_X1 U1765 ( .A(n1540), .B(n2020), .Z(n421) );
  AOI221_X1 U1766 ( .B1(n1537), .B2(B[11]), .C1(n1536), .C2(B[10]), .A(n2021), 
        .ZN(n2020) );
  OAI22_X1 U1767 ( .A1(n1620), .A2(n1976), .B1(n1621), .B2(n1538), .ZN(n2021)
         );
  INV_X1 U1768 ( .A(n387), .ZN(n395) );
  INV_X1 U1769 ( .A(n374), .ZN(n368) );
  XOR2_X1 U1770 ( .A(n1540), .B(n2022), .Z(n374) );
  AOI221_X1 U1771 ( .B1(n1537), .B2(B[17]), .C1(n1536), .C2(B[16]), .A(n2023), 
        .ZN(n2022) );
  OAI22_X1 U1772 ( .A1(n1644), .A2(n1976), .B1(n1645), .B2(n1538), .ZN(n2023)
         );
  INV_X1 U1773 ( .A(n356), .ZN(n360) );
  INV_X1 U1774 ( .A(n2024), .ZN(n351) );
  OAI222_X1 U1775 ( .A1(n2025), .A2(n2026), .B1(n2025), .B2(n2027), .C1(n2027), 
        .C2(n2026), .ZN(n326) );
  INV_X1 U1776 ( .A(n550), .ZN(n2027) );
  XNOR2_X1 U1777 ( .A(n1674), .B(n2028), .ZN(n2026) );
  AOI221_X1 U1778 ( .B1(B[21]), .B2(n1558), .C1(B[20]), .C2(n1559), .A(n2029), 
        .ZN(n2028) );
  OAI22_X1 U1779 ( .A1(n1561), .A2(n1660), .B1(n1563), .B2(n1661), .ZN(n2029)
         );
  INV_X1 U1780 ( .A(B[19]), .ZN(n1661) );
  INV_X1 U1781 ( .A(n1377), .ZN(n1660) );
  AOI222_X1 U1782 ( .A1(n2030), .A2(n2031), .B1(n2030), .B2(n564), .C1(n564), 
        .C2(n2031), .ZN(n2025) );
  XNOR2_X1 U1783 ( .A(A[2]), .B(n2032), .ZN(n2031) );
  AOI221_X1 U1784 ( .B1(B[20]), .B2(n1558), .C1(B[19]), .C2(n1559), .A(n2033), 
        .ZN(n2032) );
  OAI22_X1 U1785 ( .A1(n1561), .A2(n1656), .B1(n1563), .B2(n1657), .ZN(n2033)
         );
  INV_X1 U1786 ( .A(B[18]), .ZN(n1657) );
  INV_X1 U1787 ( .A(n1378), .ZN(n1656) );
  INV_X1 U1788 ( .A(n2034), .ZN(n2030) );
  AOI222_X1 U1789 ( .A1(n2035), .A2(n2036), .B1(n2035), .B2(n576), .C1(n576), 
        .C2(n2036), .ZN(n2034) );
  XNOR2_X1 U1790 ( .A(A[2]), .B(n2037), .ZN(n2036) );
  AOI221_X1 U1791 ( .B1(B[19]), .B2(n1558), .C1(B[18]), .C2(n1559), .A(n2038), 
        .ZN(n2037) );
  OAI22_X1 U1792 ( .A1(n1561), .A2(n1652), .B1(n1563), .B2(n1653), .ZN(n2038)
         );
  INV_X1 U1793 ( .A(B[17]), .ZN(n1653) );
  INV_X1 U1794 ( .A(n1379), .ZN(n1652) );
  OAI222_X1 U1795 ( .A1(n2039), .A2(n2040), .B1(n2039), .B2(n2041), .C1(n2041), 
        .C2(n2040), .ZN(n2035) );
  INV_X1 U1796 ( .A(n588), .ZN(n2041) );
  XNOR2_X1 U1797 ( .A(n1674), .B(n2042), .ZN(n2040) );
  AOI221_X1 U1798 ( .B1(B[18]), .B2(n1558), .C1(B[17]), .C2(n1559), .A(n2043), 
        .ZN(n2042) );
  OAI22_X1 U1799 ( .A1(n1561), .A2(n1648), .B1(n1563), .B2(n1649), .ZN(n2043)
         );
  INV_X1 U1800 ( .A(B[16]), .ZN(n1649) );
  INV_X1 U1801 ( .A(n1380), .ZN(n1648) );
  AOI222_X1 U1802 ( .A1(n2044), .A2(n2045), .B1(n2044), .B2(n600), .C1(n600), 
        .C2(n2045), .ZN(n2039) );
  XNOR2_X1 U1803 ( .A(A[2]), .B(n2046), .ZN(n2045) );
  AOI221_X1 U1804 ( .B1(B[17]), .B2(n1558), .C1(B[16]), .C2(n1559), .A(n2047), 
        .ZN(n2046) );
  OAI22_X1 U1805 ( .A1(n1561), .A2(n1644), .B1(n1563), .B2(n1645), .ZN(n2047)
         );
  INV_X1 U1806 ( .A(B[15]), .ZN(n1645) );
  INV_X1 U1807 ( .A(n1381), .ZN(n1644) );
  OAI222_X1 U1808 ( .A1(n2048), .A2(n2049), .B1(n2048), .B2(n2050), .C1(n2050), 
        .C2(n2049), .ZN(n2044) );
  INV_X1 U1809 ( .A(n610), .ZN(n2050) );
  XNOR2_X1 U1810 ( .A(n1674), .B(n2051), .ZN(n2049) );
  AOI221_X1 U1811 ( .B1(B[16]), .B2(n1558), .C1(B[15]), .C2(n1559), .A(n2052), 
        .ZN(n2051) );
  OAI22_X1 U1812 ( .A1(n1561), .A2(n1640), .B1(n1563), .B2(n1641), .ZN(n2052)
         );
  INV_X1 U1813 ( .A(B[14]), .ZN(n1641) );
  INV_X1 U1814 ( .A(n1382), .ZN(n1640) );
  AOI222_X1 U1815 ( .A1(n2053), .A2(n2054), .B1(n2053), .B2(n620), .C1(n620), 
        .C2(n2054), .ZN(n2048) );
  XNOR2_X1 U1816 ( .A(A[2]), .B(n2055), .ZN(n2054) );
  AOI221_X1 U1817 ( .B1(B[15]), .B2(n1558), .C1(B[14]), .C2(n1559), .A(n2056), 
        .ZN(n2055) );
  OAI22_X1 U1818 ( .A1(n1561), .A2(n1636), .B1(n1563), .B2(n1637), .ZN(n2056)
         );
  INV_X1 U1819 ( .A(B[13]), .ZN(n1637) );
  INV_X1 U1820 ( .A(n1383), .ZN(n1636) );
  OAI222_X1 U1821 ( .A1(n2057), .A2(n2058), .B1(n2057), .B2(n2059), .C1(n2059), 
        .C2(n2058), .ZN(n2053) );
  INV_X1 U1822 ( .A(n630), .ZN(n2059) );
  XNOR2_X1 U1823 ( .A(n1674), .B(n2060), .ZN(n2058) );
  AOI221_X1 U1824 ( .B1(B[14]), .B2(n1558), .C1(B[13]), .C2(n1559), .A(n2061), 
        .ZN(n2060) );
  OAI22_X1 U1825 ( .A1(n1561), .A2(n1632), .B1(n1563), .B2(n1633), .ZN(n2061)
         );
  INV_X1 U1826 ( .A(B[12]), .ZN(n1633) );
  INV_X1 U1827 ( .A(n1384), .ZN(n1632) );
  AOI222_X1 U1828 ( .A1(n2062), .A2(n2063), .B1(n2062), .B2(n638), .C1(n638), 
        .C2(n2063), .ZN(n2057) );
  XNOR2_X1 U1829 ( .A(A[2]), .B(n2064), .ZN(n2063) );
  AOI221_X1 U1830 ( .B1(B[13]), .B2(n1558), .C1(B[12]), .C2(n1559), .A(n2065), 
        .ZN(n2064) );
  OAI22_X1 U1831 ( .A1(n1561), .A2(n1628), .B1(n1563), .B2(n1629), .ZN(n2065)
         );
  INV_X1 U1832 ( .A(B[11]), .ZN(n1629) );
  INV_X1 U1833 ( .A(n1385), .ZN(n1628) );
  OAI222_X1 U1834 ( .A1(n2066), .A2(n2067), .B1(n2066), .B2(n2068), .C1(n2068), 
        .C2(n2067), .ZN(n2062) );
  INV_X1 U1835 ( .A(n646), .ZN(n2068) );
  XNOR2_X1 U1836 ( .A(n1674), .B(n2069), .ZN(n2067) );
  AOI221_X1 U1837 ( .B1(B[12]), .B2(n1558), .C1(B[11]), .C2(n1559), .A(n2070), 
        .ZN(n2069) );
  OAI22_X1 U1838 ( .A1(n1561), .A2(n1624), .B1(n1563), .B2(n1625), .ZN(n2070)
         );
  INV_X1 U1839 ( .A(B[10]), .ZN(n1625) );
  INV_X1 U1840 ( .A(n1386), .ZN(n1624) );
  AOI222_X1 U1841 ( .A1(n2071), .A2(n2072), .B1(n2071), .B2(n654), .C1(n654), 
        .C2(n2072), .ZN(n2066) );
  XNOR2_X1 U1842 ( .A(A[2]), .B(n2073), .ZN(n2072) );
  AOI221_X1 U1843 ( .B1(B[11]), .B2(n1558), .C1(B[10]), .C2(n1559), .A(n2074), 
        .ZN(n2073) );
  OAI22_X1 U1844 ( .A1(n1561), .A2(n1620), .B1(n1563), .B2(n1621), .ZN(n2074)
         );
  INV_X1 U1845 ( .A(B[9]), .ZN(n1621) );
  INV_X1 U1846 ( .A(n1387), .ZN(n1620) );
  OAI222_X1 U1847 ( .A1(n2075), .A2(n2076), .B1(n2075), .B2(n2077), .C1(n2077), 
        .C2(n2076), .ZN(n2071) );
  INV_X1 U1848 ( .A(n660), .ZN(n2077) );
  XNOR2_X1 U1849 ( .A(n1674), .B(n2078), .ZN(n2076) );
  AOI221_X1 U1850 ( .B1(B[10]), .B2(n1558), .C1(B[9]), .C2(n1559), .A(n2079), 
        .ZN(n2078) );
  OAI22_X1 U1851 ( .A1(n1561), .A2(n1616), .B1(n1563), .B2(n1617), .ZN(n2079)
         );
  INV_X1 U1852 ( .A(B[8]), .ZN(n1617) );
  INV_X1 U1853 ( .A(n1388), .ZN(n1616) );
  AOI222_X1 U1854 ( .A1(n2080), .A2(n2081), .B1(n2080), .B2(n666), .C1(n666), 
        .C2(n2081), .ZN(n2075) );
  XNOR2_X1 U1855 ( .A(A[2]), .B(n2082), .ZN(n2081) );
  AOI221_X1 U1856 ( .B1(B[9]), .B2(n1558), .C1(B[8]), .C2(n1559), .A(n2083), 
        .ZN(n2082) );
  OAI22_X1 U1857 ( .A1(n1561), .A2(n1612), .B1(n1563), .B2(n1613), .ZN(n2083)
         );
  INV_X1 U1858 ( .A(B[7]), .ZN(n1613) );
  INV_X1 U1859 ( .A(n1389), .ZN(n1612) );
  OAI222_X1 U1860 ( .A1(n2084), .A2(n2085), .B1(n2084), .B2(n2086), .C1(n2086), 
        .C2(n2085), .ZN(n2080) );
  INV_X1 U1861 ( .A(n672), .ZN(n2086) );
  XNOR2_X1 U1862 ( .A(n1674), .B(n2087), .ZN(n2085) );
  AOI221_X1 U1863 ( .B1(B[8]), .B2(n1558), .C1(B[7]), .C2(n1559), .A(n2088), 
        .ZN(n2087) );
  OAI22_X1 U1864 ( .A1(n1561), .A2(n1608), .B1(n1563), .B2(n1609), .ZN(n2088)
         );
  INV_X1 U1865 ( .A(B[6]), .ZN(n1609) );
  INV_X1 U1866 ( .A(n1390), .ZN(n1608) );
  AOI222_X1 U1867 ( .A1(n2089), .A2(n2090), .B1(n2089), .B2(n676), .C1(n676), 
        .C2(n2090), .ZN(n2084) );
  XNOR2_X1 U1868 ( .A(A[2]), .B(n2091), .ZN(n2090) );
  AOI221_X1 U1869 ( .B1(B[7]), .B2(n1558), .C1(B[6]), .C2(n1559), .A(n2092), 
        .ZN(n2091) );
  OAI22_X1 U1870 ( .A1(n1561), .A2(n1604), .B1(n1563), .B2(n1605), .ZN(n2092)
         );
  INV_X1 U1871 ( .A(B[5]), .ZN(n1605) );
  INV_X1 U1872 ( .A(n1391), .ZN(n1604) );
  OAI222_X1 U1873 ( .A1(n2093), .A2(n2094), .B1(n2093), .B2(n2095), .C1(n2095), 
        .C2(n2094), .ZN(n2089) );
  INV_X1 U1874 ( .A(n680), .ZN(n2095) );
  XNOR2_X1 U1875 ( .A(n1674), .B(n2096), .ZN(n2094) );
  AOI221_X1 U1876 ( .B1(B[6]), .B2(n1558), .C1(B[5]), .C2(n1559), .A(n2097), 
        .ZN(n2096) );
  OAI22_X1 U1877 ( .A1(n1561), .A2(n1600), .B1(n1563), .B2(n1601), .ZN(n2097)
         );
  INV_X1 U1878 ( .A(B[4]), .ZN(n1601) );
  INV_X1 U1879 ( .A(n1392), .ZN(n1600) );
  AOI222_X1 U1880 ( .A1(n2098), .A2(n2099), .B1(n2098), .B2(n684), .C1(n684), 
        .C2(n2099), .ZN(n2093) );
  XNOR2_X1 U1881 ( .A(A[2]), .B(n2100), .ZN(n2099) );
  AOI221_X1 U1882 ( .B1(B[5]), .B2(n1558), .C1(B[4]), .C2(n1559), .A(n2101), 
        .ZN(n2100) );
  OAI22_X1 U1883 ( .A1(n1561), .A2(n1596), .B1(n1563), .B2(n1597), .ZN(n2101)
         );
  INV_X1 U1884 ( .A(B[3]), .ZN(n1597) );
  INV_X1 U1885 ( .A(n1393), .ZN(n1596) );
  OAI222_X1 U1886 ( .A1(n2102), .A2(n2103), .B1(n2102), .B2(n2104), .C1(n2104), 
        .C2(n2103), .ZN(n2098) );
  INV_X1 U1887 ( .A(n686), .ZN(n2104) );
  XNOR2_X1 U1888 ( .A(n1674), .B(n2105), .ZN(n2103) );
  AOI221_X1 U1889 ( .B1(B[4]), .B2(n1558), .C1(B[3]), .C2(n1559), .A(n2106), 
        .ZN(n2105) );
  OAI22_X1 U1890 ( .A1(n1561), .A2(n1592), .B1(n1563), .B2(n1593), .ZN(n2106)
         );
  INV_X1 U1891 ( .A(B[2]), .ZN(n1593) );
  INV_X1 U1892 ( .A(n1394), .ZN(n1592) );
  AOI222_X1 U1893 ( .A1(n2107), .A2(n2108), .B1(n2107), .B2(n688), .C1(n688), 
        .C2(n2108), .ZN(n2102) );
  XNOR2_X1 U1894 ( .A(A[2]), .B(n2109), .ZN(n2108) );
  AOI221_X1 U1895 ( .B1(B[3]), .B2(n1558), .C1(B[2]), .C2(n1559), .A(n2110), 
        .ZN(n2109) );
  OAI22_X1 U1896 ( .A1(n1561), .A2(n1589), .B1(n1563), .B2(n1578), .ZN(n2110)
         );
  INV_X1 U1897 ( .A(B[1]), .ZN(n1578) );
  INV_X1 U1898 ( .A(n1395), .ZN(n1589) );
  AND2_X1 U1899 ( .A1(n2114), .A2(n2115), .ZN(n2107) );
  AOI211_X1 U1900 ( .C1(B[1]), .C2(n1558), .A(n2116), .B(B[0]), .ZN(n2115) );
  INV_X1 U1901 ( .A(n2117), .ZN(n2116) );
  AOI22_X1 U1902 ( .A1(n1558), .A2(B[2]), .B1(n2118), .B2(n1397), .ZN(n2117)
         );
  INV_X1 U1903 ( .A(A[0]), .ZN(n2112) );
  AOI221_X1 U1904 ( .B1(B[1]), .B2(n1559), .C1(n1396), .C2(n2118), .A(n1674), 
        .ZN(n2114) );
  INV_X1 U1905 ( .A(n1561), .ZN(n2118) );
  XNOR2_X1 U1906 ( .A(A[1]), .B(n1674), .ZN(n2111) );
  INV_X1 U1907 ( .A(A[2]), .ZN(n1674) );
  INV_X1 U1908 ( .A(A[1]), .ZN(n2113) );
  AOI21_X1 U1909 ( .B1(n2119), .B2(n2120), .A(n2121), .ZN(PRODUCT[47]) );
  OAI22_X1 U1910 ( .A1(n2122), .A2(n2123), .B1(n2122), .B2(n2124), .ZN(n2121)
         );
  INV_X1 U1911 ( .A(n2120), .ZN(n2124) );
  AOI222_X1 U1912 ( .A1(n2024), .A2(n303), .B1(n2123), .B2(n303), .C1(n2024), 
        .C2(n2123), .ZN(n2122) );
  XOR2_X1 U1913 ( .A(n1541), .B(n2125), .Z(n2024) );
  AOI221_X1 U1914 ( .B1(n1537), .B2(B[23]), .C1(n1536), .C2(B[22]), .A(n2126), 
        .ZN(n2125) );
  OAI22_X1 U1915 ( .A1(n1567), .A2(n1976), .B1(n1568), .B2(n1538), .ZN(n2126)
         );
  INV_X1 U1916 ( .A(B[21]), .ZN(n1568) );
  INV_X1 U1917 ( .A(n1375), .ZN(n1567) );
  XOR2_X1 U1918 ( .A(n2127), .B(n1541), .Z(n2120) );
  OAI221_X1 U1919 ( .B1(n1556), .B2(n1539), .C1(n1556), .C2(n1976), .A(n2128), 
        .ZN(n2127) );
  OAI21_X1 U1920 ( .B1(n1537), .B2(n1536), .A(n1554), .ZN(n2128) );
  INV_X1 U1921 ( .A(n2123), .ZN(n2119) );
  XOR2_X1 U1922 ( .A(A[23]), .B(n2129), .Z(n2123) );
  AOI221_X1 U1923 ( .B1(n1537), .B2(n1554), .C1(n1536), .C2(n1554), .A(n2130), 
        .ZN(n2129) );
  OAI22_X1 U1924 ( .A1(n1571), .A2(n1976), .B1(n1572), .B2(n1538), .ZN(n2130)
         );
  NAND3_X1 U1925 ( .A1(n2131), .A2(n2132), .A3(n2133), .ZN(n1980) );
  INV_X1 U1926 ( .A(B[22]), .ZN(n1572) );
  INV_X1 U1927 ( .A(n1374), .ZN(n1571) );
  XNOR2_X1 U1928 ( .A(A[21]), .B(A[22]), .ZN(n2133) );
  INV_X1 U1929 ( .A(n2131), .ZN(n2134) );
  XOR2_X1 U1930 ( .A(A[21]), .B(n1543), .Z(n2131) );
  XNOR2_X1 U1931 ( .A(A[22]), .B(n1541), .ZN(n2132) );
endmodule


module iir_filter_DW02_mult_4 ( A, B, PRODUCT, TC );
  input [23:0] A;
  input [23:0] B;
  output [47:0] PRODUCT;
  input TC;
  wire   n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n351, n352, n353, n354, n355, n356, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n906, n907, n908, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134;

  FA_X1 U182 ( .A(n351), .B(n352), .CI(n304), .CO(n303), .S(PRODUCT[44]) );
  FA_X1 U183 ( .A(n353), .B(n354), .CI(n305), .CO(n304), .S(PRODUCT[43]) );
  FA_X1 U184 ( .A(n355), .B(n358), .CI(n306), .CO(n305), .S(PRODUCT[42]) );
  FA_X1 U185 ( .A(n359), .B(n361), .CI(n307), .CO(n306), .S(PRODUCT[41]) );
  FA_X1 U186 ( .A(n362), .B(n364), .CI(n308), .CO(n307), .S(PRODUCT[40]) );
  FA_X1 U187 ( .A(n365), .B(n370), .CI(n309), .CO(n308), .S(PRODUCT[39]) );
  FA_X1 U188 ( .A(n371), .B(n375), .CI(n310), .CO(n309), .S(PRODUCT[38]) );
  FA_X1 U189 ( .A(n376), .B(n381), .CI(n311), .CO(n310), .S(PRODUCT[37]) );
  FA_X1 U190 ( .A(n382), .B(n389), .CI(n312), .CO(n311), .S(PRODUCT[36]) );
  FA_X1 U191 ( .A(n390), .B(n396), .CI(n313), .CO(n312), .S(PRODUCT[35]) );
  FA_X1 U192 ( .A(n397), .B(n403), .CI(n314), .CO(n313), .S(PRODUCT[34]) );
  FA_X1 U193 ( .A(n404), .B(n413), .CI(n315), .CO(n314), .S(PRODUCT[33]) );
  FA_X1 U194 ( .A(n414), .B(n422), .CI(n316), .CO(n315), .S(PRODUCT[32]) );
  FA_X1 U195 ( .A(n423), .B(n432), .CI(n317), .CO(n316), .S(PRODUCT[31]) );
  FA_X1 U196 ( .A(n433), .B(n444), .CI(n318), .CO(n317), .S(PRODUCT[30]) );
  FA_X1 U197 ( .A(n445), .B(n455), .CI(n319), .CO(n318), .S(PRODUCT[29]) );
  FA_X1 U198 ( .A(n456), .B(n467), .CI(n320), .CO(n319), .S(PRODUCT[28]) );
  FA_X1 U199 ( .A(n468), .B(n481), .CI(n321), .CO(n320), .S(PRODUCT[27]) );
  FA_X1 U200 ( .A(n482), .B(n494), .CI(n322), .CO(n321), .S(PRODUCT[26]) );
  FA_X1 U201 ( .A(n495), .B(n507), .CI(n323), .CO(n322), .S(PRODUCT[25]) );
  FA_X1 U202 ( .A(n508), .B(n906), .CI(n324), .CO(n323), .S(PRODUCT[24]) );
  FA_X1 U203 ( .A(n907), .B(n522), .CI(n325), .CO(n324), .S(PRODUCT[23]) );
  FA_X1 U204 ( .A(n908), .B(n536), .CI(n326), .CO(n325), .S(PRODUCT[22]) );
  FA_X1 U235 ( .A(n356), .B(n749), .CI(n729), .CO(n352), .S(n353) );
  FA_X1 U236 ( .A(n730), .B(n360), .CI(n750), .CO(n354), .S(n355) );
  FA_X1 U238 ( .A(n360), .B(n731), .CI(n751), .CO(n358), .S(n359) );
  FA_X1 U240 ( .A(n752), .B(n363), .CI(n366), .CO(n361), .S(n362) );
  FA_X1 U241 ( .A(n368), .B(n775), .CI(n732), .CO(n356), .S(n363) );
  FA_X1 U242 ( .A(n776), .B(n753), .CI(n367), .CO(n364), .S(n365) );
  FA_X1 U243 ( .A(n733), .B(n374), .CI(n372), .CO(n366), .S(n367) );
  FA_X1 U245 ( .A(n373), .B(n377), .CI(n777), .CO(n370), .S(n371) );
  FA_X1 U246 ( .A(n374), .B(n379), .CI(n754), .CO(n372), .S(n373) );
  FA_X1 U248 ( .A(n778), .B(n378), .CI(n383), .CO(n375), .S(n376) );
  FA_X1 U249 ( .A(n385), .B(n380), .CI(n755), .CO(n377), .S(n378) );
  FA_X1 U250 ( .A(n387), .B(n801), .CI(n734), .CO(n379), .S(n380) );
  FA_X1 U251 ( .A(n802), .B(n779), .CI(n384), .CO(n381), .S(n382) );
  FA_X1 U252 ( .A(n386), .B(n393), .CI(n391), .CO(n383), .S(n384) );
  FA_X1 U253 ( .A(n735), .B(n395), .CI(n756), .CO(n385), .S(n386) );
  FA_X1 U255 ( .A(n392), .B(n398), .CI(n803), .CO(n389), .S(n390) );
  FA_X1 U256 ( .A(n394), .B(n400), .CI(n780), .CO(n391), .S(n392) );
  FA_X1 U257 ( .A(n395), .B(n736), .CI(n757), .CO(n393), .S(n394) );
  FA_X1 U259 ( .A(n804), .B(n399), .CI(n405), .CO(n396), .S(n397) );
  FA_X1 U260 ( .A(n407), .B(n401), .CI(n781), .CO(n398), .S(n399) );
  FA_X1 U261 ( .A(n758), .B(n402), .CI(n409), .CO(n400), .S(n401) );
  FA_X1 U262 ( .A(n411), .B(n827), .CI(n737), .CO(n387), .S(n402) );
  FA_X1 U263 ( .A(n828), .B(n805), .CI(n406), .CO(n403), .S(n404) );
  FA_X1 U264 ( .A(n408), .B(n417), .CI(n415), .CO(n405), .S(n406) );
  FA_X1 U265 ( .A(n410), .B(n759), .CI(n782), .CO(n407), .S(n408) );
  FA_X1 U266 ( .A(n738), .B(n421), .CI(n419), .CO(n409), .S(n410) );
  FA_X1 U268 ( .A(n416), .B(n424), .CI(n829), .CO(n413), .S(n414) );
  FA_X1 U269 ( .A(n418), .B(n426), .CI(n806), .CO(n415), .S(n416) );
  FA_X1 U270 ( .A(n420), .B(n428), .CI(n783), .CO(n417), .S(n418) );
  FA_X1 U271 ( .A(n421), .B(n430), .CI(n760), .CO(n419), .S(n420) );
  FA_X1 U273 ( .A(n830), .B(n425), .CI(n434), .CO(n422), .S(n423) );
  FA_X1 U274 ( .A(n436), .B(n427), .CI(n807), .CO(n424), .S(n425) );
  FA_X1 U275 ( .A(n784), .B(n429), .CI(n438), .CO(n426), .S(n427) );
  FA_X1 U276 ( .A(n440), .B(n431), .CI(n761), .CO(n428), .S(n429) );
  FA_X1 U277 ( .A(n442), .B(n853), .CI(n739), .CO(n430), .S(n431) );
  FA_X1 U278 ( .A(n854), .B(n831), .CI(n435), .CO(n432), .S(n433) );
  FA_X1 U279 ( .A(n437), .B(n448), .CI(n446), .CO(n434), .S(n435) );
  FA_X1 U280 ( .A(n439), .B(n785), .CI(n808), .CO(n436), .S(n437) );
  FA_X1 U281 ( .A(n441), .B(n452), .CI(n450), .CO(n438), .S(n439) );
  FA_X1 U282 ( .A(n740), .B(n454), .CI(n762), .CO(n440), .S(n441) );
  FA_X1 U284 ( .A(n447), .B(n457), .CI(n855), .CO(n444), .S(n445) );
  FA_X1 U285 ( .A(n449), .B(n459), .CI(n832), .CO(n446), .S(n447) );
  FA_X1 U286 ( .A(n451), .B(n461), .CI(n809), .CO(n448), .S(n449) );
  FA_X1 U287 ( .A(n453), .B(n463), .CI(n786), .CO(n450), .S(n451) );
  FA_X1 U288 ( .A(n454), .B(n465), .CI(n763), .CO(n452), .S(n453) );
  FA_X1 U290 ( .A(n856), .B(n458), .CI(n469), .CO(n455), .S(n456) );
  FA_X1 U291 ( .A(n471), .B(n460), .CI(n833), .CO(n457), .S(n458) );
  FA_X1 U292 ( .A(n810), .B(n462), .CI(n473), .CO(n459), .S(n460) );
  FA_X1 U293 ( .A(n475), .B(n464), .CI(n787), .CO(n461), .S(n462) );
  FA_X1 U294 ( .A(n764), .B(n466), .CI(n477), .CO(n463), .S(n464) );
  FA_X1 U295 ( .A(n479), .B(n879), .CI(n741), .CO(n465), .S(n466) );
  FA_X1 U296 ( .A(n880), .B(n857), .CI(n470), .CO(n467), .S(n468) );
  FA_X1 U297 ( .A(n472), .B(n485), .CI(n483), .CO(n469), .S(n470) );
  FA_X1 U298 ( .A(n474), .B(n811), .CI(n834), .CO(n471), .S(n472) );
  FA_X1 U299 ( .A(n476), .B(n489), .CI(n487), .CO(n473), .S(n474) );
  FA_X1 U300 ( .A(n478), .B(n765), .CI(n788), .CO(n475), .S(n476) );
  FA_X1 U301 ( .A(n742), .B(n493), .CI(n491), .CO(n477), .S(n478) );
  FA_X1 U303 ( .A(n484), .B(n858), .CI(n881), .CO(n481), .S(n482) );
  FA_X1 U304 ( .A(n486), .B(n498), .CI(n496), .CO(n483), .S(n484) );
  FA_X1 U305 ( .A(n488), .B(n812), .CI(n835), .CO(n485), .S(n486) );
  FA_X1 U306 ( .A(n490), .B(n502), .CI(n500), .CO(n487), .S(n488) );
  FA_X1 U307 ( .A(n492), .B(n504), .CI(n789), .CO(n489), .S(n490) );
  FA_X1 U308 ( .A(n743), .B(n493), .CI(n766), .CO(n491), .S(n492) );
  FA_X1 U310 ( .A(n497), .B(n509), .CI(n882), .CO(n494), .S(n495) );
  FA_X1 U311 ( .A(n499), .B(n511), .CI(n859), .CO(n496), .S(n497) );
  FA_X1 U312 ( .A(n501), .B(n513), .CI(n836), .CO(n498), .S(n499) );
  FA_X1 U313 ( .A(n503), .B(n515), .CI(n813), .CO(n500), .S(n501) );
  FA_X1 U314 ( .A(n505), .B(n517), .CI(n790), .CO(n502), .S(n503) );
  FA_X1 U315 ( .A(n506), .B(n744), .CI(n767), .CO(n504), .S(n505) );
  FA_X1 U318 ( .A(n883), .B(n510), .CI(n521), .CO(n507), .S(n508) );
  FA_X1 U319 ( .A(n860), .B(n512), .CI(n523), .CO(n509), .S(n510) );
  FA_X1 U320 ( .A(n837), .B(n514), .CI(n525), .CO(n511), .S(n512) );
  FA_X1 U321 ( .A(n814), .B(n516), .CI(n527), .CO(n513), .S(n514) );
  FA_X1 U322 ( .A(n791), .B(n518), .CI(n529), .CO(n515), .S(n516) );
  FA_X1 U323 ( .A(n768), .B(n520), .CI(n531), .CO(n517), .S(n518) );
  HA_X1 U324 ( .A(n533), .B(n745), .CO(n519), .S(n520) );
  FA_X1 U325 ( .A(n884), .B(n524), .CI(n535), .CO(n521), .S(n522) );
  FA_X1 U326 ( .A(n861), .B(n526), .CI(n537), .CO(n523), .S(n524) );
  FA_X1 U327 ( .A(n838), .B(n528), .CI(n539), .CO(n525), .S(n526) );
  FA_X1 U328 ( .A(n815), .B(n530), .CI(n541), .CO(n527), .S(n528) );
  FA_X1 U329 ( .A(n792), .B(n532), .CI(n543), .CO(n529), .S(n530) );
  FA_X1 U330 ( .A(n769), .B(n534), .CI(n545), .CO(n531), .S(n532) );
  HA_X1 U331 ( .A(n547), .B(n746), .CO(n533), .S(n534) );
  FA_X1 U332 ( .A(n885), .B(n538), .CI(n549), .CO(n535), .S(n536) );
  FA_X1 U333 ( .A(n862), .B(n540), .CI(n551), .CO(n537), .S(n538) );
  FA_X1 U334 ( .A(n839), .B(n542), .CI(n553), .CO(n539), .S(n540) );
  FA_X1 U335 ( .A(n816), .B(n544), .CI(n555), .CO(n541), .S(n542) );
  FA_X1 U336 ( .A(n793), .B(n546), .CI(n557), .CO(n543), .S(n544) );
  FA_X1 U337 ( .A(n770), .B(n548), .CI(n559), .CO(n545), .S(n546) );
  HA_X1 U338 ( .A(n561), .B(n747), .CO(n547), .S(n548) );
  FA_X1 U339 ( .A(n886), .B(n552), .CI(n563), .CO(n549), .S(n550) );
  FA_X1 U340 ( .A(n863), .B(n554), .CI(n565), .CO(n551), .S(n552) );
  FA_X1 U341 ( .A(n840), .B(n556), .CI(n567), .CO(n553), .S(n554) );
  FA_X1 U342 ( .A(n817), .B(n558), .CI(n569), .CO(n555), .S(n556) );
  FA_X1 U343 ( .A(n794), .B(n560), .CI(n571), .CO(n557), .S(n558) );
  FA_X1 U344 ( .A(n771), .B(n562), .CI(n573), .CO(n559), .S(n560) );
  HA_X1 U345 ( .A(n748), .B(n1540), .CO(n561), .S(n562) );
  FA_X1 U346 ( .A(n887), .B(n566), .CI(n575), .CO(n563), .S(n564) );
  FA_X1 U347 ( .A(n864), .B(n568), .CI(n577), .CO(n565), .S(n566) );
  FA_X1 U348 ( .A(n841), .B(n570), .CI(n579), .CO(n567), .S(n568) );
  FA_X1 U349 ( .A(n818), .B(n572), .CI(n581), .CO(n569), .S(n570) );
  FA_X1 U350 ( .A(n795), .B(n574), .CI(n583), .CO(n571), .S(n572) );
  HA_X1 U351 ( .A(n585), .B(n772), .CO(n573), .S(n574) );
  FA_X1 U352 ( .A(n888), .B(n578), .CI(n587), .CO(n575), .S(n576) );
  FA_X1 U353 ( .A(n865), .B(n580), .CI(n589), .CO(n577), .S(n578) );
  FA_X1 U354 ( .A(n842), .B(n582), .CI(n591), .CO(n579), .S(n580) );
  FA_X1 U355 ( .A(n819), .B(n584), .CI(n593), .CO(n581), .S(n582) );
  FA_X1 U356 ( .A(n796), .B(n586), .CI(n595), .CO(n583), .S(n584) );
  HA_X1 U357 ( .A(n597), .B(n773), .CO(n585), .S(n586) );
  FA_X1 U358 ( .A(n889), .B(n590), .CI(n599), .CO(n587), .S(n588) );
  FA_X1 U359 ( .A(n866), .B(n592), .CI(n601), .CO(n589), .S(n590) );
  FA_X1 U360 ( .A(n843), .B(n594), .CI(n603), .CO(n591), .S(n592) );
  FA_X1 U361 ( .A(n820), .B(n596), .CI(n605), .CO(n593), .S(n594) );
  FA_X1 U362 ( .A(n797), .B(n598), .CI(n607), .CO(n595), .S(n596) );
  HA_X1 U363 ( .A(n774), .B(n1542), .CO(n597), .S(n598) );
  FA_X1 U364 ( .A(n890), .B(n602), .CI(n609), .CO(n599), .S(n600) );
  FA_X1 U365 ( .A(n867), .B(n604), .CI(n611), .CO(n601), .S(n602) );
  FA_X1 U366 ( .A(n844), .B(n606), .CI(n613), .CO(n603), .S(n604) );
  FA_X1 U367 ( .A(n821), .B(n608), .CI(n615), .CO(n605), .S(n606) );
  HA_X1 U368 ( .A(n617), .B(n798), .CO(n607), .S(n608) );
  FA_X1 U369 ( .A(n891), .B(n612), .CI(n619), .CO(n609), .S(n610) );
  FA_X1 U370 ( .A(n868), .B(n614), .CI(n621), .CO(n611), .S(n612) );
  FA_X1 U371 ( .A(n845), .B(n616), .CI(n623), .CO(n613), .S(n614) );
  FA_X1 U372 ( .A(n822), .B(n618), .CI(n625), .CO(n615), .S(n616) );
  HA_X1 U373 ( .A(n627), .B(n799), .CO(n617), .S(n618) );
  FA_X1 U374 ( .A(n892), .B(n622), .CI(n629), .CO(n619), .S(n620) );
  FA_X1 U375 ( .A(n869), .B(n624), .CI(n631), .CO(n621), .S(n622) );
  FA_X1 U376 ( .A(n846), .B(n626), .CI(n633), .CO(n623), .S(n624) );
  FA_X1 U377 ( .A(n823), .B(n628), .CI(n635), .CO(n625), .S(n626) );
  HA_X1 U378 ( .A(n800), .B(n1544), .CO(n627), .S(n628) );
  FA_X1 U379 ( .A(n893), .B(n632), .CI(n637), .CO(n629), .S(n630) );
  FA_X1 U380 ( .A(n870), .B(n634), .CI(n639), .CO(n631), .S(n632) );
  FA_X1 U381 ( .A(n847), .B(n636), .CI(n641), .CO(n633), .S(n634) );
  HA_X1 U382 ( .A(n643), .B(n824), .CO(n635), .S(n636) );
  FA_X1 U383 ( .A(n894), .B(n640), .CI(n645), .CO(n637), .S(n638) );
  FA_X1 U384 ( .A(n871), .B(n642), .CI(n647), .CO(n639), .S(n640) );
  FA_X1 U385 ( .A(n848), .B(n644), .CI(n649), .CO(n641), .S(n642) );
  HA_X1 U386 ( .A(n651), .B(n825), .CO(n643), .S(n644) );
  FA_X1 U387 ( .A(n895), .B(n648), .CI(n653), .CO(n645), .S(n646) );
  FA_X1 U388 ( .A(n872), .B(n650), .CI(n655), .CO(n647), .S(n648) );
  FA_X1 U389 ( .A(n849), .B(n652), .CI(n657), .CO(n649), .S(n650) );
  HA_X1 U390 ( .A(n826), .B(n1546), .CO(n651), .S(n652) );
  FA_X1 U391 ( .A(n896), .B(n656), .CI(n659), .CO(n653), .S(n654) );
  FA_X1 U392 ( .A(n873), .B(n658), .CI(n661), .CO(n655), .S(n656) );
  HA_X1 U393 ( .A(n663), .B(n850), .CO(n657), .S(n658) );
  FA_X1 U394 ( .A(n897), .B(n662), .CI(n665), .CO(n659), .S(n660) );
  FA_X1 U395 ( .A(n874), .B(n664), .CI(n667), .CO(n661), .S(n662) );
  HA_X1 U396 ( .A(n669), .B(n851), .CO(n663), .S(n664) );
  FA_X1 U397 ( .A(n898), .B(n668), .CI(n671), .CO(n665), .S(n666) );
  FA_X1 U398 ( .A(n875), .B(n670), .CI(n673), .CO(n667), .S(n668) );
  HA_X1 U399 ( .A(n852), .B(n1548), .CO(n669), .S(n670) );
  FA_X1 U400 ( .A(n899), .B(n674), .CI(n675), .CO(n671), .S(n672) );
  HA_X1 U401 ( .A(n677), .B(n876), .CO(n673), .S(n674) );
  FA_X1 U402 ( .A(n900), .B(n678), .CI(n679), .CO(n675), .S(n676) );
  HA_X1 U403 ( .A(n681), .B(n877), .CO(n677), .S(n678) );
  FA_X1 U404 ( .A(n901), .B(n682), .CI(n683), .CO(n679), .S(n680) );
  HA_X1 U405 ( .A(n878), .B(n1550), .CO(n681), .S(n682) );
  HA_X1 U406 ( .A(n685), .B(n902), .CO(n683), .S(n684) );
  HA_X1 U407 ( .A(n687), .B(n903), .CO(n685), .S(n686) );
  HA_X1 U408 ( .A(n904), .B(n1552), .CO(n687), .S(n688) );
  FA_X1 U1112 ( .A(B[22]), .B(n1554), .CI(n706), .CO(n1374), .S(n1375) );
  FA_X1 U1113 ( .A(B[21]), .B(B[22]), .CI(n707), .CO(n706), .S(n1376) );
  FA_X1 U1114 ( .A(B[20]), .B(B[21]), .CI(n708), .CO(n707), .S(n1377) );
  FA_X1 U1115 ( .A(B[19]), .B(B[20]), .CI(n709), .CO(n708), .S(n1378) );
  FA_X1 U1116 ( .A(B[18]), .B(B[19]), .CI(n710), .CO(n709), .S(n1379) );
  FA_X1 U1117 ( .A(B[17]), .B(B[18]), .CI(n711), .CO(n710), .S(n1380) );
  FA_X1 U1118 ( .A(B[16]), .B(B[17]), .CI(n712), .CO(n711), .S(n1381) );
  FA_X1 U1119 ( .A(B[15]), .B(B[16]), .CI(n713), .CO(n712), .S(n1382) );
  FA_X1 U1120 ( .A(B[14]), .B(B[15]), .CI(n714), .CO(n713), .S(n1383) );
  FA_X1 U1121 ( .A(B[13]), .B(B[14]), .CI(n715), .CO(n714), .S(n1384) );
  FA_X1 U1122 ( .A(B[12]), .B(B[13]), .CI(n716), .CO(n715), .S(n1385) );
  FA_X1 U1123 ( .A(B[11]), .B(B[12]), .CI(n717), .CO(n716), .S(n1386) );
  FA_X1 U1124 ( .A(B[10]), .B(B[11]), .CI(n718), .CO(n717), .S(n1387) );
  FA_X1 U1125 ( .A(B[9]), .B(B[10]), .CI(n719), .CO(n718), .S(n1388) );
  FA_X1 U1126 ( .A(B[8]), .B(B[9]), .CI(n720), .CO(n719), .S(n1389) );
  FA_X1 U1127 ( .A(B[7]), .B(B[8]), .CI(n721), .CO(n720), .S(n1390) );
  FA_X1 U1128 ( .A(B[6]), .B(B[7]), .CI(n722), .CO(n721), .S(n1391) );
  FA_X1 U1129 ( .A(B[5]), .B(B[6]), .CI(n723), .CO(n722), .S(n1392) );
  FA_X1 U1130 ( .A(B[4]), .B(B[5]), .CI(n724), .CO(n723), .S(n1393) );
  FA_X1 U1131 ( .A(B[3]), .B(B[4]), .CI(n725), .CO(n724), .S(n1394) );
  FA_X1 U1132 ( .A(B[2]), .B(B[3]), .CI(n726), .CO(n725), .S(n1395) );
  FA_X1 U1133 ( .A(B[1]), .B(B[2]), .CI(n727), .CO(n726), .S(n1396) );
  HA_X1 U1134 ( .A(B[0]), .B(B[1]), .CO(n727), .S(n1397) );
  OR2_X1 U1138 ( .A1(n2134), .A2(n2133), .ZN(n1534) );
  INV_X1 U1139 ( .A(n1555), .ZN(n1554) );
  INV_X1 U1140 ( .A(n1534), .ZN(n1536) );
  INV_X1 U1141 ( .A(n1535), .ZN(n1537) );
  BUF_X1 U1142 ( .A(n1980), .Z(n1538) );
  BUF_X1 U1143 ( .A(n1980), .Z(n1539) );
  NAND3_X1 U1144 ( .A1(n1673), .A2(n1672), .A3(n1671), .ZN(n1586) );
  NAND3_X1 U1145 ( .A1(n1854), .A2(n1853), .A3(n1852), .ZN(n1804) );
  NAND3_X1 U1146 ( .A1(n1794), .A2(n1793), .A3(n1792), .ZN(n1744) );
  NAND3_X1 U1147 ( .A1(n1734), .A2(n1733), .A3(n1732), .ZN(n1684) );
  NAND3_X1 U1148 ( .A1(n2111), .A2(n2112), .A3(n2113), .ZN(n1563) );
  NAND2_X1 U1149 ( .A1(n1911), .A2(n1913), .ZN(n1857) );
  NAND2_X1 U1150 ( .A1(n1851), .A2(n1853), .ZN(n1797) );
  NAND2_X1 U1151 ( .A1(n1791), .A2(n1793), .ZN(n1737) );
  NAND2_X1 U1152 ( .A1(n1731), .A2(n1733), .ZN(n1677) );
  INV_X1 U1153 ( .A(n1553), .ZN(n1552) );
  INV_X1 U1154 ( .A(n1549), .ZN(n1548) );
  INV_X1 U1155 ( .A(n1551), .ZN(n1550) );
  NAND3_X1 U1156 ( .A1(n1914), .A2(n1913), .A3(n1912), .ZN(n1864) );
  NAND3_X1 U1157 ( .A1(n1974), .A2(n1973), .A3(n1972), .ZN(n1924) );
  NAND2_X1 U1158 ( .A1(n2134), .A2(n2132), .ZN(n1976) );
  NAND2_X1 U1159 ( .A1(n1971), .A2(n1973), .ZN(n1917) );
  INV_X1 U1160 ( .A(n1547), .ZN(n1546) );
  INV_X1 U1161 ( .A(n1541), .ZN(n1540) );
  INV_X1 U1162 ( .A(n1543), .ZN(n1542) );
  INV_X1 U1163 ( .A(n1545), .ZN(n1544) );
  OR2_X1 U1164 ( .A1(n2132), .A2(n2131), .ZN(n1535) );
  NAND2_X1 U1165 ( .A1(A[0]), .A2(n2111), .ZN(n1561) );
  INV_X1 U1166 ( .A(A[5]), .ZN(n1553) );
  INV_X1 U1167 ( .A(A[11]), .ZN(n1549) );
  INV_X1 U1168 ( .A(A[8]), .ZN(n1551) );
  INV_X1 U1169 ( .A(A[14]), .ZN(n1547) );
  INV_X1 U1170 ( .A(A[17]), .ZN(n1545) );
  INV_X1 U1171 ( .A(A[23]), .ZN(n1541) );
  INV_X1 U1172 ( .A(A[20]), .ZN(n1543) );
  NOR2_X4 U1173 ( .A1(n1670), .A2(n1671), .ZN(n1581) );
  NOR2_X4 U1174 ( .A1(n1672), .A2(n1673), .ZN(n1582) );
  NAND2_X2 U1175 ( .A1(n1670), .A2(n1672), .ZN(n1576) );
  NOR2_X4 U1176 ( .A1(n1731), .A2(n1732), .ZN(n1680) );
  NOR2_X4 U1177 ( .A1(n1733), .A2(n1734), .ZN(n1681) );
  NOR2_X4 U1178 ( .A1(n1791), .A2(n1792), .ZN(n1740) );
  NOR2_X4 U1179 ( .A1(n1793), .A2(n1794), .ZN(n1741) );
  NOR2_X4 U1180 ( .A1(n1851), .A2(n1852), .ZN(n1800) );
  NOR2_X4 U1181 ( .A1(n1853), .A2(n1854), .ZN(n1801) );
  NOR2_X4 U1182 ( .A1(n1911), .A2(n1912), .ZN(n1860) );
  NOR2_X4 U1183 ( .A1(n1913), .A2(n1914), .ZN(n1861) );
  NOR2_X4 U1184 ( .A1(n1971), .A2(n1972), .ZN(n1920) );
  NOR2_X4 U1185 ( .A1(n1973), .A2(n1974), .ZN(n1921) );
  INV_X2 U1186 ( .A(B[0]), .ZN(n1574) );
  NOR2_X4 U1187 ( .A1(n2112), .A2(n2111), .ZN(n1558) );
  NOR2_X4 U1188 ( .A1(n2113), .A2(A[0]), .ZN(n1559) );
  INV_X1 U1189 ( .A(B[23]), .ZN(n1555) );
  INV_X1 U1190 ( .A(B[23]), .ZN(n1556) );
  XNOR2_X1 U1191 ( .A(A[2]), .B(n1557), .ZN(n908) );
  AOI221_X1 U1192 ( .B1(B[22]), .B2(n1558), .C1(B[21]), .C2(n1559), .A(n1560), 
        .ZN(n1557) );
  OAI22_X1 U1193 ( .A1(n1561), .A2(n1562), .B1(n1563), .B2(n1564), .ZN(n1560)
         );
  XNOR2_X1 U1194 ( .A(A[2]), .B(n1565), .ZN(n907) );
  AOI221_X1 U1195 ( .B1(B[23]), .B2(n1558), .C1(n1559), .C2(B[22]), .A(n1566), 
        .ZN(n1565) );
  OAI22_X1 U1196 ( .A1(n1561), .A2(n1567), .B1(n1568), .B2(n1563), .ZN(n1566)
         );
  XNOR2_X1 U1197 ( .A(A[2]), .B(n1569), .ZN(n906) );
  AOI221_X1 U1198 ( .B1(B[23]), .B2(n1558), .C1(n1554), .C2(n1559), .A(n1570), 
        .ZN(n1569) );
  OAI22_X1 U1199 ( .A1(n1561), .A2(n1571), .B1(n1572), .B2(n1563), .ZN(n1570)
         );
  XNOR2_X1 U1200 ( .A(n1573), .B(n1553), .ZN(n904) );
  OAI22_X1 U1201 ( .A1(n1574), .A2(n1575), .B1(n1576), .B2(n1574), .ZN(n1573)
         );
  XNOR2_X1 U1202 ( .A(n1577), .B(n1553), .ZN(n903) );
  OAI222_X1 U1203 ( .A1(n1575), .A2(n1578), .B1(n1574), .B2(n1579), .C1(n1576), 
        .C2(n1580), .ZN(n1577) );
  INV_X1 U1204 ( .A(n1581), .ZN(n1579) );
  INV_X1 U1205 ( .A(n1582), .ZN(n1575) );
  XNOR2_X1 U1206 ( .A(n1552), .B(n1583), .ZN(n902) );
  AOI221_X1 U1207 ( .B1(B[2]), .B2(n1582), .C1(B[1]), .C2(n1581), .A(n1584), 
        .ZN(n1583) );
  OAI22_X1 U1208 ( .A1(n1576), .A2(n1585), .B1(n1574), .B2(n1586), .ZN(n1584)
         );
  XNOR2_X1 U1209 ( .A(n1552), .B(n1587), .ZN(n901) );
  AOI221_X1 U1210 ( .B1(B[3]), .B2(n1582), .C1(B[2]), .C2(n1581), .A(n1588), 
        .ZN(n1587) );
  OAI22_X1 U1211 ( .A1(n1576), .A2(n1589), .B1(n1578), .B2(n1586), .ZN(n1588)
         );
  XNOR2_X1 U1212 ( .A(n1552), .B(n1590), .ZN(n900) );
  AOI221_X1 U1213 ( .B1(B[4]), .B2(n1582), .C1(B[3]), .C2(n1581), .A(n1591), 
        .ZN(n1590) );
  OAI22_X1 U1214 ( .A1(n1576), .A2(n1592), .B1(n1593), .B2(n1586), .ZN(n1591)
         );
  XNOR2_X1 U1215 ( .A(n1552), .B(n1594), .ZN(n899) );
  AOI221_X1 U1216 ( .B1(B[5]), .B2(n1582), .C1(B[4]), .C2(n1581), .A(n1595), 
        .ZN(n1594) );
  OAI22_X1 U1217 ( .A1(n1576), .A2(n1596), .B1(n1586), .B2(n1597), .ZN(n1595)
         );
  XNOR2_X1 U1218 ( .A(n1552), .B(n1598), .ZN(n898) );
  AOI221_X1 U1219 ( .B1(B[6]), .B2(n1582), .C1(B[5]), .C2(n1581), .A(n1599), 
        .ZN(n1598) );
  OAI22_X1 U1220 ( .A1(n1576), .A2(n1600), .B1(n1586), .B2(n1601), .ZN(n1599)
         );
  XNOR2_X1 U1221 ( .A(n1552), .B(n1602), .ZN(n897) );
  AOI221_X1 U1222 ( .B1(B[7]), .B2(n1582), .C1(B[6]), .C2(n1581), .A(n1603), 
        .ZN(n1602) );
  OAI22_X1 U1223 ( .A1(n1576), .A2(n1604), .B1(n1586), .B2(n1605), .ZN(n1603)
         );
  XNOR2_X1 U1224 ( .A(n1552), .B(n1606), .ZN(n896) );
  AOI221_X1 U1225 ( .B1(B[8]), .B2(n1582), .C1(B[7]), .C2(n1581), .A(n1607), 
        .ZN(n1606) );
  OAI22_X1 U1226 ( .A1(n1576), .A2(n1608), .B1(n1586), .B2(n1609), .ZN(n1607)
         );
  XNOR2_X1 U1227 ( .A(n1552), .B(n1610), .ZN(n895) );
  AOI221_X1 U1228 ( .B1(B[9]), .B2(n1582), .C1(B[8]), .C2(n1581), .A(n1611), 
        .ZN(n1610) );
  OAI22_X1 U1229 ( .A1(n1576), .A2(n1612), .B1(n1586), .B2(n1613), .ZN(n1611)
         );
  XNOR2_X1 U1230 ( .A(n1552), .B(n1614), .ZN(n894) );
  AOI221_X1 U1231 ( .B1(B[10]), .B2(n1582), .C1(B[9]), .C2(n1581), .A(n1615), 
        .ZN(n1614) );
  OAI22_X1 U1232 ( .A1(n1576), .A2(n1616), .B1(n1586), .B2(n1617), .ZN(n1615)
         );
  XNOR2_X1 U1233 ( .A(n1552), .B(n1618), .ZN(n893) );
  AOI221_X1 U1234 ( .B1(B[11]), .B2(n1582), .C1(B[10]), .C2(n1581), .A(n1619), 
        .ZN(n1618) );
  OAI22_X1 U1235 ( .A1(n1576), .A2(n1620), .B1(n1586), .B2(n1621), .ZN(n1619)
         );
  XNOR2_X1 U1236 ( .A(n1552), .B(n1622), .ZN(n892) );
  AOI221_X1 U1237 ( .B1(B[12]), .B2(n1582), .C1(B[11]), .C2(n1581), .A(n1623), 
        .ZN(n1622) );
  OAI22_X1 U1238 ( .A1(n1576), .A2(n1624), .B1(n1586), .B2(n1625), .ZN(n1623)
         );
  XNOR2_X1 U1239 ( .A(n1552), .B(n1626), .ZN(n891) );
  AOI221_X1 U1240 ( .B1(B[13]), .B2(n1582), .C1(B[12]), .C2(n1581), .A(n1627), 
        .ZN(n1626) );
  OAI22_X1 U1241 ( .A1(n1576), .A2(n1628), .B1(n1586), .B2(n1629), .ZN(n1627)
         );
  XNOR2_X1 U1242 ( .A(n1552), .B(n1630), .ZN(n890) );
  AOI221_X1 U1243 ( .B1(B[14]), .B2(n1582), .C1(B[13]), .C2(n1581), .A(n1631), 
        .ZN(n1630) );
  OAI22_X1 U1244 ( .A1(n1576), .A2(n1632), .B1(n1586), .B2(n1633), .ZN(n1631)
         );
  XNOR2_X1 U1245 ( .A(n1552), .B(n1634), .ZN(n889) );
  AOI221_X1 U1246 ( .B1(B[15]), .B2(n1582), .C1(B[14]), .C2(n1581), .A(n1635), 
        .ZN(n1634) );
  OAI22_X1 U1247 ( .A1(n1576), .A2(n1636), .B1(n1586), .B2(n1637), .ZN(n1635)
         );
  XNOR2_X1 U1248 ( .A(n1552), .B(n1638), .ZN(n888) );
  AOI221_X1 U1249 ( .B1(B[16]), .B2(n1582), .C1(B[15]), .C2(n1581), .A(n1639), 
        .ZN(n1638) );
  OAI22_X1 U1250 ( .A1(n1576), .A2(n1640), .B1(n1586), .B2(n1641), .ZN(n1639)
         );
  XNOR2_X1 U1251 ( .A(n1552), .B(n1642), .ZN(n887) );
  AOI221_X1 U1252 ( .B1(B[17]), .B2(n1582), .C1(B[16]), .C2(n1581), .A(n1643), 
        .ZN(n1642) );
  OAI22_X1 U1253 ( .A1(n1576), .A2(n1644), .B1(n1586), .B2(n1645), .ZN(n1643)
         );
  XNOR2_X1 U1254 ( .A(n1552), .B(n1646), .ZN(n886) );
  AOI221_X1 U1255 ( .B1(B[18]), .B2(n1582), .C1(B[17]), .C2(n1581), .A(n1647), 
        .ZN(n1646) );
  OAI22_X1 U1256 ( .A1(n1576), .A2(n1648), .B1(n1586), .B2(n1649), .ZN(n1647)
         );
  XNOR2_X1 U1257 ( .A(n1552), .B(n1650), .ZN(n885) );
  AOI221_X1 U1258 ( .B1(B[19]), .B2(n1582), .C1(B[18]), .C2(n1581), .A(n1651), 
        .ZN(n1650) );
  OAI22_X1 U1259 ( .A1(n1576), .A2(n1652), .B1(n1586), .B2(n1653), .ZN(n1651)
         );
  XNOR2_X1 U1260 ( .A(A[5]), .B(n1654), .ZN(n884) );
  AOI221_X1 U1261 ( .B1(n1582), .B2(B[20]), .C1(B[19]), .C2(n1581), .A(n1655), 
        .ZN(n1654) );
  OAI22_X1 U1262 ( .A1(n1576), .A2(n1656), .B1(n1586), .B2(n1657), .ZN(n1655)
         );
  XNOR2_X1 U1263 ( .A(A[5]), .B(n1658), .ZN(n883) );
  AOI221_X1 U1264 ( .B1(n1582), .B2(B[21]), .C1(n1581), .C2(B[20]), .A(n1659), 
        .ZN(n1658) );
  OAI22_X1 U1265 ( .A1(n1576), .A2(n1660), .B1(n1586), .B2(n1661), .ZN(n1659)
         );
  XNOR2_X1 U1266 ( .A(A[5]), .B(n1662), .ZN(n882) );
  AOI221_X1 U1267 ( .B1(n1582), .B2(B[22]), .C1(n1581), .C2(B[21]), .A(n1663), 
        .ZN(n1662) );
  OAI22_X1 U1268 ( .A1(n1562), .A2(n1576), .B1(n1564), .B2(n1586), .ZN(n1663)
         );
  XNOR2_X1 U1269 ( .A(A[5]), .B(n1664), .ZN(n881) );
  AOI221_X1 U1270 ( .B1(n1582), .B2(B[23]), .C1(n1581), .C2(B[22]), .A(n1665), 
        .ZN(n1664) );
  OAI22_X1 U1271 ( .A1(n1567), .A2(n1576), .B1(n1568), .B2(n1586), .ZN(n1665)
         );
  XNOR2_X1 U1272 ( .A(A[5]), .B(n1666), .ZN(n880) );
  AOI221_X1 U1273 ( .B1(n1582), .B2(B[23]), .C1(n1581), .C2(n1554), .A(n1667), 
        .ZN(n1666) );
  OAI22_X1 U1274 ( .A1(n1571), .A2(n1576), .B1(n1572), .B2(n1586), .ZN(n1667)
         );
  XNOR2_X1 U1275 ( .A(n1552), .B(n1668), .ZN(n879) );
  OAI221_X1 U1276 ( .B1(n1556), .B2(n1586), .C1(n1556), .C2(n1576), .A(n1669), 
        .ZN(n1668) );
  OAI21_X1 U1277 ( .B1(n1582), .B2(n1581), .A(n1554), .ZN(n1669) );
  INV_X1 U1278 ( .A(n1673), .ZN(n1670) );
  XNOR2_X1 U1279 ( .A(A[3]), .B(A[4]), .ZN(n1671) );
  XNOR2_X1 U1280 ( .A(A[4]), .B(n1553), .ZN(n1672) );
  XOR2_X1 U1281 ( .A(A[3]), .B(n1674), .Z(n1673) );
  XNOR2_X1 U1282 ( .A(n1675), .B(n1551), .ZN(n878) );
  OAI22_X1 U1283 ( .A1(n1574), .A2(n1676), .B1(n1574), .B2(n1677), .ZN(n1675)
         );
  XNOR2_X1 U1284 ( .A(n1678), .B(n1551), .ZN(n877) );
  OAI222_X1 U1285 ( .A1(n1578), .A2(n1676), .B1(n1574), .B2(n1679), .C1(n1580), 
        .C2(n1677), .ZN(n1678) );
  INV_X1 U1286 ( .A(n1680), .ZN(n1679) );
  INV_X1 U1287 ( .A(n1681), .ZN(n1676) );
  XNOR2_X1 U1288 ( .A(n1550), .B(n1682), .ZN(n876) );
  AOI221_X1 U1289 ( .B1(n1681), .B2(B[2]), .C1(n1680), .C2(B[1]), .A(n1683), 
        .ZN(n1682) );
  OAI22_X1 U1290 ( .A1(n1585), .A2(n1677), .B1(n1574), .B2(n1684), .ZN(n1683)
         );
  XNOR2_X1 U1291 ( .A(n1550), .B(n1685), .ZN(n875) );
  AOI221_X1 U1292 ( .B1(n1681), .B2(B[3]), .C1(n1680), .C2(B[2]), .A(n1686), 
        .ZN(n1685) );
  OAI22_X1 U1293 ( .A1(n1589), .A2(n1677), .B1(n1578), .B2(n1684), .ZN(n1686)
         );
  XNOR2_X1 U1294 ( .A(n1550), .B(n1687), .ZN(n874) );
  AOI221_X1 U1295 ( .B1(n1681), .B2(B[4]), .C1(n1680), .C2(B[3]), .A(n1688), 
        .ZN(n1687) );
  OAI22_X1 U1296 ( .A1(n1592), .A2(n1677), .B1(n1593), .B2(n1684), .ZN(n1688)
         );
  XNOR2_X1 U1297 ( .A(n1550), .B(n1689), .ZN(n873) );
  AOI221_X1 U1298 ( .B1(n1681), .B2(B[5]), .C1(n1680), .C2(B[4]), .A(n1690), 
        .ZN(n1689) );
  OAI22_X1 U1299 ( .A1(n1596), .A2(n1677), .B1(n1597), .B2(n1684), .ZN(n1690)
         );
  XNOR2_X1 U1300 ( .A(n1550), .B(n1691), .ZN(n872) );
  AOI221_X1 U1301 ( .B1(n1681), .B2(B[6]), .C1(n1680), .C2(B[5]), .A(n1692), 
        .ZN(n1691) );
  OAI22_X1 U1302 ( .A1(n1600), .A2(n1677), .B1(n1601), .B2(n1684), .ZN(n1692)
         );
  XNOR2_X1 U1303 ( .A(n1550), .B(n1693), .ZN(n871) );
  AOI221_X1 U1304 ( .B1(n1681), .B2(B[7]), .C1(n1680), .C2(B[6]), .A(n1694), 
        .ZN(n1693) );
  OAI22_X1 U1305 ( .A1(n1604), .A2(n1677), .B1(n1605), .B2(n1684), .ZN(n1694)
         );
  XNOR2_X1 U1306 ( .A(n1550), .B(n1695), .ZN(n870) );
  AOI221_X1 U1307 ( .B1(n1681), .B2(B[8]), .C1(n1680), .C2(B[7]), .A(n1696), 
        .ZN(n1695) );
  OAI22_X1 U1308 ( .A1(n1608), .A2(n1677), .B1(n1609), .B2(n1684), .ZN(n1696)
         );
  XNOR2_X1 U1309 ( .A(n1550), .B(n1697), .ZN(n869) );
  AOI221_X1 U1310 ( .B1(n1681), .B2(B[9]), .C1(n1680), .C2(B[8]), .A(n1698), 
        .ZN(n1697) );
  OAI22_X1 U1311 ( .A1(n1612), .A2(n1677), .B1(n1613), .B2(n1684), .ZN(n1698)
         );
  XNOR2_X1 U1312 ( .A(n1550), .B(n1699), .ZN(n868) );
  AOI221_X1 U1313 ( .B1(n1681), .B2(B[10]), .C1(n1680), .C2(B[9]), .A(n1700), 
        .ZN(n1699) );
  OAI22_X1 U1314 ( .A1(n1616), .A2(n1677), .B1(n1617), .B2(n1684), .ZN(n1700)
         );
  XNOR2_X1 U1315 ( .A(n1550), .B(n1701), .ZN(n867) );
  AOI221_X1 U1316 ( .B1(n1681), .B2(B[11]), .C1(n1680), .C2(B[10]), .A(n1702), 
        .ZN(n1701) );
  OAI22_X1 U1317 ( .A1(n1620), .A2(n1677), .B1(n1621), .B2(n1684), .ZN(n1702)
         );
  XNOR2_X1 U1318 ( .A(n1550), .B(n1703), .ZN(n866) );
  AOI221_X1 U1319 ( .B1(n1681), .B2(B[12]), .C1(n1680), .C2(B[11]), .A(n1704), 
        .ZN(n1703) );
  OAI22_X1 U1320 ( .A1(n1624), .A2(n1677), .B1(n1625), .B2(n1684), .ZN(n1704)
         );
  XNOR2_X1 U1321 ( .A(n1550), .B(n1705), .ZN(n865) );
  AOI221_X1 U1322 ( .B1(n1681), .B2(B[13]), .C1(n1680), .C2(B[12]), .A(n1706), 
        .ZN(n1705) );
  OAI22_X1 U1323 ( .A1(n1628), .A2(n1677), .B1(n1629), .B2(n1684), .ZN(n1706)
         );
  XNOR2_X1 U1324 ( .A(n1550), .B(n1707), .ZN(n864) );
  AOI221_X1 U1325 ( .B1(n1681), .B2(B[14]), .C1(n1680), .C2(B[13]), .A(n1708), 
        .ZN(n1707) );
  OAI22_X1 U1326 ( .A1(n1632), .A2(n1677), .B1(n1633), .B2(n1684), .ZN(n1708)
         );
  XNOR2_X1 U1327 ( .A(n1550), .B(n1709), .ZN(n863) );
  AOI221_X1 U1328 ( .B1(n1681), .B2(B[15]), .C1(n1680), .C2(B[14]), .A(n1710), 
        .ZN(n1709) );
  OAI22_X1 U1329 ( .A1(n1636), .A2(n1677), .B1(n1637), .B2(n1684), .ZN(n1710)
         );
  XNOR2_X1 U1330 ( .A(n1550), .B(n1711), .ZN(n862) );
  AOI221_X1 U1331 ( .B1(n1681), .B2(B[16]), .C1(n1680), .C2(B[15]), .A(n1712), 
        .ZN(n1711) );
  OAI22_X1 U1332 ( .A1(n1640), .A2(n1677), .B1(n1641), .B2(n1684), .ZN(n1712)
         );
  XNOR2_X1 U1333 ( .A(n1550), .B(n1713), .ZN(n861) );
  AOI221_X1 U1334 ( .B1(n1681), .B2(B[17]), .C1(n1680), .C2(B[16]), .A(n1714), 
        .ZN(n1713) );
  OAI22_X1 U1335 ( .A1(n1644), .A2(n1677), .B1(n1645), .B2(n1684), .ZN(n1714)
         );
  XNOR2_X1 U1336 ( .A(n1550), .B(n1715), .ZN(n860) );
  AOI221_X1 U1337 ( .B1(n1681), .B2(B[18]), .C1(n1680), .C2(B[17]), .A(n1716), 
        .ZN(n1715) );
  OAI22_X1 U1338 ( .A1(n1648), .A2(n1677), .B1(n1649), .B2(n1684), .ZN(n1716)
         );
  XNOR2_X1 U1339 ( .A(n1550), .B(n1717), .ZN(n859) );
  AOI221_X1 U1340 ( .B1(n1681), .B2(B[19]), .C1(n1680), .C2(B[18]), .A(n1718), 
        .ZN(n1717) );
  OAI22_X1 U1341 ( .A1(n1652), .A2(n1677), .B1(n1653), .B2(n1684), .ZN(n1718)
         );
  XNOR2_X1 U1342 ( .A(A[8]), .B(n1719), .ZN(n858) );
  AOI221_X1 U1343 ( .B1(n1681), .B2(B[20]), .C1(n1680), .C2(B[19]), .A(n1720), 
        .ZN(n1719) );
  OAI22_X1 U1344 ( .A1(n1656), .A2(n1677), .B1(n1657), .B2(n1684), .ZN(n1720)
         );
  XNOR2_X1 U1345 ( .A(A[8]), .B(n1721), .ZN(n857) );
  AOI221_X1 U1346 ( .B1(n1681), .B2(B[21]), .C1(n1680), .C2(B[20]), .A(n1722), 
        .ZN(n1721) );
  OAI22_X1 U1347 ( .A1(n1660), .A2(n1677), .B1(n1661), .B2(n1684), .ZN(n1722)
         );
  XNOR2_X1 U1348 ( .A(A[8]), .B(n1723), .ZN(n856) );
  AOI221_X1 U1349 ( .B1(n1681), .B2(B[22]), .C1(n1680), .C2(B[21]), .A(n1724), 
        .ZN(n1723) );
  OAI22_X1 U1350 ( .A1(n1562), .A2(n1677), .B1(n1564), .B2(n1684), .ZN(n1724)
         );
  XNOR2_X1 U1351 ( .A(A[8]), .B(n1725), .ZN(n855) );
  AOI221_X1 U1352 ( .B1(n1681), .B2(B[23]), .C1(n1680), .C2(B[22]), .A(n1726), 
        .ZN(n1725) );
  OAI22_X1 U1353 ( .A1(n1567), .A2(n1677), .B1(n1568), .B2(n1684), .ZN(n1726)
         );
  XNOR2_X1 U1354 ( .A(A[8]), .B(n1727), .ZN(n854) );
  AOI221_X1 U1355 ( .B1(n1681), .B2(B[23]), .C1(n1680), .C2(n1554), .A(n1728), 
        .ZN(n1727) );
  OAI22_X1 U1356 ( .A1(n1571), .A2(n1677), .B1(n1572), .B2(n1684), .ZN(n1728)
         );
  XNOR2_X1 U1357 ( .A(n1550), .B(n1729), .ZN(n853) );
  OAI221_X1 U1358 ( .B1(n1555), .B2(n1684), .C1(n1556), .C2(n1677), .A(n1730), 
        .ZN(n1729) );
  OAI21_X1 U1359 ( .B1(n1681), .B2(n1680), .A(n1554), .ZN(n1730) );
  INV_X1 U1360 ( .A(n1734), .ZN(n1731) );
  XNOR2_X1 U1361 ( .A(A[6]), .B(A[7]), .ZN(n1732) );
  XNOR2_X1 U1362 ( .A(A[7]), .B(n1551), .ZN(n1733) );
  XOR2_X1 U1363 ( .A(A[6]), .B(n1553), .Z(n1734) );
  XNOR2_X1 U1364 ( .A(n1735), .B(n1549), .ZN(n852) );
  OAI22_X1 U1365 ( .A1(n1574), .A2(n1736), .B1(n1574), .B2(n1737), .ZN(n1735)
         );
  XNOR2_X1 U1366 ( .A(n1738), .B(n1549), .ZN(n851) );
  OAI222_X1 U1367 ( .A1(n1578), .A2(n1736), .B1(n1574), .B2(n1739), .C1(n1580), 
        .C2(n1737), .ZN(n1738) );
  INV_X1 U1368 ( .A(n1740), .ZN(n1739) );
  INV_X1 U1369 ( .A(n1741), .ZN(n1736) );
  XNOR2_X1 U1370 ( .A(n1548), .B(n1742), .ZN(n850) );
  AOI221_X1 U1371 ( .B1(n1741), .B2(B[2]), .C1(n1740), .C2(B[1]), .A(n1743), 
        .ZN(n1742) );
  OAI22_X1 U1372 ( .A1(n1585), .A2(n1737), .B1(n1574), .B2(n1744), .ZN(n1743)
         );
  XNOR2_X1 U1373 ( .A(n1548), .B(n1745), .ZN(n849) );
  AOI221_X1 U1374 ( .B1(n1741), .B2(B[3]), .C1(n1740), .C2(B[2]), .A(n1746), 
        .ZN(n1745) );
  OAI22_X1 U1375 ( .A1(n1589), .A2(n1737), .B1(n1578), .B2(n1744), .ZN(n1746)
         );
  XNOR2_X1 U1376 ( .A(n1548), .B(n1747), .ZN(n848) );
  AOI221_X1 U1377 ( .B1(n1741), .B2(B[4]), .C1(n1740), .C2(B[3]), .A(n1748), 
        .ZN(n1747) );
  OAI22_X1 U1378 ( .A1(n1592), .A2(n1737), .B1(n1593), .B2(n1744), .ZN(n1748)
         );
  XNOR2_X1 U1379 ( .A(n1548), .B(n1749), .ZN(n847) );
  AOI221_X1 U1380 ( .B1(n1741), .B2(B[5]), .C1(n1740), .C2(B[4]), .A(n1750), 
        .ZN(n1749) );
  OAI22_X1 U1381 ( .A1(n1596), .A2(n1737), .B1(n1597), .B2(n1744), .ZN(n1750)
         );
  XNOR2_X1 U1382 ( .A(n1548), .B(n1751), .ZN(n846) );
  AOI221_X1 U1383 ( .B1(n1741), .B2(B[6]), .C1(n1740), .C2(B[5]), .A(n1752), 
        .ZN(n1751) );
  OAI22_X1 U1384 ( .A1(n1600), .A2(n1737), .B1(n1601), .B2(n1744), .ZN(n1752)
         );
  XNOR2_X1 U1385 ( .A(n1548), .B(n1753), .ZN(n845) );
  AOI221_X1 U1386 ( .B1(n1741), .B2(B[7]), .C1(n1740), .C2(B[6]), .A(n1754), 
        .ZN(n1753) );
  OAI22_X1 U1387 ( .A1(n1604), .A2(n1737), .B1(n1605), .B2(n1744), .ZN(n1754)
         );
  XNOR2_X1 U1388 ( .A(n1548), .B(n1755), .ZN(n844) );
  AOI221_X1 U1389 ( .B1(n1741), .B2(B[8]), .C1(n1740), .C2(B[7]), .A(n1756), 
        .ZN(n1755) );
  OAI22_X1 U1390 ( .A1(n1608), .A2(n1737), .B1(n1609), .B2(n1744), .ZN(n1756)
         );
  XNOR2_X1 U1391 ( .A(n1548), .B(n1757), .ZN(n843) );
  AOI221_X1 U1392 ( .B1(n1741), .B2(B[9]), .C1(n1740), .C2(B[8]), .A(n1758), 
        .ZN(n1757) );
  OAI22_X1 U1393 ( .A1(n1612), .A2(n1737), .B1(n1613), .B2(n1744), .ZN(n1758)
         );
  XNOR2_X1 U1394 ( .A(n1548), .B(n1759), .ZN(n842) );
  AOI221_X1 U1395 ( .B1(n1741), .B2(B[10]), .C1(n1740), .C2(B[9]), .A(n1760), 
        .ZN(n1759) );
  OAI22_X1 U1396 ( .A1(n1616), .A2(n1737), .B1(n1617), .B2(n1744), .ZN(n1760)
         );
  XNOR2_X1 U1397 ( .A(n1548), .B(n1761), .ZN(n841) );
  AOI221_X1 U1398 ( .B1(n1741), .B2(B[11]), .C1(n1740), .C2(B[10]), .A(n1762), 
        .ZN(n1761) );
  OAI22_X1 U1399 ( .A1(n1620), .A2(n1737), .B1(n1621), .B2(n1744), .ZN(n1762)
         );
  XNOR2_X1 U1400 ( .A(n1548), .B(n1763), .ZN(n840) );
  AOI221_X1 U1401 ( .B1(n1741), .B2(B[12]), .C1(n1740), .C2(B[11]), .A(n1764), 
        .ZN(n1763) );
  OAI22_X1 U1402 ( .A1(n1624), .A2(n1737), .B1(n1625), .B2(n1744), .ZN(n1764)
         );
  XNOR2_X1 U1403 ( .A(n1548), .B(n1765), .ZN(n839) );
  AOI221_X1 U1404 ( .B1(n1741), .B2(B[13]), .C1(n1740), .C2(B[12]), .A(n1766), 
        .ZN(n1765) );
  OAI22_X1 U1405 ( .A1(n1628), .A2(n1737), .B1(n1629), .B2(n1744), .ZN(n1766)
         );
  XNOR2_X1 U1406 ( .A(n1548), .B(n1767), .ZN(n838) );
  AOI221_X1 U1407 ( .B1(n1741), .B2(B[14]), .C1(n1740), .C2(B[13]), .A(n1768), 
        .ZN(n1767) );
  OAI22_X1 U1408 ( .A1(n1632), .A2(n1737), .B1(n1633), .B2(n1744), .ZN(n1768)
         );
  XNOR2_X1 U1409 ( .A(n1548), .B(n1769), .ZN(n837) );
  AOI221_X1 U1410 ( .B1(n1741), .B2(B[15]), .C1(n1740), .C2(B[14]), .A(n1770), 
        .ZN(n1769) );
  OAI22_X1 U1411 ( .A1(n1636), .A2(n1737), .B1(n1637), .B2(n1744), .ZN(n1770)
         );
  XNOR2_X1 U1412 ( .A(n1548), .B(n1771), .ZN(n836) );
  AOI221_X1 U1413 ( .B1(n1741), .B2(B[16]), .C1(n1740), .C2(B[15]), .A(n1772), 
        .ZN(n1771) );
  OAI22_X1 U1414 ( .A1(n1640), .A2(n1737), .B1(n1641), .B2(n1744), .ZN(n1772)
         );
  XNOR2_X1 U1415 ( .A(n1548), .B(n1773), .ZN(n835) );
  AOI221_X1 U1416 ( .B1(n1741), .B2(B[17]), .C1(n1740), .C2(B[16]), .A(n1774), 
        .ZN(n1773) );
  OAI22_X1 U1417 ( .A1(n1644), .A2(n1737), .B1(n1645), .B2(n1744), .ZN(n1774)
         );
  XNOR2_X1 U1418 ( .A(n1548), .B(n1775), .ZN(n834) );
  AOI221_X1 U1419 ( .B1(n1741), .B2(B[18]), .C1(n1740), .C2(B[17]), .A(n1776), 
        .ZN(n1775) );
  OAI22_X1 U1420 ( .A1(n1648), .A2(n1737), .B1(n1649), .B2(n1744), .ZN(n1776)
         );
  XNOR2_X1 U1421 ( .A(n1548), .B(n1777), .ZN(n833) );
  AOI221_X1 U1422 ( .B1(n1741), .B2(B[19]), .C1(n1740), .C2(B[18]), .A(n1778), 
        .ZN(n1777) );
  OAI22_X1 U1423 ( .A1(n1652), .A2(n1737), .B1(n1653), .B2(n1744), .ZN(n1778)
         );
  XNOR2_X1 U1424 ( .A(n1548), .B(n1779), .ZN(n832) );
  AOI221_X1 U1425 ( .B1(n1741), .B2(B[20]), .C1(n1740), .C2(B[19]), .A(n1780), 
        .ZN(n1779) );
  OAI22_X1 U1426 ( .A1(n1656), .A2(n1737), .B1(n1657), .B2(n1744), .ZN(n1780)
         );
  XNOR2_X1 U1427 ( .A(A[11]), .B(n1781), .ZN(n831) );
  AOI221_X1 U1428 ( .B1(n1741), .B2(B[21]), .C1(n1740), .C2(B[20]), .A(n1782), 
        .ZN(n1781) );
  OAI22_X1 U1429 ( .A1(n1660), .A2(n1737), .B1(n1661), .B2(n1744), .ZN(n1782)
         );
  XNOR2_X1 U1430 ( .A(A[11]), .B(n1783), .ZN(n830) );
  AOI221_X1 U1431 ( .B1(n1741), .B2(B[22]), .C1(n1740), .C2(B[21]), .A(n1784), 
        .ZN(n1783) );
  OAI22_X1 U1432 ( .A1(n1562), .A2(n1737), .B1(n1564), .B2(n1744), .ZN(n1784)
         );
  XNOR2_X1 U1433 ( .A(A[11]), .B(n1785), .ZN(n829) );
  AOI221_X1 U1434 ( .B1(n1741), .B2(B[23]), .C1(n1740), .C2(B[22]), .A(n1786), 
        .ZN(n1785) );
  OAI22_X1 U1435 ( .A1(n1567), .A2(n1737), .B1(n1568), .B2(n1744), .ZN(n1786)
         );
  XNOR2_X1 U1436 ( .A(A[11]), .B(n1787), .ZN(n828) );
  AOI221_X1 U1437 ( .B1(n1741), .B2(B[23]), .C1(n1740), .C2(n1554), .A(n1788), 
        .ZN(n1787) );
  OAI22_X1 U1438 ( .A1(n1571), .A2(n1737), .B1(n1572), .B2(n1744), .ZN(n1788)
         );
  XNOR2_X1 U1439 ( .A(A[11]), .B(n1789), .ZN(n827) );
  OAI221_X1 U1440 ( .B1(n1556), .B2(n1744), .C1(n1556), .C2(n1737), .A(n1790), 
        .ZN(n1789) );
  OAI21_X1 U1441 ( .B1(n1741), .B2(n1740), .A(n1554), .ZN(n1790) );
  INV_X1 U1442 ( .A(n1794), .ZN(n1791) );
  XNOR2_X1 U1443 ( .A(A[10]), .B(A[9]), .ZN(n1792) );
  XNOR2_X1 U1444 ( .A(A[10]), .B(n1549), .ZN(n1793) );
  XOR2_X1 U1445 ( .A(A[9]), .B(n1551), .Z(n1794) );
  XNOR2_X1 U1446 ( .A(n1795), .B(n1547), .ZN(n826) );
  OAI22_X1 U1447 ( .A1(n1574), .A2(n1796), .B1(n1574), .B2(n1797), .ZN(n1795)
         );
  XNOR2_X1 U1448 ( .A(n1798), .B(n1547), .ZN(n825) );
  OAI222_X1 U1449 ( .A1(n1578), .A2(n1796), .B1(n1574), .B2(n1799), .C1(n1580), 
        .C2(n1797), .ZN(n1798) );
  INV_X1 U1450 ( .A(n1800), .ZN(n1799) );
  INV_X1 U1451 ( .A(n1801), .ZN(n1796) );
  XNOR2_X1 U1452 ( .A(n1546), .B(n1802), .ZN(n824) );
  AOI221_X1 U1453 ( .B1(n1801), .B2(B[2]), .C1(n1800), .C2(B[1]), .A(n1803), 
        .ZN(n1802) );
  OAI22_X1 U1454 ( .A1(n1585), .A2(n1797), .B1(n1574), .B2(n1804), .ZN(n1803)
         );
  XNOR2_X1 U1455 ( .A(n1546), .B(n1805), .ZN(n823) );
  AOI221_X1 U1456 ( .B1(n1801), .B2(B[3]), .C1(n1800), .C2(B[2]), .A(n1806), 
        .ZN(n1805) );
  OAI22_X1 U1457 ( .A1(n1589), .A2(n1797), .B1(n1578), .B2(n1804), .ZN(n1806)
         );
  XNOR2_X1 U1458 ( .A(n1546), .B(n1807), .ZN(n822) );
  AOI221_X1 U1459 ( .B1(n1801), .B2(B[4]), .C1(n1800), .C2(B[3]), .A(n1808), 
        .ZN(n1807) );
  OAI22_X1 U1460 ( .A1(n1592), .A2(n1797), .B1(n1593), .B2(n1804), .ZN(n1808)
         );
  XNOR2_X1 U1461 ( .A(n1546), .B(n1809), .ZN(n821) );
  AOI221_X1 U1462 ( .B1(n1801), .B2(B[5]), .C1(n1800), .C2(B[4]), .A(n1810), 
        .ZN(n1809) );
  OAI22_X1 U1463 ( .A1(n1596), .A2(n1797), .B1(n1597), .B2(n1804), .ZN(n1810)
         );
  XNOR2_X1 U1464 ( .A(n1546), .B(n1811), .ZN(n820) );
  AOI221_X1 U1465 ( .B1(n1801), .B2(B[6]), .C1(n1800), .C2(B[5]), .A(n1812), 
        .ZN(n1811) );
  OAI22_X1 U1466 ( .A1(n1600), .A2(n1797), .B1(n1601), .B2(n1804), .ZN(n1812)
         );
  XNOR2_X1 U1467 ( .A(n1546), .B(n1813), .ZN(n819) );
  AOI221_X1 U1468 ( .B1(n1801), .B2(B[7]), .C1(n1800), .C2(B[6]), .A(n1814), 
        .ZN(n1813) );
  OAI22_X1 U1469 ( .A1(n1604), .A2(n1797), .B1(n1605), .B2(n1804), .ZN(n1814)
         );
  XNOR2_X1 U1470 ( .A(n1546), .B(n1815), .ZN(n818) );
  AOI221_X1 U1471 ( .B1(n1801), .B2(B[8]), .C1(n1800), .C2(B[7]), .A(n1816), 
        .ZN(n1815) );
  OAI22_X1 U1472 ( .A1(n1608), .A2(n1797), .B1(n1609), .B2(n1804), .ZN(n1816)
         );
  XNOR2_X1 U1473 ( .A(n1546), .B(n1817), .ZN(n817) );
  AOI221_X1 U1474 ( .B1(n1801), .B2(B[9]), .C1(n1800), .C2(B[8]), .A(n1818), 
        .ZN(n1817) );
  OAI22_X1 U1475 ( .A1(n1612), .A2(n1797), .B1(n1613), .B2(n1804), .ZN(n1818)
         );
  XNOR2_X1 U1476 ( .A(n1546), .B(n1819), .ZN(n816) );
  AOI221_X1 U1477 ( .B1(n1801), .B2(B[10]), .C1(n1800), .C2(B[9]), .A(n1820), 
        .ZN(n1819) );
  OAI22_X1 U1478 ( .A1(n1616), .A2(n1797), .B1(n1617), .B2(n1804), .ZN(n1820)
         );
  XNOR2_X1 U1479 ( .A(n1546), .B(n1821), .ZN(n815) );
  AOI221_X1 U1480 ( .B1(n1801), .B2(B[11]), .C1(n1800), .C2(B[10]), .A(n1822), 
        .ZN(n1821) );
  OAI22_X1 U1481 ( .A1(n1620), .A2(n1797), .B1(n1621), .B2(n1804), .ZN(n1822)
         );
  XNOR2_X1 U1482 ( .A(n1546), .B(n1823), .ZN(n814) );
  AOI221_X1 U1483 ( .B1(n1801), .B2(B[12]), .C1(n1800), .C2(B[11]), .A(n1824), 
        .ZN(n1823) );
  OAI22_X1 U1484 ( .A1(n1624), .A2(n1797), .B1(n1625), .B2(n1804), .ZN(n1824)
         );
  XNOR2_X1 U1485 ( .A(n1546), .B(n1825), .ZN(n813) );
  AOI221_X1 U1486 ( .B1(n1801), .B2(B[13]), .C1(n1800), .C2(B[12]), .A(n1826), 
        .ZN(n1825) );
  OAI22_X1 U1487 ( .A1(n1628), .A2(n1797), .B1(n1629), .B2(n1804), .ZN(n1826)
         );
  XNOR2_X1 U1488 ( .A(n1546), .B(n1827), .ZN(n812) );
  AOI221_X1 U1489 ( .B1(n1801), .B2(B[14]), .C1(n1800), .C2(B[13]), .A(n1828), 
        .ZN(n1827) );
  OAI22_X1 U1490 ( .A1(n1632), .A2(n1797), .B1(n1633), .B2(n1804), .ZN(n1828)
         );
  XNOR2_X1 U1491 ( .A(n1546), .B(n1829), .ZN(n811) );
  AOI221_X1 U1492 ( .B1(n1801), .B2(B[15]), .C1(n1800), .C2(B[14]), .A(n1830), 
        .ZN(n1829) );
  OAI22_X1 U1493 ( .A1(n1636), .A2(n1797), .B1(n1637), .B2(n1804), .ZN(n1830)
         );
  XNOR2_X1 U1494 ( .A(n1546), .B(n1831), .ZN(n810) );
  AOI221_X1 U1495 ( .B1(n1801), .B2(B[16]), .C1(n1800), .C2(B[15]), .A(n1832), 
        .ZN(n1831) );
  OAI22_X1 U1496 ( .A1(n1640), .A2(n1797), .B1(n1641), .B2(n1804), .ZN(n1832)
         );
  XNOR2_X1 U1497 ( .A(n1546), .B(n1833), .ZN(n809) );
  AOI221_X1 U1498 ( .B1(n1801), .B2(B[17]), .C1(n1800), .C2(B[16]), .A(n1834), 
        .ZN(n1833) );
  OAI22_X1 U1499 ( .A1(n1644), .A2(n1797), .B1(n1645), .B2(n1804), .ZN(n1834)
         );
  XNOR2_X1 U1500 ( .A(n1546), .B(n1835), .ZN(n808) );
  AOI221_X1 U1501 ( .B1(n1801), .B2(B[18]), .C1(n1800), .C2(B[17]), .A(n1836), 
        .ZN(n1835) );
  OAI22_X1 U1502 ( .A1(n1648), .A2(n1797), .B1(n1649), .B2(n1804), .ZN(n1836)
         );
  XNOR2_X1 U1503 ( .A(n1546), .B(n1837), .ZN(n807) );
  AOI221_X1 U1504 ( .B1(n1801), .B2(B[19]), .C1(n1800), .C2(B[18]), .A(n1838), 
        .ZN(n1837) );
  OAI22_X1 U1505 ( .A1(n1652), .A2(n1797), .B1(n1653), .B2(n1804), .ZN(n1838)
         );
  XNOR2_X1 U1506 ( .A(n1546), .B(n1839), .ZN(n806) );
  AOI221_X1 U1507 ( .B1(n1801), .B2(B[20]), .C1(n1800), .C2(B[19]), .A(n1840), 
        .ZN(n1839) );
  OAI22_X1 U1508 ( .A1(n1656), .A2(n1797), .B1(n1657), .B2(n1804), .ZN(n1840)
         );
  XNOR2_X1 U1509 ( .A(A[14]), .B(n1841), .ZN(n805) );
  AOI221_X1 U1510 ( .B1(n1801), .B2(B[21]), .C1(n1800), .C2(B[20]), .A(n1842), 
        .ZN(n1841) );
  OAI22_X1 U1511 ( .A1(n1660), .A2(n1797), .B1(n1661), .B2(n1804), .ZN(n1842)
         );
  XNOR2_X1 U1512 ( .A(A[14]), .B(n1843), .ZN(n804) );
  AOI221_X1 U1513 ( .B1(n1801), .B2(B[22]), .C1(n1800), .C2(B[21]), .A(n1844), 
        .ZN(n1843) );
  OAI22_X1 U1514 ( .A1(n1562), .A2(n1797), .B1(n1564), .B2(n1804), .ZN(n1844)
         );
  XNOR2_X1 U1515 ( .A(A[14]), .B(n1845), .ZN(n803) );
  AOI221_X1 U1516 ( .B1(n1801), .B2(B[23]), .C1(n1800), .C2(B[22]), .A(n1846), 
        .ZN(n1845) );
  OAI22_X1 U1517 ( .A1(n1567), .A2(n1797), .B1(n1568), .B2(n1804), .ZN(n1846)
         );
  XNOR2_X1 U1518 ( .A(A[14]), .B(n1847), .ZN(n802) );
  AOI221_X1 U1519 ( .B1(n1801), .B2(B[23]), .C1(n1800), .C2(n1554), .A(n1848), 
        .ZN(n1847) );
  OAI22_X1 U1520 ( .A1(n1571), .A2(n1797), .B1(n1572), .B2(n1804), .ZN(n1848)
         );
  XNOR2_X1 U1521 ( .A(A[14]), .B(n1849), .ZN(n801) );
  OAI221_X1 U1522 ( .B1(n1556), .B2(n1804), .C1(n1556), .C2(n1797), .A(n1850), 
        .ZN(n1849) );
  OAI21_X1 U1523 ( .B1(n1801), .B2(n1800), .A(n1554), .ZN(n1850) );
  INV_X1 U1524 ( .A(n1854), .ZN(n1851) );
  XNOR2_X1 U1525 ( .A(A[12]), .B(A[13]), .ZN(n1852) );
  XNOR2_X1 U1526 ( .A(A[13]), .B(n1547), .ZN(n1853) );
  XOR2_X1 U1527 ( .A(A[12]), .B(n1549), .Z(n1854) );
  XNOR2_X1 U1528 ( .A(n1855), .B(n1545), .ZN(n800) );
  OAI22_X1 U1529 ( .A1(n1574), .A2(n1856), .B1(n1574), .B2(n1857), .ZN(n1855)
         );
  XNOR2_X1 U1530 ( .A(n1858), .B(n1545), .ZN(n799) );
  OAI222_X1 U1531 ( .A1(n1578), .A2(n1856), .B1(n1574), .B2(n1859), .C1(n1580), 
        .C2(n1857), .ZN(n1858) );
  INV_X1 U1532 ( .A(n1860), .ZN(n1859) );
  INV_X1 U1533 ( .A(n1861), .ZN(n1856) );
  XNOR2_X1 U1534 ( .A(n1544), .B(n1862), .ZN(n798) );
  AOI221_X1 U1535 ( .B1(n1861), .B2(B[2]), .C1(n1860), .C2(B[1]), .A(n1863), 
        .ZN(n1862) );
  OAI22_X1 U1536 ( .A1(n1585), .A2(n1857), .B1(n1574), .B2(n1864), .ZN(n1863)
         );
  XNOR2_X1 U1537 ( .A(n1544), .B(n1865), .ZN(n797) );
  AOI221_X1 U1538 ( .B1(n1861), .B2(B[3]), .C1(n1860), .C2(B[2]), .A(n1866), 
        .ZN(n1865) );
  OAI22_X1 U1539 ( .A1(n1589), .A2(n1857), .B1(n1578), .B2(n1864), .ZN(n1866)
         );
  XNOR2_X1 U1540 ( .A(n1544), .B(n1867), .ZN(n796) );
  AOI221_X1 U1541 ( .B1(n1861), .B2(B[4]), .C1(n1860), .C2(B[3]), .A(n1868), 
        .ZN(n1867) );
  OAI22_X1 U1542 ( .A1(n1592), .A2(n1857), .B1(n1593), .B2(n1864), .ZN(n1868)
         );
  XNOR2_X1 U1543 ( .A(n1544), .B(n1869), .ZN(n795) );
  AOI221_X1 U1544 ( .B1(n1861), .B2(B[5]), .C1(n1860), .C2(B[4]), .A(n1870), 
        .ZN(n1869) );
  OAI22_X1 U1545 ( .A1(n1596), .A2(n1857), .B1(n1597), .B2(n1864), .ZN(n1870)
         );
  XNOR2_X1 U1546 ( .A(n1544), .B(n1871), .ZN(n794) );
  AOI221_X1 U1547 ( .B1(n1861), .B2(B[6]), .C1(n1860), .C2(B[5]), .A(n1872), 
        .ZN(n1871) );
  OAI22_X1 U1548 ( .A1(n1600), .A2(n1857), .B1(n1601), .B2(n1864), .ZN(n1872)
         );
  XNOR2_X1 U1549 ( .A(n1544), .B(n1873), .ZN(n793) );
  AOI221_X1 U1550 ( .B1(n1861), .B2(B[7]), .C1(n1860), .C2(B[6]), .A(n1874), 
        .ZN(n1873) );
  OAI22_X1 U1551 ( .A1(n1604), .A2(n1857), .B1(n1605), .B2(n1864), .ZN(n1874)
         );
  XNOR2_X1 U1552 ( .A(n1544), .B(n1875), .ZN(n792) );
  AOI221_X1 U1553 ( .B1(n1861), .B2(B[8]), .C1(n1860), .C2(B[7]), .A(n1876), 
        .ZN(n1875) );
  OAI22_X1 U1554 ( .A1(n1608), .A2(n1857), .B1(n1609), .B2(n1864), .ZN(n1876)
         );
  XNOR2_X1 U1555 ( .A(n1544), .B(n1877), .ZN(n791) );
  AOI221_X1 U1556 ( .B1(n1861), .B2(B[9]), .C1(n1860), .C2(B[8]), .A(n1878), 
        .ZN(n1877) );
  OAI22_X1 U1557 ( .A1(n1612), .A2(n1857), .B1(n1613), .B2(n1864), .ZN(n1878)
         );
  XNOR2_X1 U1558 ( .A(n1544), .B(n1879), .ZN(n790) );
  AOI221_X1 U1559 ( .B1(n1861), .B2(B[10]), .C1(n1860), .C2(B[9]), .A(n1880), 
        .ZN(n1879) );
  OAI22_X1 U1560 ( .A1(n1616), .A2(n1857), .B1(n1617), .B2(n1864), .ZN(n1880)
         );
  XNOR2_X1 U1561 ( .A(n1544), .B(n1881), .ZN(n789) );
  AOI221_X1 U1562 ( .B1(n1861), .B2(B[11]), .C1(n1860), .C2(B[10]), .A(n1882), 
        .ZN(n1881) );
  OAI22_X1 U1563 ( .A1(n1620), .A2(n1857), .B1(n1621), .B2(n1864), .ZN(n1882)
         );
  XNOR2_X1 U1564 ( .A(n1544), .B(n1883), .ZN(n788) );
  AOI221_X1 U1565 ( .B1(n1861), .B2(B[12]), .C1(n1860), .C2(B[11]), .A(n1884), 
        .ZN(n1883) );
  OAI22_X1 U1566 ( .A1(n1624), .A2(n1857), .B1(n1625), .B2(n1864), .ZN(n1884)
         );
  XNOR2_X1 U1567 ( .A(n1544), .B(n1885), .ZN(n787) );
  AOI221_X1 U1568 ( .B1(n1861), .B2(B[13]), .C1(n1860), .C2(B[12]), .A(n1886), 
        .ZN(n1885) );
  OAI22_X1 U1569 ( .A1(n1628), .A2(n1857), .B1(n1629), .B2(n1864), .ZN(n1886)
         );
  XNOR2_X1 U1570 ( .A(n1544), .B(n1887), .ZN(n786) );
  AOI221_X1 U1571 ( .B1(n1861), .B2(B[14]), .C1(n1860), .C2(B[13]), .A(n1888), 
        .ZN(n1887) );
  OAI22_X1 U1572 ( .A1(n1632), .A2(n1857), .B1(n1633), .B2(n1864), .ZN(n1888)
         );
  XNOR2_X1 U1573 ( .A(n1544), .B(n1889), .ZN(n785) );
  AOI221_X1 U1574 ( .B1(n1861), .B2(B[15]), .C1(n1860), .C2(B[14]), .A(n1890), 
        .ZN(n1889) );
  OAI22_X1 U1575 ( .A1(n1636), .A2(n1857), .B1(n1637), .B2(n1864), .ZN(n1890)
         );
  XNOR2_X1 U1576 ( .A(n1544), .B(n1891), .ZN(n784) );
  AOI221_X1 U1577 ( .B1(n1861), .B2(B[16]), .C1(n1860), .C2(B[15]), .A(n1892), 
        .ZN(n1891) );
  OAI22_X1 U1578 ( .A1(n1640), .A2(n1857), .B1(n1641), .B2(n1864), .ZN(n1892)
         );
  XNOR2_X1 U1579 ( .A(n1544), .B(n1893), .ZN(n783) );
  AOI221_X1 U1580 ( .B1(n1861), .B2(B[17]), .C1(n1860), .C2(B[16]), .A(n1894), 
        .ZN(n1893) );
  OAI22_X1 U1581 ( .A1(n1644), .A2(n1857), .B1(n1645), .B2(n1864), .ZN(n1894)
         );
  XNOR2_X1 U1582 ( .A(n1544), .B(n1895), .ZN(n782) );
  AOI221_X1 U1583 ( .B1(n1861), .B2(B[18]), .C1(n1860), .C2(B[17]), .A(n1896), 
        .ZN(n1895) );
  OAI22_X1 U1584 ( .A1(n1648), .A2(n1857), .B1(n1649), .B2(n1864), .ZN(n1896)
         );
  XNOR2_X1 U1585 ( .A(n1544), .B(n1897), .ZN(n781) );
  AOI221_X1 U1586 ( .B1(n1861), .B2(B[19]), .C1(n1860), .C2(B[18]), .A(n1898), 
        .ZN(n1897) );
  OAI22_X1 U1587 ( .A1(n1652), .A2(n1857), .B1(n1653), .B2(n1864), .ZN(n1898)
         );
  XNOR2_X1 U1588 ( .A(n1544), .B(n1899), .ZN(n780) );
  AOI221_X1 U1589 ( .B1(n1861), .B2(B[20]), .C1(n1860), .C2(B[19]), .A(n1900), 
        .ZN(n1899) );
  OAI22_X1 U1590 ( .A1(n1656), .A2(n1857), .B1(n1657), .B2(n1864), .ZN(n1900)
         );
  XNOR2_X1 U1591 ( .A(A[17]), .B(n1901), .ZN(n779) );
  AOI221_X1 U1592 ( .B1(n1861), .B2(B[21]), .C1(n1860), .C2(B[20]), .A(n1902), 
        .ZN(n1901) );
  OAI22_X1 U1593 ( .A1(n1660), .A2(n1857), .B1(n1661), .B2(n1864), .ZN(n1902)
         );
  XNOR2_X1 U1594 ( .A(A[17]), .B(n1903), .ZN(n778) );
  AOI221_X1 U1595 ( .B1(n1861), .B2(B[22]), .C1(n1860), .C2(B[21]), .A(n1904), 
        .ZN(n1903) );
  OAI22_X1 U1596 ( .A1(n1562), .A2(n1857), .B1(n1564), .B2(n1864), .ZN(n1904)
         );
  XNOR2_X1 U1597 ( .A(A[17]), .B(n1905), .ZN(n777) );
  AOI221_X1 U1598 ( .B1(n1861), .B2(B[23]), .C1(n1860), .C2(B[22]), .A(n1906), 
        .ZN(n1905) );
  OAI22_X1 U1599 ( .A1(n1567), .A2(n1857), .B1(n1568), .B2(n1864), .ZN(n1906)
         );
  XNOR2_X1 U1600 ( .A(A[17]), .B(n1907), .ZN(n776) );
  AOI221_X1 U1601 ( .B1(n1861), .B2(B[23]), .C1(n1860), .C2(n1554), .A(n1908), 
        .ZN(n1907) );
  OAI22_X1 U1602 ( .A1(n1571), .A2(n1857), .B1(n1572), .B2(n1864), .ZN(n1908)
         );
  XNOR2_X1 U1603 ( .A(A[17]), .B(n1909), .ZN(n775) );
  OAI221_X1 U1604 ( .B1(n1556), .B2(n1864), .C1(n1556), .C2(n1857), .A(n1910), 
        .ZN(n1909) );
  OAI21_X1 U1605 ( .B1(n1861), .B2(n1860), .A(n1554), .ZN(n1910) );
  INV_X1 U1606 ( .A(n1914), .ZN(n1911) );
  XNOR2_X1 U1607 ( .A(A[15]), .B(A[16]), .ZN(n1912) );
  XNOR2_X1 U1608 ( .A(A[16]), .B(n1545), .ZN(n1913) );
  XOR2_X1 U1609 ( .A(A[15]), .B(n1547), .Z(n1914) );
  XNOR2_X1 U1610 ( .A(n1915), .B(n1543), .ZN(n774) );
  OAI22_X1 U1611 ( .A1(n1574), .A2(n1916), .B1(n1574), .B2(n1917), .ZN(n1915)
         );
  XNOR2_X1 U1612 ( .A(n1918), .B(n1543), .ZN(n773) );
  OAI222_X1 U1613 ( .A1(n1578), .A2(n1916), .B1(n1574), .B2(n1919), .C1(n1580), 
        .C2(n1917), .ZN(n1918) );
  INV_X1 U1614 ( .A(n1920), .ZN(n1919) );
  INV_X1 U1615 ( .A(n1921), .ZN(n1916) );
  XNOR2_X1 U1616 ( .A(n1542), .B(n1922), .ZN(n772) );
  AOI221_X1 U1617 ( .B1(n1921), .B2(B[2]), .C1(n1920), .C2(B[1]), .A(n1923), 
        .ZN(n1922) );
  OAI22_X1 U1618 ( .A1(n1585), .A2(n1917), .B1(n1574), .B2(n1924), .ZN(n1923)
         );
  XNOR2_X1 U1619 ( .A(n1542), .B(n1925), .ZN(n771) );
  AOI221_X1 U1620 ( .B1(n1921), .B2(B[3]), .C1(n1920), .C2(B[2]), .A(n1926), 
        .ZN(n1925) );
  OAI22_X1 U1621 ( .A1(n1589), .A2(n1917), .B1(n1578), .B2(n1924), .ZN(n1926)
         );
  XNOR2_X1 U1622 ( .A(n1542), .B(n1927), .ZN(n770) );
  AOI221_X1 U1623 ( .B1(n1921), .B2(B[4]), .C1(n1920), .C2(B[3]), .A(n1928), 
        .ZN(n1927) );
  OAI22_X1 U1624 ( .A1(n1592), .A2(n1917), .B1(n1593), .B2(n1924), .ZN(n1928)
         );
  XNOR2_X1 U1625 ( .A(n1542), .B(n1929), .ZN(n769) );
  AOI221_X1 U1626 ( .B1(n1921), .B2(B[5]), .C1(n1920), .C2(B[4]), .A(n1930), 
        .ZN(n1929) );
  OAI22_X1 U1627 ( .A1(n1596), .A2(n1917), .B1(n1597), .B2(n1924), .ZN(n1930)
         );
  XNOR2_X1 U1628 ( .A(n1542), .B(n1931), .ZN(n768) );
  AOI221_X1 U1629 ( .B1(n1921), .B2(B[6]), .C1(n1920), .C2(B[5]), .A(n1932), 
        .ZN(n1931) );
  OAI22_X1 U1630 ( .A1(n1600), .A2(n1917), .B1(n1601), .B2(n1924), .ZN(n1932)
         );
  XNOR2_X1 U1631 ( .A(n1542), .B(n1933), .ZN(n767) );
  AOI221_X1 U1632 ( .B1(n1921), .B2(B[7]), .C1(n1920), .C2(B[6]), .A(n1934), 
        .ZN(n1933) );
  OAI22_X1 U1633 ( .A1(n1604), .A2(n1917), .B1(n1605), .B2(n1924), .ZN(n1934)
         );
  XNOR2_X1 U1634 ( .A(n1542), .B(n1935), .ZN(n766) );
  AOI221_X1 U1635 ( .B1(n1921), .B2(B[8]), .C1(n1920), .C2(B[7]), .A(n1936), 
        .ZN(n1935) );
  OAI22_X1 U1636 ( .A1(n1608), .A2(n1917), .B1(n1609), .B2(n1924), .ZN(n1936)
         );
  XNOR2_X1 U1637 ( .A(n1542), .B(n1937), .ZN(n765) );
  AOI221_X1 U1638 ( .B1(n1921), .B2(B[9]), .C1(n1920), .C2(B[8]), .A(n1938), 
        .ZN(n1937) );
  OAI22_X1 U1639 ( .A1(n1612), .A2(n1917), .B1(n1613), .B2(n1924), .ZN(n1938)
         );
  XNOR2_X1 U1640 ( .A(n1542), .B(n1939), .ZN(n764) );
  AOI221_X1 U1641 ( .B1(n1921), .B2(B[10]), .C1(n1920), .C2(B[9]), .A(n1940), 
        .ZN(n1939) );
  OAI22_X1 U1642 ( .A1(n1616), .A2(n1917), .B1(n1617), .B2(n1924), .ZN(n1940)
         );
  XNOR2_X1 U1643 ( .A(n1542), .B(n1941), .ZN(n763) );
  AOI221_X1 U1644 ( .B1(n1921), .B2(B[11]), .C1(n1920), .C2(B[10]), .A(n1942), 
        .ZN(n1941) );
  OAI22_X1 U1645 ( .A1(n1620), .A2(n1917), .B1(n1621), .B2(n1924), .ZN(n1942)
         );
  XNOR2_X1 U1646 ( .A(n1542), .B(n1943), .ZN(n762) );
  AOI221_X1 U1647 ( .B1(n1921), .B2(B[12]), .C1(n1920), .C2(B[11]), .A(n1944), 
        .ZN(n1943) );
  OAI22_X1 U1648 ( .A1(n1624), .A2(n1917), .B1(n1625), .B2(n1924), .ZN(n1944)
         );
  XNOR2_X1 U1649 ( .A(n1542), .B(n1945), .ZN(n761) );
  AOI221_X1 U1650 ( .B1(n1921), .B2(B[13]), .C1(n1920), .C2(B[12]), .A(n1946), 
        .ZN(n1945) );
  OAI22_X1 U1651 ( .A1(n1628), .A2(n1917), .B1(n1629), .B2(n1924), .ZN(n1946)
         );
  XNOR2_X1 U1652 ( .A(n1542), .B(n1947), .ZN(n760) );
  AOI221_X1 U1653 ( .B1(n1921), .B2(B[14]), .C1(n1920), .C2(B[13]), .A(n1948), 
        .ZN(n1947) );
  OAI22_X1 U1654 ( .A1(n1632), .A2(n1917), .B1(n1633), .B2(n1924), .ZN(n1948)
         );
  XNOR2_X1 U1655 ( .A(n1542), .B(n1949), .ZN(n759) );
  AOI221_X1 U1656 ( .B1(n1921), .B2(B[15]), .C1(n1920), .C2(B[14]), .A(n1950), 
        .ZN(n1949) );
  OAI22_X1 U1657 ( .A1(n1636), .A2(n1917), .B1(n1637), .B2(n1924), .ZN(n1950)
         );
  XNOR2_X1 U1658 ( .A(n1542), .B(n1951), .ZN(n758) );
  AOI221_X1 U1659 ( .B1(n1921), .B2(B[16]), .C1(n1920), .C2(B[15]), .A(n1952), 
        .ZN(n1951) );
  OAI22_X1 U1660 ( .A1(n1640), .A2(n1917), .B1(n1641), .B2(n1924), .ZN(n1952)
         );
  XNOR2_X1 U1661 ( .A(n1542), .B(n1953), .ZN(n757) );
  AOI221_X1 U1662 ( .B1(n1921), .B2(B[17]), .C1(n1920), .C2(B[16]), .A(n1954), 
        .ZN(n1953) );
  OAI22_X1 U1663 ( .A1(n1644), .A2(n1917), .B1(n1645), .B2(n1924), .ZN(n1954)
         );
  XNOR2_X1 U1664 ( .A(n1542), .B(n1955), .ZN(n756) );
  AOI221_X1 U1665 ( .B1(n1921), .B2(B[18]), .C1(n1920), .C2(B[17]), .A(n1956), 
        .ZN(n1955) );
  OAI22_X1 U1666 ( .A1(n1648), .A2(n1917), .B1(n1649), .B2(n1924), .ZN(n1956)
         );
  XNOR2_X1 U1667 ( .A(n1542), .B(n1957), .ZN(n755) );
  AOI221_X1 U1668 ( .B1(n1921), .B2(B[19]), .C1(n1920), .C2(B[18]), .A(n1958), 
        .ZN(n1957) );
  OAI22_X1 U1669 ( .A1(n1652), .A2(n1917), .B1(n1653), .B2(n1924), .ZN(n1958)
         );
  XNOR2_X1 U1670 ( .A(n1542), .B(n1959), .ZN(n754) );
  AOI221_X1 U1671 ( .B1(n1921), .B2(B[20]), .C1(n1920), .C2(B[19]), .A(n1960), 
        .ZN(n1959) );
  OAI22_X1 U1672 ( .A1(n1656), .A2(n1917), .B1(n1657), .B2(n1924), .ZN(n1960)
         );
  XNOR2_X1 U1673 ( .A(A[20]), .B(n1961), .ZN(n753) );
  AOI221_X1 U1674 ( .B1(n1921), .B2(B[21]), .C1(n1920), .C2(B[20]), .A(n1962), 
        .ZN(n1961) );
  OAI22_X1 U1675 ( .A1(n1660), .A2(n1917), .B1(n1661), .B2(n1924), .ZN(n1962)
         );
  XNOR2_X1 U1676 ( .A(A[20]), .B(n1963), .ZN(n752) );
  AOI221_X1 U1677 ( .B1(n1921), .B2(B[22]), .C1(n1920), .C2(B[21]), .A(n1964), 
        .ZN(n1963) );
  OAI22_X1 U1678 ( .A1(n1562), .A2(n1917), .B1(n1564), .B2(n1924), .ZN(n1964)
         );
  XNOR2_X1 U1679 ( .A(A[20]), .B(n1965), .ZN(n751) );
  AOI221_X1 U1680 ( .B1(n1921), .B2(n1554), .C1(n1920), .C2(B[22]), .A(n1966), 
        .ZN(n1965) );
  OAI22_X1 U1681 ( .A1(n1567), .A2(n1917), .B1(n1568), .B2(n1924), .ZN(n1966)
         );
  XNOR2_X1 U1682 ( .A(A[20]), .B(n1967), .ZN(n750) );
  AOI221_X1 U1683 ( .B1(n1921), .B2(B[23]), .C1(n1920), .C2(n1554), .A(n1968), 
        .ZN(n1967) );
  OAI22_X1 U1684 ( .A1(n1571), .A2(n1917), .B1(n1572), .B2(n1924), .ZN(n1968)
         );
  XNOR2_X1 U1685 ( .A(A[20]), .B(n1969), .ZN(n749) );
  OAI221_X1 U1686 ( .B1(n1556), .B2(n1924), .C1(n1556), .C2(n1917), .A(n1970), 
        .ZN(n1969) );
  OAI21_X1 U1687 ( .B1(n1921), .B2(n1920), .A(n1554), .ZN(n1970) );
  INV_X1 U1688 ( .A(n1974), .ZN(n1971) );
  XNOR2_X1 U1689 ( .A(A[18]), .B(A[19]), .ZN(n1972) );
  XNOR2_X1 U1690 ( .A(A[19]), .B(n1543), .ZN(n1973) );
  XOR2_X1 U1691 ( .A(A[18]), .B(n1545), .Z(n1974) );
  XNOR2_X1 U1692 ( .A(n1975), .B(n1541), .ZN(n748) );
  OAI22_X1 U1693 ( .A1(n1574), .A2(n1535), .B1(n1574), .B2(n1976), .ZN(n1975)
         );
  XNOR2_X1 U1694 ( .A(n1977), .B(n1541), .ZN(n747) );
  OAI222_X1 U1695 ( .A1(n1578), .A2(n1535), .B1(n1574), .B2(n1534), .C1(n1580), 
        .C2(n1976), .ZN(n1977) );
  INV_X1 U1696 ( .A(n1397), .ZN(n1580) );
  XNOR2_X1 U1697 ( .A(n1540), .B(n1978), .ZN(n746) );
  AOI221_X1 U1698 ( .B1(n1537), .B2(B[2]), .C1(n1536), .C2(B[1]), .A(n1979), 
        .ZN(n1978) );
  OAI22_X1 U1699 ( .A1(n1585), .A2(n1976), .B1(n1574), .B2(n1538), .ZN(n1979)
         );
  INV_X1 U1700 ( .A(n1396), .ZN(n1585) );
  XNOR2_X1 U1701 ( .A(n1540), .B(n1981), .ZN(n745) );
  AOI221_X1 U1702 ( .B1(n1537), .B2(B[3]), .C1(n1536), .C2(B[2]), .A(n1982), 
        .ZN(n1981) );
  OAI22_X1 U1703 ( .A1(n1589), .A2(n1976), .B1(n1578), .B2(n1539), .ZN(n1982)
         );
  XNOR2_X1 U1704 ( .A(n1540), .B(n1983), .ZN(n744) );
  AOI221_X1 U1705 ( .B1(n1537), .B2(B[4]), .C1(n1536), .C2(B[3]), .A(n1984), 
        .ZN(n1983) );
  OAI22_X1 U1706 ( .A1(n1592), .A2(n1976), .B1(n1593), .B2(n1539), .ZN(n1984)
         );
  XNOR2_X1 U1707 ( .A(n1540), .B(n1985), .ZN(n743) );
  AOI221_X1 U1708 ( .B1(n1537), .B2(B[5]), .C1(n1536), .C2(B[4]), .A(n1986), 
        .ZN(n1985) );
  OAI22_X1 U1709 ( .A1(n1596), .A2(n1976), .B1(n1597), .B2(n1539), .ZN(n1986)
         );
  XNOR2_X1 U1710 ( .A(n1540), .B(n1987), .ZN(n742) );
  AOI221_X1 U1711 ( .B1(n1537), .B2(B[6]), .C1(n1536), .C2(B[5]), .A(n1988), 
        .ZN(n1987) );
  OAI22_X1 U1712 ( .A1(n1600), .A2(n1976), .B1(n1601), .B2(n1539), .ZN(n1988)
         );
  XNOR2_X1 U1713 ( .A(n1540), .B(n1989), .ZN(n741) );
  AOI221_X1 U1714 ( .B1(n1537), .B2(B[7]), .C1(n1536), .C2(B[6]), .A(n1990), 
        .ZN(n1989) );
  OAI22_X1 U1715 ( .A1(n1604), .A2(n1976), .B1(n1605), .B2(n1539), .ZN(n1990)
         );
  XNOR2_X1 U1716 ( .A(n1540), .B(n1991), .ZN(n740) );
  AOI221_X1 U1717 ( .B1(n1537), .B2(B[9]), .C1(n1536), .C2(B[8]), .A(n1992), 
        .ZN(n1991) );
  OAI22_X1 U1718 ( .A1(n1612), .A2(n1976), .B1(n1613), .B2(n1539), .ZN(n1992)
         );
  XNOR2_X1 U1719 ( .A(n1540), .B(n1993), .ZN(n739) );
  AOI221_X1 U1720 ( .B1(n1537), .B2(B[10]), .C1(n1536), .C2(B[9]), .A(n1994), 
        .ZN(n1993) );
  OAI22_X1 U1721 ( .A1(n1616), .A2(n1976), .B1(n1617), .B2(n1539), .ZN(n1994)
         );
  XNOR2_X1 U1722 ( .A(n1540), .B(n1995), .ZN(n738) );
  AOI221_X1 U1723 ( .B1(n1537), .B2(B[12]), .C1(n1536), .C2(B[11]), .A(n1996), 
        .ZN(n1995) );
  OAI22_X1 U1724 ( .A1(n1624), .A2(n1976), .B1(n1625), .B2(n1539), .ZN(n1996)
         );
  XNOR2_X1 U1725 ( .A(n1540), .B(n1997), .ZN(n737) );
  AOI221_X1 U1726 ( .B1(n1537), .B2(B[13]), .C1(n1536), .C2(B[12]), .A(n1998), 
        .ZN(n1997) );
  OAI22_X1 U1727 ( .A1(n1628), .A2(n1976), .B1(n1629), .B2(n1539), .ZN(n1998)
         );
  XNOR2_X1 U1728 ( .A(n1540), .B(n1999), .ZN(n736) );
  AOI221_X1 U1729 ( .B1(n1537), .B2(B[14]), .C1(n1536), .C2(B[13]), .A(n2000), 
        .ZN(n1999) );
  OAI22_X1 U1730 ( .A1(n1632), .A2(n1976), .B1(n1633), .B2(n1539), .ZN(n2000)
         );
  XNOR2_X1 U1731 ( .A(n1540), .B(n2001), .ZN(n735) );
  AOI221_X1 U1732 ( .B1(n1537), .B2(B[15]), .C1(n1536), .C2(B[14]), .A(n2002), 
        .ZN(n2001) );
  OAI22_X1 U1733 ( .A1(n1636), .A2(n1976), .B1(n1637), .B2(n1539), .ZN(n2002)
         );
  XNOR2_X1 U1734 ( .A(n1540), .B(n2003), .ZN(n734) );
  AOI221_X1 U1735 ( .B1(n1537), .B2(B[16]), .C1(n1536), .C2(B[15]), .A(n2004), 
        .ZN(n2003) );
  OAI22_X1 U1736 ( .A1(n1640), .A2(n1976), .B1(n1641), .B2(n1538), .ZN(n2004)
         );
  XNOR2_X1 U1737 ( .A(n1540), .B(n2005), .ZN(n733) );
  AOI221_X1 U1738 ( .B1(n1537), .B2(B[18]), .C1(n1536), .C2(B[17]), .A(n2006), 
        .ZN(n2005) );
  OAI22_X1 U1739 ( .A1(n1648), .A2(n1976), .B1(n1649), .B2(n1538), .ZN(n2006)
         );
  XNOR2_X1 U1740 ( .A(n1540), .B(n2007), .ZN(n732) );
  AOI221_X1 U1741 ( .B1(n1537), .B2(B[19]), .C1(n1536), .C2(B[18]), .A(n2008), 
        .ZN(n2007) );
  OAI22_X1 U1742 ( .A1(n1652), .A2(n1976), .B1(n1653), .B2(n1538), .ZN(n2008)
         );
  XNOR2_X1 U1743 ( .A(n1540), .B(n2009), .ZN(n731) );
  AOI221_X1 U1744 ( .B1(n1537), .B2(B[20]), .C1(n1536), .C2(B[19]), .A(n2010), 
        .ZN(n2009) );
  OAI22_X1 U1745 ( .A1(n1656), .A2(n1976), .B1(n1657), .B2(n1538), .ZN(n2010)
         );
  XNOR2_X1 U1746 ( .A(A[23]), .B(n2011), .ZN(n730) );
  AOI221_X1 U1747 ( .B1(n1537), .B2(B[21]), .C1(n1536), .C2(B[20]), .A(n2012), 
        .ZN(n2011) );
  OAI22_X1 U1748 ( .A1(n1660), .A2(n1976), .B1(n1661), .B2(n1538), .ZN(n2012)
         );
  XNOR2_X1 U1749 ( .A(A[23]), .B(n2013), .ZN(n729) );
  AOI221_X1 U1750 ( .B1(n1537), .B2(B[22]), .C1(n1536), .C2(B[21]), .A(n2014), 
        .ZN(n2013) );
  OAI22_X1 U1751 ( .A1(n1562), .A2(n1976), .B1(n1564), .B2(n1538), .ZN(n2014)
         );
  INV_X1 U1752 ( .A(B[20]), .ZN(n1564) );
  INV_X1 U1753 ( .A(n1376), .ZN(n1562) );
  XNOR2_X1 U1754 ( .A(n519), .B(n2015), .ZN(n506) );
  INV_X1 U1755 ( .A(n493), .ZN(n479) );
  NOR2_X1 U1756 ( .A1(n2015), .A2(n519), .ZN(n493) );
  XOR2_X1 U1757 ( .A(n2016), .B(n1674), .Z(n2015) );
  OAI221_X1 U1758 ( .B1(n1563), .B2(n1556), .C1(n1561), .C2(n1556), .A(n2017), 
        .ZN(n2016) );
  OAI21_X1 U1759 ( .B1(n1558), .B2(n1559), .A(n1554), .ZN(n2017) );
  INV_X1 U1760 ( .A(n454), .ZN(n442) );
  XOR2_X1 U1761 ( .A(n1540), .B(n2018), .Z(n454) );
  AOI221_X1 U1762 ( .B1(n1537), .B2(B[8]), .C1(n1536), .C2(B[7]), .A(n2019), 
        .ZN(n2018) );
  OAI22_X1 U1763 ( .A1(n1608), .A2(n1976), .B1(n1609), .B2(n1538), .ZN(n2019)
         );
  INV_X1 U1764 ( .A(n421), .ZN(n411) );
  XOR2_X1 U1765 ( .A(n1540), .B(n2020), .Z(n421) );
  AOI221_X1 U1766 ( .B1(n1537), .B2(B[11]), .C1(n1536), .C2(B[10]), .A(n2021), 
        .ZN(n2020) );
  OAI22_X1 U1767 ( .A1(n1620), .A2(n1976), .B1(n1621), .B2(n1538), .ZN(n2021)
         );
  INV_X1 U1768 ( .A(n387), .ZN(n395) );
  INV_X1 U1769 ( .A(n374), .ZN(n368) );
  XOR2_X1 U1770 ( .A(n1540), .B(n2022), .Z(n374) );
  AOI221_X1 U1771 ( .B1(n1537), .B2(B[17]), .C1(n1536), .C2(B[16]), .A(n2023), 
        .ZN(n2022) );
  OAI22_X1 U1772 ( .A1(n1644), .A2(n1976), .B1(n1645), .B2(n1538), .ZN(n2023)
         );
  INV_X1 U1773 ( .A(n356), .ZN(n360) );
  INV_X1 U1774 ( .A(n2024), .ZN(n351) );
  OAI222_X1 U1775 ( .A1(n2025), .A2(n2026), .B1(n2025), .B2(n2027), .C1(n2027), 
        .C2(n2026), .ZN(n326) );
  INV_X1 U1776 ( .A(n550), .ZN(n2027) );
  XNOR2_X1 U1777 ( .A(n1674), .B(n2028), .ZN(n2026) );
  AOI221_X1 U1778 ( .B1(B[21]), .B2(n1558), .C1(B[20]), .C2(n1559), .A(n2029), 
        .ZN(n2028) );
  OAI22_X1 U1779 ( .A1(n1561), .A2(n1660), .B1(n1563), .B2(n1661), .ZN(n2029)
         );
  INV_X1 U1780 ( .A(B[19]), .ZN(n1661) );
  INV_X1 U1781 ( .A(n1377), .ZN(n1660) );
  AOI222_X1 U1782 ( .A1(n2030), .A2(n2031), .B1(n2030), .B2(n564), .C1(n564), 
        .C2(n2031), .ZN(n2025) );
  XNOR2_X1 U1783 ( .A(A[2]), .B(n2032), .ZN(n2031) );
  AOI221_X1 U1784 ( .B1(B[20]), .B2(n1558), .C1(B[19]), .C2(n1559), .A(n2033), 
        .ZN(n2032) );
  OAI22_X1 U1785 ( .A1(n1561), .A2(n1656), .B1(n1563), .B2(n1657), .ZN(n2033)
         );
  INV_X1 U1786 ( .A(B[18]), .ZN(n1657) );
  INV_X1 U1787 ( .A(n1378), .ZN(n1656) );
  INV_X1 U1788 ( .A(n2034), .ZN(n2030) );
  AOI222_X1 U1789 ( .A1(n2035), .A2(n2036), .B1(n2035), .B2(n576), .C1(n576), 
        .C2(n2036), .ZN(n2034) );
  XNOR2_X1 U1790 ( .A(A[2]), .B(n2037), .ZN(n2036) );
  AOI221_X1 U1791 ( .B1(B[19]), .B2(n1558), .C1(B[18]), .C2(n1559), .A(n2038), 
        .ZN(n2037) );
  OAI22_X1 U1792 ( .A1(n1561), .A2(n1652), .B1(n1563), .B2(n1653), .ZN(n2038)
         );
  INV_X1 U1793 ( .A(B[17]), .ZN(n1653) );
  INV_X1 U1794 ( .A(n1379), .ZN(n1652) );
  OAI222_X1 U1795 ( .A1(n2039), .A2(n2040), .B1(n2039), .B2(n2041), .C1(n2041), 
        .C2(n2040), .ZN(n2035) );
  INV_X1 U1796 ( .A(n588), .ZN(n2041) );
  XNOR2_X1 U1797 ( .A(n1674), .B(n2042), .ZN(n2040) );
  AOI221_X1 U1798 ( .B1(B[18]), .B2(n1558), .C1(B[17]), .C2(n1559), .A(n2043), 
        .ZN(n2042) );
  OAI22_X1 U1799 ( .A1(n1561), .A2(n1648), .B1(n1563), .B2(n1649), .ZN(n2043)
         );
  INV_X1 U1800 ( .A(B[16]), .ZN(n1649) );
  INV_X1 U1801 ( .A(n1380), .ZN(n1648) );
  AOI222_X1 U1802 ( .A1(n2044), .A2(n2045), .B1(n2044), .B2(n600), .C1(n600), 
        .C2(n2045), .ZN(n2039) );
  XNOR2_X1 U1803 ( .A(A[2]), .B(n2046), .ZN(n2045) );
  AOI221_X1 U1804 ( .B1(B[17]), .B2(n1558), .C1(B[16]), .C2(n1559), .A(n2047), 
        .ZN(n2046) );
  OAI22_X1 U1805 ( .A1(n1561), .A2(n1644), .B1(n1563), .B2(n1645), .ZN(n2047)
         );
  INV_X1 U1806 ( .A(B[15]), .ZN(n1645) );
  INV_X1 U1807 ( .A(n1381), .ZN(n1644) );
  OAI222_X1 U1808 ( .A1(n2048), .A2(n2049), .B1(n2048), .B2(n2050), .C1(n2050), 
        .C2(n2049), .ZN(n2044) );
  INV_X1 U1809 ( .A(n610), .ZN(n2050) );
  XNOR2_X1 U1810 ( .A(n1674), .B(n2051), .ZN(n2049) );
  AOI221_X1 U1811 ( .B1(B[16]), .B2(n1558), .C1(B[15]), .C2(n1559), .A(n2052), 
        .ZN(n2051) );
  OAI22_X1 U1812 ( .A1(n1561), .A2(n1640), .B1(n1563), .B2(n1641), .ZN(n2052)
         );
  INV_X1 U1813 ( .A(B[14]), .ZN(n1641) );
  INV_X1 U1814 ( .A(n1382), .ZN(n1640) );
  AOI222_X1 U1815 ( .A1(n2053), .A2(n2054), .B1(n2053), .B2(n620), .C1(n620), 
        .C2(n2054), .ZN(n2048) );
  XNOR2_X1 U1816 ( .A(A[2]), .B(n2055), .ZN(n2054) );
  AOI221_X1 U1817 ( .B1(B[15]), .B2(n1558), .C1(B[14]), .C2(n1559), .A(n2056), 
        .ZN(n2055) );
  OAI22_X1 U1818 ( .A1(n1561), .A2(n1636), .B1(n1563), .B2(n1637), .ZN(n2056)
         );
  INV_X1 U1819 ( .A(B[13]), .ZN(n1637) );
  INV_X1 U1820 ( .A(n1383), .ZN(n1636) );
  OAI222_X1 U1821 ( .A1(n2057), .A2(n2058), .B1(n2057), .B2(n2059), .C1(n2059), 
        .C2(n2058), .ZN(n2053) );
  INV_X1 U1822 ( .A(n630), .ZN(n2059) );
  XNOR2_X1 U1823 ( .A(n1674), .B(n2060), .ZN(n2058) );
  AOI221_X1 U1824 ( .B1(B[14]), .B2(n1558), .C1(B[13]), .C2(n1559), .A(n2061), 
        .ZN(n2060) );
  OAI22_X1 U1825 ( .A1(n1561), .A2(n1632), .B1(n1563), .B2(n1633), .ZN(n2061)
         );
  INV_X1 U1826 ( .A(B[12]), .ZN(n1633) );
  INV_X1 U1827 ( .A(n1384), .ZN(n1632) );
  AOI222_X1 U1828 ( .A1(n2062), .A2(n2063), .B1(n2062), .B2(n638), .C1(n638), 
        .C2(n2063), .ZN(n2057) );
  XNOR2_X1 U1829 ( .A(A[2]), .B(n2064), .ZN(n2063) );
  AOI221_X1 U1830 ( .B1(B[13]), .B2(n1558), .C1(B[12]), .C2(n1559), .A(n2065), 
        .ZN(n2064) );
  OAI22_X1 U1831 ( .A1(n1561), .A2(n1628), .B1(n1563), .B2(n1629), .ZN(n2065)
         );
  INV_X1 U1832 ( .A(B[11]), .ZN(n1629) );
  INV_X1 U1833 ( .A(n1385), .ZN(n1628) );
  OAI222_X1 U1834 ( .A1(n2066), .A2(n2067), .B1(n2066), .B2(n2068), .C1(n2068), 
        .C2(n2067), .ZN(n2062) );
  INV_X1 U1835 ( .A(n646), .ZN(n2068) );
  XNOR2_X1 U1836 ( .A(n1674), .B(n2069), .ZN(n2067) );
  AOI221_X1 U1837 ( .B1(B[12]), .B2(n1558), .C1(B[11]), .C2(n1559), .A(n2070), 
        .ZN(n2069) );
  OAI22_X1 U1838 ( .A1(n1561), .A2(n1624), .B1(n1563), .B2(n1625), .ZN(n2070)
         );
  INV_X1 U1839 ( .A(B[10]), .ZN(n1625) );
  INV_X1 U1840 ( .A(n1386), .ZN(n1624) );
  AOI222_X1 U1841 ( .A1(n2071), .A2(n2072), .B1(n2071), .B2(n654), .C1(n654), 
        .C2(n2072), .ZN(n2066) );
  XNOR2_X1 U1842 ( .A(A[2]), .B(n2073), .ZN(n2072) );
  AOI221_X1 U1843 ( .B1(B[11]), .B2(n1558), .C1(B[10]), .C2(n1559), .A(n2074), 
        .ZN(n2073) );
  OAI22_X1 U1844 ( .A1(n1561), .A2(n1620), .B1(n1563), .B2(n1621), .ZN(n2074)
         );
  INV_X1 U1845 ( .A(B[9]), .ZN(n1621) );
  INV_X1 U1846 ( .A(n1387), .ZN(n1620) );
  OAI222_X1 U1847 ( .A1(n2075), .A2(n2076), .B1(n2075), .B2(n2077), .C1(n2077), 
        .C2(n2076), .ZN(n2071) );
  INV_X1 U1848 ( .A(n660), .ZN(n2077) );
  XNOR2_X1 U1849 ( .A(n1674), .B(n2078), .ZN(n2076) );
  AOI221_X1 U1850 ( .B1(B[10]), .B2(n1558), .C1(B[9]), .C2(n1559), .A(n2079), 
        .ZN(n2078) );
  OAI22_X1 U1851 ( .A1(n1561), .A2(n1616), .B1(n1563), .B2(n1617), .ZN(n2079)
         );
  INV_X1 U1852 ( .A(B[8]), .ZN(n1617) );
  INV_X1 U1853 ( .A(n1388), .ZN(n1616) );
  AOI222_X1 U1854 ( .A1(n2080), .A2(n2081), .B1(n2080), .B2(n666), .C1(n666), 
        .C2(n2081), .ZN(n2075) );
  XNOR2_X1 U1855 ( .A(A[2]), .B(n2082), .ZN(n2081) );
  AOI221_X1 U1856 ( .B1(B[9]), .B2(n1558), .C1(B[8]), .C2(n1559), .A(n2083), 
        .ZN(n2082) );
  OAI22_X1 U1857 ( .A1(n1561), .A2(n1612), .B1(n1563), .B2(n1613), .ZN(n2083)
         );
  INV_X1 U1858 ( .A(B[7]), .ZN(n1613) );
  INV_X1 U1859 ( .A(n1389), .ZN(n1612) );
  OAI222_X1 U1860 ( .A1(n2084), .A2(n2085), .B1(n2084), .B2(n2086), .C1(n2086), 
        .C2(n2085), .ZN(n2080) );
  INV_X1 U1861 ( .A(n672), .ZN(n2086) );
  XNOR2_X1 U1862 ( .A(n1674), .B(n2087), .ZN(n2085) );
  AOI221_X1 U1863 ( .B1(B[8]), .B2(n1558), .C1(B[7]), .C2(n1559), .A(n2088), 
        .ZN(n2087) );
  OAI22_X1 U1864 ( .A1(n1561), .A2(n1608), .B1(n1563), .B2(n1609), .ZN(n2088)
         );
  INV_X1 U1865 ( .A(B[6]), .ZN(n1609) );
  INV_X1 U1866 ( .A(n1390), .ZN(n1608) );
  AOI222_X1 U1867 ( .A1(n2089), .A2(n2090), .B1(n2089), .B2(n676), .C1(n676), 
        .C2(n2090), .ZN(n2084) );
  XNOR2_X1 U1868 ( .A(A[2]), .B(n2091), .ZN(n2090) );
  AOI221_X1 U1869 ( .B1(B[7]), .B2(n1558), .C1(B[6]), .C2(n1559), .A(n2092), 
        .ZN(n2091) );
  OAI22_X1 U1870 ( .A1(n1561), .A2(n1604), .B1(n1563), .B2(n1605), .ZN(n2092)
         );
  INV_X1 U1871 ( .A(B[5]), .ZN(n1605) );
  INV_X1 U1872 ( .A(n1391), .ZN(n1604) );
  OAI222_X1 U1873 ( .A1(n2093), .A2(n2094), .B1(n2093), .B2(n2095), .C1(n2095), 
        .C2(n2094), .ZN(n2089) );
  INV_X1 U1874 ( .A(n680), .ZN(n2095) );
  XNOR2_X1 U1875 ( .A(n1674), .B(n2096), .ZN(n2094) );
  AOI221_X1 U1876 ( .B1(B[6]), .B2(n1558), .C1(B[5]), .C2(n1559), .A(n2097), 
        .ZN(n2096) );
  OAI22_X1 U1877 ( .A1(n1561), .A2(n1600), .B1(n1563), .B2(n1601), .ZN(n2097)
         );
  INV_X1 U1878 ( .A(B[4]), .ZN(n1601) );
  INV_X1 U1879 ( .A(n1392), .ZN(n1600) );
  AOI222_X1 U1880 ( .A1(n2098), .A2(n2099), .B1(n2098), .B2(n684), .C1(n684), 
        .C2(n2099), .ZN(n2093) );
  XNOR2_X1 U1881 ( .A(A[2]), .B(n2100), .ZN(n2099) );
  AOI221_X1 U1882 ( .B1(B[5]), .B2(n1558), .C1(B[4]), .C2(n1559), .A(n2101), 
        .ZN(n2100) );
  OAI22_X1 U1883 ( .A1(n1561), .A2(n1596), .B1(n1563), .B2(n1597), .ZN(n2101)
         );
  INV_X1 U1884 ( .A(B[3]), .ZN(n1597) );
  INV_X1 U1885 ( .A(n1393), .ZN(n1596) );
  OAI222_X1 U1886 ( .A1(n2102), .A2(n2103), .B1(n2102), .B2(n2104), .C1(n2104), 
        .C2(n2103), .ZN(n2098) );
  INV_X1 U1887 ( .A(n686), .ZN(n2104) );
  XNOR2_X1 U1888 ( .A(n1674), .B(n2105), .ZN(n2103) );
  AOI221_X1 U1889 ( .B1(B[4]), .B2(n1558), .C1(B[3]), .C2(n1559), .A(n2106), 
        .ZN(n2105) );
  OAI22_X1 U1890 ( .A1(n1561), .A2(n1592), .B1(n1563), .B2(n1593), .ZN(n2106)
         );
  INV_X1 U1891 ( .A(B[2]), .ZN(n1593) );
  INV_X1 U1892 ( .A(n1394), .ZN(n1592) );
  AOI222_X1 U1893 ( .A1(n2107), .A2(n2108), .B1(n2107), .B2(n688), .C1(n688), 
        .C2(n2108), .ZN(n2102) );
  XNOR2_X1 U1894 ( .A(A[2]), .B(n2109), .ZN(n2108) );
  AOI221_X1 U1895 ( .B1(B[3]), .B2(n1558), .C1(B[2]), .C2(n1559), .A(n2110), 
        .ZN(n2109) );
  OAI22_X1 U1896 ( .A1(n1561), .A2(n1589), .B1(n1563), .B2(n1578), .ZN(n2110)
         );
  INV_X1 U1897 ( .A(B[1]), .ZN(n1578) );
  INV_X1 U1898 ( .A(n1395), .ZN(n1589) );
  AND2_X1 U1899 ( .A1(n2114), .A2(n2115), .ZN(n2107) );
  AOI211_X1 U1900 ( .C1(B[1]), .C2(n1558), .A(n2116), .B(B[0]), .ZN(n2115) );
  INV_X1 U1901 ( .A(n2117), .ZN(n2116) );
  AOI22_X1 U1902 ( .A1(n1558), .A2(B[2]), .B1(n2118), .B2(n1397), .ZN(n2117)
         );
  INV_X1 U1903 ( .A(A[0]), .ZN(n2112) );
  AOI221_X1 U1904 ( .B1(B[1]), .B2(n1559), .C1(n1396), .C2(n2118), .A(n1674), 
        .ZN(n2114) );
  INV_X1 U1905 ( .A(n1561), .ZN(n2118) );
  XNOR2_X1 U1906 ( .A(A[1]), .B(n1674), .ZN(n2111) );
  INV_X1 U1907 ( .A(A[2]), .ZN(n1674) );
  INV_X1 U1908 ( .A(A[1]), .ZN(n2113) );
  AOI21_X1 U1909 ( .B1(n2119), .B2(n2120), .A(n2121), .ZN(PRODUCT[47]) );
  OAI22_X1 U1910 ( .A1(n2122), .A2(n2123), .B1(n2122), .B2(n2124), .ZN(n2121)
         );
  INV_X1 U1911 ( .A(n2120), .ZN(n2124) );
  AOI222_X1 U1912 ( .A1(n2024), .A2(n303), .B1(n2123), .B2(n303), .C1(n2024), 
        .C2(n2123), .ZN(n2122) );
  XOR2_X1 U1913 ( .A(n1541), .B(n2125), .Z(n2024) );
  AOI221_X1 U1914 ( .B1(n1537), .B2(B[23]), .C1(n1536), .C2(B[22]), .A(n2126), 
        .ZN(n2125) );
  OAI22_X1 U1915 ( .A1(n1567), .A2(n1976), .B1(n1568), .B2(n1538), .ZN(n2126)
         );
  INV_X1 U1916 ( .A(B[21]), .ZN(n1568) );
  INV_X1 U1917 ( .A(n1375), .ZN(n1567) );
  XOR2_X1 U1918 ( .A(n2127), .B(n1541), .Z(n2120) );
  OAI221_X1 U1919 ( .B1(n1556), .B2(n1539), .C1(n1556), .C2(n1976), .A(n2128), 
        .ZN(n2127) );
  OAI21_X1 U1920 ( .B1(n1537), .B2(n1536), .A(n1554), .ZN(n2128) );
  INV_X1 U1921 ( .A(n2123), .ZN(n2119) );
  XOR2_X1 U1922 ( .A(A[23]), .B(n2129), .Z(n2123) );
  AOI221_X1 U1923 ( .B1(n1537), .B2(n1554), .C1(n1536), .C2(n1554), .A(n2130), 
        .ZN(n2129) );
  OAI22_X1 U1924 ( .A1(n1571), .A2(n1976), .B1(n1572), .B2(n1538), .ZN(n2130)
         );
  NAND3_X1 U1925 ( .A1(n2131), .A2(n2132), .A3(n2133), .ZN(n1980) );
  INV_X1 U1926 ( .A(B[22]), .ZN(n1572) );
  INV_X1 U1927 ( .A(n1374), .ZN(n1571) );
  XNOR2_X1 U1928 ( .A(A[21]), .B(A[22]), .ZN(n2133) );
  INV_X1 U1929 ( .A(n2131), .ZN(n2134) );
  XOR2_X1 U1930 ( .A(A[21]), .B(n1543), .Z(n2131) );
  XNOR2_X1 U1931 ( .A(A[22]), .B(n1541), .ZN(n2132) );
endmodule


module iir_filter_DW02_mult_3 ( A, B, PRODUCT, TC );
  input [23:0] A;
  input [23:0] B;
  output [47:0] PRODUCT;
  input TC;
  wire   n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n351, n352, n353, n354, n355, n356, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n906, n907, n908, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134;

  FA_X1 U182 ( .A(n351), .B(n352), .CI(n304), .CO(n303), .S(PRODUCT[44]) );
  FA_X1 U183 ( .A(n353), .B(n354), .CI(n305), .CO(n304), .S(PRODUCT[43]) );
  FA_X1 U184 ( .A(n355), .B(n358), .CI(n306), .CO(n305), .S(PRODUCT[42]) );
  FA_X1 U185 ( .A(n359), .B(n361), .CI(n307), .CO(n306), .S(PRODUCT[41]) );
  FA_X1 U186 ( .A(n362), .B(n364), .CI(n308), .CO(n307), .S(PRODUCT[40]) );
  FA_X1 U187 ( .A(n365), .B(n370), .CI(n309), .CO(n308), .S(PRODUCT[39]) );
  FA_X1 U188 ( .A(n371), .B(n375), .CI(n310), .CO(n309), .S(PRODUCT[38]) );
  FA_X1 U189 ( .A(n376), .B(n381), .CI(n311), .CO(n310), .S(PRODUCT[37]) );
  FA_X1 U190 ( .A(n382), .B(n389), .CI(n312), .CO(n311), .S(PRODUCT[36]) );
  FA_X1 U191 ( .A(n390), .B(n396), .CI(n313), .CO(n312), .S(PRODUCT[35]) );
  FA_X1 U192 ( .A(n397), .B(n403), .CI(n314), .CO(n313), .S(PRODUCT[34]) );
  FA_X1 U193 ( .A(n404), .B(n413), .CI(n315), .CO(n314), .S(PRODUCT[33]) );
  FA_X1 U194 ( .A(n414), .B(n422), .CI(n316), .CO(n315), .S(PRODUCT[32]) );
  FA_X1 U195 ( .A(n423), .B(n432), .CI(n317), .CO(n316), .S(PRODUCT[31]) );
  FA_X1 U196 ( .A(n433), .B(n444), .CI(n318), .CO(n317), .S(PRODUCT[30]) );
  FA_X1 U197 ( .A(n445), .B(n455), .CI(n319), .CO(n318), .S(PRODUCT[29]) );
  FA_X1 U198 ( .A(n456), .B(n467), .CI(n320), .CO(n319), .S(PRODUCT[28]) );
  FA_X1 U199 ( .A(n468), .B(n481), .CI(n321), .CO(n320), .S(PRODUCT[27]) );
  FA_X1 U200 ( .A(n482), .B(n494), .CI(n322), .CO(n321), .S(PRODUCT[26]) );
  FA_X1 U201 ( .A(n495), .B(n507), .CI(n323), .CO(n322), .S(PRODUCT[25]) );
  FA_X1 U202 ( .A(n508), .B(n906), .CI(n324), .CO(n323), .S(PRODUCT[24]) );
  FA_X1 U203 ( .A(n907), .B(n522), .CI(n325), .CO(n324), .S(PRODUCT[23]) );
  FA_X1 U204 ( .A(n908), .B(n536), .CI(n326), .CO(n325), .S(PRODUCT[22]) );
  FA_X1 U235 ( .A(n356), .B(n749), .CI(n729), .CO(n352), .S(n353) );
  FA_X1 U236 ( .A(n730), .B(n360), .CI(n750), .CO(n354), .S(n355) );
  FA_X1 U238 ( .A(n360), .B(n731), .CI(n751), .CO(n358), .S(n359) );
  FA_X1 U240 ( .A(n752), .B(n363), .CI(n366), .CO(n361), .S(n362) );
  FA_X1 U241 ( .A(n368), .B(n775), .CI(n732), .CO(n356), .S(n363) );
  FA_X1 U242 ( .A(n776), .B(n753), .CI(n367), .CO(n364), .S(n365) );
  FA_X1 U243 ( .A(n733), .B(n374), .CI(n372), .CO(n366), .S(n367) );
  FA_X1 U245 ( .A(n373), .B(n377), .CI(n777), .CO(n370), .S(n371) );
  FA_X1 U246 ( .A(n374), .B(n379), .CI(n754), .CO(n372), .S(n373) );
  FA_X1 U248 ( .A(n778), .B(n378), .CI(n383), .CO(n375), .S(n376) );
  FA_X1 U249 ( .A(n385), .B(n380), .CI(n755), .CO(n377), .S(n378) );
  FA_X1 U250 ( .A(n387), .B(n801), .CI(n734), .CO(n379), .S(n380) );
  FA_X1 U251 ( .A(n802), .B(n779), .CI(n384), .CO(n381), .S(n382) );
  FA_X1 U252 ( .A(n386), .B(n393), .CI(n391), .CO(n383), .S(n384) );
  FA_X1 U253 ( .A(n735), .B(n395), .CI(n756), .CO(n385), .S(n386) );
  FA_X1 U255 ( .A(n392), .B(n398), .CI(n803), .CO(n389), .S(n390) );
  FA_X1 U256 ( .A(n394), .B(n400), .CI(n780), .CO(n391), .S(n392) );
  FA_X1 U257 ( .A(n395), .B(n736), .CI(n757), .CO(n393), .S(n394) );
  FA_X1 U259 ( .A(n804), .B(n399), .CI(n405), .CO(n396), .S(n397) );
  FA_X1 U260 ( .A(n407), .B(n401), .CI(n781), .CO(n398), .S(n399) );
  FA_X1 U261 ( .A(n758), .B(n402), .CI(n409), .CO(n400), .S(n401) );
  FA_X1 U262 ( .A(n411), .B(n827), .CI(n737), .CO(n387), .S(n402) );
  FA_X1 U263 ( .A(n828), .B(n805), .CI(n406), .CO(n403), .S(n404) );
  FA_X1 U264 ( .A(n408), .B(n417), .CI(n415), .CO(n405), .S(n406) );
  FA_X1 U265 ( .A(n410), .B(n759), .CI(n782), .CO(n407), .S(n408) );
  FA_X1 U266 ( .A(n738), .B(n421), .CI(n419), .CO(n409), .S(n410) );
  FA_X1 U268 ( .A(n416), .B(n424), .CI(n829), .CO(n413), .S(n414) );
  FA_X1 U269 ( .A(n418), .B(n426), .CI(n806), .CO(n415), .S(n416) );
  FA_X1 U270 ( .A(n420), .B(n428), .CI(n783), .CO(n417), .S(n418) );
  FA_X1 U271 ( .A(n421), .B(n430), .CI(n760), .CO(n419), .S(n420) );
  FA_X1 U273 ( .A(n830), .B(n425), .CI(n434), .CO(n422), .S(n423) );
  FA_X1 U274 ( .A(n436), .B(n427), .CI(n807), .CO(n424), .S(n425) );
  FA_X1 U275 ( .A(n784), .B(n429), .CI(n438), .CO(n426), .S(n427) );
  FA_X1 U276 ( .A(n440), .B(n431), .CI(n761), .CO(n428), .S(n429) );
  FA_X1 U277 ( .A(n442), .B(n853), .CI(n739), .CO(n430), .S(n431) );
  FA_X1 U278 ( .A(n854), .B(n831), .CI(n435), .CO(n432), .S(n433) );
  FA_X1 U279 ( .A(n437), .B(n448), .CI(n446), .CO(n434), .S(n435) );
  FA_X1 U280 ( .A(n439), .B(n785), .CI(n808), .CO(n436), .S(n437) );
  FA_X1 U281 ( .A(n441), .B(n452), .CI(n450), .CO(n438), .S(n439) );
  FA_X1 U282 ( .A(n740), .B(n454), .CI(n762), .CO(n440), .S(n441) );
  FA_X1 U284 ( .A(n447), .B(n457), .CI(n855), .CO(n444), .S(n445) );
  FA_X1 U285 ( .A(n449), .B(n459), .CI(n832), .CO(n446), .S(n447) );
  FA_X1 U286 ( .A(n451), .B(n461), .CI(n809), .CO(n448), .S(n449) );
  FA_X1 U287 ( .A(n453), .B(n463), .CI(n786), .CO(n450), .S(n451) );
  FA_X1 U288 ( .A(n454), .B(n465), .CI(n763), .CO(n452), .S(n453) );
  FA_X1 U290 ( .A(n856), .B(n458), .CI(n469), .CO(n455), .S(n456) );
  FA_X1 U291 ( .A(n471), .B(n460), .CI(n833), .CO(n457), .S(n458) );
  FA_X1 U292 ( .A(n810), .B(n462), .CI(n473), .CO(n459), .S(n460) );
  FA_X1 U293 ( .A(n475), .B(n464), .CI(n787), .CO(n461), .S(n462) );
  FA_X1 U294 ( .A(n764), .B(n466), .CI(n477), .CO(n463), .S(n464) );
  FA_X1 U295 ( .A(n479), .B(n879), .CI(n741), .CO(n465), .S(n466) );
  FA_X1 U296 ( .A(n880), .B(n857), .CI(n470), .CO(n467), .S(n468) );
  FA_X1 U297 ( .A(n472), .B(n485), .CI(n483), .CO(n469), .S(n470) );
  FA_X1 U298 ( .A(n474), .B(n811), .CI(n834), .CO(n471), .S(n472) );
  FA_X1 U299 ( .A(n476), .B(n489), .CI(n487), .CO(n473), .S(n474) );
  FA_X1 U300 ( .A(n478), .B(n765), .CI(n788), .CO(n475), .S(n476) );
  FA_X1 U301 ( .A(n742), .B(n493), .CI(n491), .CO(n477), .S(n478) );
  FA_X1 U303 ( .A(n484), .B(n858), .CI(n881), .CO(n481), .S(n482) );
  FA_X1 U304 ( .A(n486), .B(n498), .CI(n496), .CO(n483), .S(n484) );
  FA_X1 U305 ( .A(n488), .B(n812), .CI(n835), .CO(n485), .S(n486) );
  FA_X1 U306 ( .A(n490), .B(n502), .CI(n500), .CO(n487), .S(n488) );
  FA_X1 U307 ( .A(n492), .B(n504), .CI(n789), .CO(n489), .S(n490) );
  FA_X1 U308 ( .A(n743), .B(n493), .CI(n766), .CO(n491), .S(n492) );
  FA_X1 U310 ( .A(n497), .B(n509), .CI(n882), .CO(n494), .S(n495) );
  FA_X1 U311 ( .A(n499), .B(n511), .CI(n859), .CO(n496), .S(n497) );
  FA_X1 U312 ( .A(n501), .B(n513), .CI(n836), .CO(n498), .S(n499) );
  FA_X1 U313 ( .A(n503), .B(n515), .CI(n813), .CO(n500), .S(n501) );
  FA_X1 U314 ( .A(n505), .B(n517), .CI(n790), .CO(n502), .S(n503) );
  FA_X1 U315 ( .A(n506), .B(n744), .CI(n767), .CO(n504), .S(n505) );
  FA_X1 U318 ( .A(n883), .B(n510), .CI(n521), .CO(n507), .S(n508) );
  FA_X1 U319 ( .A(n860), .B(n512), .CI(n523), .CO(n509), .S(n510) );
  FA_X1 U320 ( .A(n837), .B(n514), .CI(n525), .CO(n511), .S(n512) );
  FA_X1 U321 ( .A(n814), .B(n516), .CI(n527), .CO(n513), .S(n514) );
  FA_X1 U322 ( .A(n791), .B(n518), .CI(n529), .CO(n515), .S(n516) );
  FA_X1 U323 ( .A(n768), .B(n520), .CI(n531), .CO(n517), .S(n518) );
  HA_X1 U324 ( .A(n533), .B(n745), .CO(n519), .S(n520) );
  FA_X1 U325 ( .A(n884), .B(n524), .CI(n535), .CO(n521), .S(n522) );
  FA_X1 U326 ( .A(n861), .B(n526), .CI(n537), .CO(n523), .S(n524) );
  FA_X1 U327 ( .A(n838), .B(n528), .CI(n539), .CO(n525), .S(n526) );
  FA_X1 U328 ( .A(n815), .B(n530), .CI(n541), .CO(n527), .S(n528) );
  FA_X1 U329 ( .A(n792), .B(n532), .CI(n543), .CO(n529), .S(n530) );
  FA_X1 U330 ( .A(n769), .B(n534), .CI(n545), .CO(n531), .S(n532) );
  HA_X1 U331 ( .A(n547), .B(n746), .CO(n533), .S(n534) );
  FA_X1 U332 ( .A(n885), .B(n538), .CI(n549), .CO(n535), .S(n536) );
  FA_X1 U333 ( .A(n862), .B(n540), .CI(n551), .CO(n537), .S(n538) );
  FA_X1 U334 ( .A(n839), .B(n542), .CI(n553), .CO(n539), .S(n540) );
  FA_X1 U335 ( .A(n816), .B(n544), .CI(n555), .CO(n541), .S(n542) );
  FA_X1 U336 ( .A(n793), .B(n546), .CI(n557), .CO(n543), .S(n544) );
  FA_X1 U337 ( .A(n770), .B(n548), .CI(n559), .CO(n545), .S(n546) );
  HA_X1 U338 ( .A(n561), .B(n747), .CO(n547), .S(n548) );
  FA_X1 U339 ( .A(n886), .B(n552), .CI(n563), .CO(n549), .S(n550) );
  FA_X1 U340 ( .A(n863), .B(n554), .CI(n565), .CO(n551), .S(n552) );
  FA_X1 U341 ( .A(n840), .B(n556), .CI(n567), .CO(n553), .S(n554) );
  FA_X1 U342 ( .A(n817), .B(n558), .CI(n569), .CO(n555), .S(n556) );
  FA_X1 U343 ( .A(n794), .B(n560), .CI(n571), .CO(n557), .S(n558) );
  FA_X1 U344 ( .A(n771), .B(n562), .CI(n573), .CO(n559), .S(n560) );
  HA_X1 U345 ( .A(n748), .B(n1540), .CO(n561), .S(n562) );
  FA_X1 U346 ( .A(n887), .B(n566), .CI(n575), .CO(n563), .S(n564) );
  FA_X1 U347 ( .A(n864), .B(n568), .CI(n577), .CO(n565), .S(n566) );
  FA_X1 U348 ( .A(n841), .B(n570), .CI(n579), .CO(n567), .S(n568) );
  FA_X1 U349 ( .A(n818), .B(n572), .CI(n581), .CO(n569), .S(n570) );
  FA_X1 U350 ( .A(n795), .B(n574), .CI(n583), .CO(n571), .S(n572) );
  HA_X1 U351 ( .A(n585), .B(n772), .CO(n573), .S(n574) );
  FA_X1 U352 ( .A(n888), .B(n578), .CI(n587), .CO(n575), .S(n576) );
  FA_X1 U353 ( .A(n865), .B(n580), .CI(n589), .CO(n577), .S(n578) );
  FA_X1 U354 ( .A(n842), .B(n582), .CI(n591), .CO(n579), .S(n580) );
  FA_X1 U355 ( .A(n819), .B(n584), .CI(n593), .CO(n581), .S(n582) );
  FA_X1 U356 ( .A(n796), .B(n586), .CI(n595), .CO(n583), .S(n584) );
  HA_X1 U357 ( .A(n597), .B(n773), .CO(n585), .S(n586) );
  FA_X1 U358 ( .A(n889), .B(n590), .CI(n599), .CO(n587), .S(n588) );
  FA_X1 U359 ( .A(n866), .B(n592), .CI(n601), .CO(n589), .S(n590) );
  FA_X1 U360 ( .A(n843), .B(n594), .CI(n603), .CO(n591), .S(n592) );
  FA_X1 U361 ( .A(n820), .B(n596), .CI(n605), .CO(n593), .S(n594) );
  FA_X1 U362 ( .A(n797), .B(n598), .CI(n607), .CO(n595), .S(n596) );
  HA_X1 U363 ( .A(n774), .B(n1542), .CO(n597), .S(n598) );
  FA_X1 U364 ( .A(n890), .B(n602), .CI(n609), .CO(n599), .S(n600) );
  FA_X1 U365 ( .A(n867), .B(n604), .CI(n611), .CO(n601), .S(n602) );
  FA_X1 U366 ( .A(n844), .B(n606), .CI(n613), .CO(n603), .S(n604) );
  FA_X1 U367 ( .A(n821), .B(n608), .CI(n615), .CO(n605), .S(n606) );
  HA_X1 U368 ( .A(n617), .B(n798), .CO(n607), .S(n608) );
  FA_X1 U369 ( .A(n891), .B(n612), .CI(n619), .CO(n609), .S(n610) );
  FA_X1 U370 ( .A(n868), .B(n614), .CI(n621), .CO(n611), .S(n612) );
  FA_X1 U371 ( .A(n845), .B(n616), .CI(n623), .CO(n613), .S(n614) );
  FA_X1 U372 ( .A(n822), .B(n618), .CI(n625), .CO(n615), .S(n616) );
  HA_X1 U373 ( .A(n627), .B(n799), .CO(n617), .S(n618) );
  FA_X1 U374 ( .A(n892), .B(n622), .CI(n629), .CO(n619), .S(n620) );
  FA_X1 U375 ( .A(n869), .B(n624), .CI(n631), .CO(n621), .S(n622) );
  FA_X1 U376 ( .A(n846), .B(n626), .CI(n633), .CO(n623), .S(n624) );
  FA_X1 U377 ( .A(n823), .B(n628), .CI(n635), .CO(n625), .S(n626) );
  HA_X1 U378 ( .A(n800), .B(n1544), .CO(n627), .S(n628) );
  FA_X1 U379 ( .A(n893), .B(n632), .CI(n637), .CO(n629), .S(n630) );
  FA_X1 U380 ( .A(n870), .B(n634), .CI(n639), .CO(n631), .S(n632) );
  FA_X1 U381 ( .A(n847), .B(n636), .CI(n641), .CO(n633), .S(n634) );
  HA_X1 U382 ( .A(n643), .B(n824), .CO(n635), .S(n636) );
  FA_X1 U383 ( .A(n894), .B(n640), .CI(n645), .CO(n637), .S(n638) );
  FA_X1 U384 ( .A(n871), .B(n642), .CI(n647), .CO(n639), .S(n640) );
  FA_X1 U385 ( .A(n848), .B(n644), .CI(n649), .CO(n641), .S(n642) );
  HA_X1 U386 ( .A(n651), .B(n825), .CO(n643), .S(n644) );
  FA_X1 U387 ( .A(n895), .B(n648), .CI(n653), .CO(n645), .S(n646) );
  FA_X1 U388 ( .A(n872), .B(n650), .CI(n655), .CO(n647), .S(n648) );
  FA_X1 U389 ( .A(n849), .B(n652), .CI(n657), .CO(n649), .S(n650) );
  HA_X1 U390 ( .A(n826), .B(n1546), .CO(n651), .S(n652) );
  FA_X1 U391 ( .A(n896), .B(n656), .CI(n659), .CO(n653), .S(n654) );
  FA_X1 U392 ( .A(n873), .B(n658), .CI(n661), .CO(n655), .S(n656) );
  HA_X1 U393 ( .A(n663), .B(n850), .CO(n657), .S(n658) );
  FA_X1 U394 ( .A(n897), .B(n662), .CI(n665), .CO(n659), .S(n660) );
  FA_X1 U395 ( .A(n874), .B(n664), .CI(n667), .CO(n661), .S(n662) );
  HA_X1 U396 ( .A(n669), .B(n851), .CO(n663), .S(n664) );
  FA_X1 U397 ( .A(n898), .B(n668), .CI(n671), .CO(n665), .S(n666) );
  FA_X1 U398 ( .A(n875), .B(n670), .CI(n673), .CO(n667), .S(n668) );
  HA_X1 U399 ( .A(n852), .B(n1548), .CO(n669), .S(n670) );
  FA_X1 U400 ( .A(n899), .B(n674), .CI(n675), .CO(n671), .S(n672) );
  HA_X1 U401 ( .A(n677), .B(n876), .CO(n673), .S(n674) );
  FA_X1 U402 ( .A(n900), .B(n678), .CI(n679), .CO(n675), .S(n676) );
  HA_X1 U403 ( .A(n681), .B(n877), .CO(n677), .S(n678) );
  FA_X1 U404 ( .A(n901), .B(n682), .CI(n683), .CO(n679), .S(n680) );
  HA_X1 U405 ( .A(n878), .B(n1550), .CO(n681), .S(n682) );
  HA_X1 U406 ( .A(n685), .B(n902), .CO(n683), .S(n684) );
  HA_X1 U407 ( .A(n687), .B(n903), .CO(n685), .S(n686) );
  HA_X1 U408 ( .A(n904), .B(n1552), .CO(n687), .S(n688) );
  FA_X1 U1112 ( .A(B[22]), .B(n1554), .CI(n706), .CO(n1374), .S(n1375) );
  FA_X1 U1113 ( .A(B[21]), .B(B[22]), .CI(n707), .CO(n706), .S(n1376) );
  FA_X1 U1114 ( .A(B[20]), .B(B[21]), .CI(n708), .CO(n707), .S(n1377) );
  FA_X1 U1115 ( .A(B[19]), .B(B[20]), .CI(n709), .CO(n708), .S(n1378) );
  FA_X1 U1116 ( .A(B[18]), .B(B[19]), .CI(n710), .CO(n709), .S(n1379) );
  FA_X1 U1117 ( .A(B[17]), .B(B[18]), .CI(n711), .CO(n710), .S(n1380) );
  FA_X1 U1118 ( .A(B[16]), .B(B[17]), .CI(n712), .CO(n711), .S(n1381) );
  FA_X1 U1119 ( .A(B[15]), .B(B[16]), .CI(n713), .CO(n712), .S(n1382) );
  FA_X1 U1120 ( .A(B[14]), .B(B[15]), .CI(n714), .CO(n713), .S(n1383) );
  FA_X1 U1121 ( .A(B[13]), .B(B[14]), .CI(n715), .CO(n714), .S(n1384) );
  FA_X1 U1122 ( .A(B[12]), .B(B[13]), .CI(n716), .CO(n715), .S(n1385) );
  FA_X1 U1123 ( .A(B[11]), .B(B[12]), .CI(n717), .CO(n716), .S(n1386) );
  FA_X1 U1124 ( .A(B[10]), .B(B[11]), .CI(n718), .CO(n717), .S(n1387) );
  FA_X1 U1125 ( .A(B[9]), .B(B[10]), .CI(n719), .CO(n718), .S(n1388) );
  FA_X1 U1126 ( .A(B[8]), .B(B[9]), .CI(n720), .CO(n719), .S(n1389) );
  FA_X1 U1127 ( .A(B[7]), .B(B[8]), .CI(n721), .CO(n720), .S(n1390) );
  FA_X1 U1128 ( .A(B[6]), .B(B[7]), .CI(n722), .CO(n721), .S(n1391) );
  FA_X1 U1129 ( .A(B[5]), .B(B[6]), .CI(n723), .CO(n722), .S(n1392) );
  FA_X1 U1130 ( .A(B[4]), .B(B[5]), .CI(n724), .CO(n723), .S(n1393) );
  FA_X1 U1131 ( .A(B[3]), .B(B[4]), .CI(n725), .CO(n724), .S(n1394) );
  FA_X1 U1132 ( .A(B[2]), .B(B[3]), .CI(n726), .CO(n725), .S(n1395) );
  FA_X1 U1133 ( .A(B[1]), .B(B[2]), .CI(n727), .CO(n726), .S(n1396) );
  HA_X1 U1134 ( .A(B[0]), .B(B[1]), .CO(n727), .S(n1397) );
  OR2_X1 U1138 ( .A1(n2134), .A2(n2133), .ZN(n1534) );
  INV_X1 U1139 ( .A(n1534), .ZN(n1536) );
  INV_X1 U1140 ( .A(n1535), .ZN(n1537) );
  BUF_X1 U1141 ( .A(n1980), .Z(n1538) );
  BUF_X1 U1142 ( .A(n1980), .Z(n1539) );
  NAND3_X1 U1143 ( .A1(n1673), .A2(n1672), .A3(n1671), .ZN(n1586) );
  NAND3_X1 U1144 ( .A1(n1854), .A2(n1853), .A3(n1852), .ZN(n1804) );
  NAND3_X1 U1145 ( .A1(n1794), .A2(n1793), .A3(n1792), .ZN(n1744) );
  NAND3_X1 U1146 ( .A1(n1734), .A2(n1733), .A3(n1732), .ZN(n1684) );
  NAND3_X1 U1147 ( .A1(n2111), .A2(n2112), .A3(n2113), .ZN(n1563) );
  NAND2_X1 U1148 ( .A1(n1911), .A2(n1913), .ZN(n1857) );
  NAND2_X1 U1149 ( .A1(n1851), .A2(n1853), .ZN(n1797) );
  NAND2_X1 U1150 ( .A1(n1791), .A2(n1793), .ZN(n1737) );
  NAND2_X1 U1151 ( .A1(n1731), .A2(n1733), .ZN(n1677) );
  INV_X1 U1152 ( .A(n1553), .ZN(n1552) );
  INV_X1 U1153 ( .A(n1549), .ZN(n1548) );
  INV_X1 U1154 ( .A(n1551), .ZN(n1550) );
  NAND3_X1 U1155 ( .A1(n1914), .A2(n1913), .A3(n1912), .ZN(n1864) );
  NAND3_X1 U1156 ( .A1(n1974), .A2(n1973), .A3(n1972), .ZN(n1924) );
  NAND2_X1 U1157 ( .A1(n2134), .A2(n2132), .ZN(n1976) );
  NAND2_X1 U1158 ( .A1(n1971), .A2(n1973), .ZN(n1917) );
  INV_X1 U1159 ( .A(n1541), .ZN(n1540) );
  INV_X1 U1160 ( .A(n1543), .ZN(n1542) );
  INV_X1 U1161 ( .A(n1545), .ZN(n1544) );
  INV_X1 U1162 ( .A(n1547), .ZN(n1546) );
  INV_X1 U1163 ( .A(n1555), .ZN(n1554) );
  OR2_X1 U1164 ( .A1(n2132), .A2(n2131), .ZN(n1535) );
  NAND2_X1 U1165 ( .A1(A[0]), .A2(n2111), .ZN(n1561) );
  INV_X2 U1166 ( .A(B[0]), .ZN(n1574) );
  INV_X1 U1167 ( .A(A[5]), .ZN(n1553) );
  INV_X1 U1168 ( .A(A[11]), .ZN(n1549) );
  INV_X1 U1169 ( .A(A[8]), .ZN(n1551) );
  INV_X1 U1170 ( .A(A[17]), .ZN(n1545) );
  INV_X1 U1171 ( .A(A[14]), .ZN(n1547) );
  INV_X1 U1172 ( .A(A[23]), .ZN(n1541) );
  INV_X1 U1173 ( .A(A[20]), .ZN(n1543) );
  NOR2_X4 U1174 ( .A1(n1670), .A2(n1671), .ZN(n1581) );
  NOR2_X4 U1175 ( .A1(n1672), .A2(n1673), .ZN(n1582) );
  NAND2_X2 U1176 ( .A1(n1670), .A2(n1672), .ZN(n1576) );
  NOR2_X4 U1177 ( .A1(n1731), .A2(n1732), .ZN(n1680) );
  NOR2_X4 U1178 ( .A1(n1733), .A2(n1734), .ZN(n1681) );
  NOR2_X4 U1179 ( .A1(n1791), .A2(n1792), .ZN(n1740) );
  NOR2_X4 U1180 ( .A1(n1793), .A2(n1794), .ZN(n1741) );
  NOR2_X4 U1181 ( .A1(n1851), .A2(n1852), .ZN(n1800) );
  NOR2_X4 U1182 ( .A1(n1853), .A2(n1854), .ZN(n1801) );
  NOR2_X4 U1183 ( .A1(n1911), .A2(n1912), .ZN(n1860) );
  NOR2_X4 U1184 ( .A1(n1913), .A2(n1914), .ZN(n1861) );
  NOR2_X4 U1185 ( .A1(n1971), .A2(n1972), .ZN(n1920) );
  NOR2_X4 U1186 ( .A1(n1973), .A2(n1974), .ZN(n1921) );
  NOR2_X4 U1187 ( .A1(n2112), .A2(n2111), .ZN(n1558) );
  NOR2_X4 U1188 ( .A1(n2113), .A2(A[0]), .ZN(n1559) );
  INV_X1 U1189 ( .A(B[23]), .ZN(n1555) );
  INV_X1 U1190 ( .A(B[23]), .ZN(n1556) );
  XNOR2_X1 U1191 ( .A(A[2]), .B(n1557), .ZN(n908) );
  AOI221_X1 U1192 ( .B1(B[22]), .B2(n1558), .C1(B[21]), .C2(n1559), .A(n1560), 
        .ZN(n1557) );
  OAI22_X1 U1193 ( .A1(n1561), .A2(n1562), .B1(n1563), .B2(n1564), .ZN(n1560)
         );
  XNOR2_X1 U1194 ( .A(A[2]), .B(n1565), .ZN(n907) );
  AOI221_X1 U1195 ( .B1(B[23]), .B2(n1558), .C1(n1559), .C2(B[22]), .A(n1566), 
        .ZN(n1565) );
  OAI22_X1 U1196 ( .A1(n1561), .A2(n1567), .B1(n1568), .B2(n1563), .ZN(n1566)
         );
  XNOR2_X1 U1197 ( .A(A[2]), .B(n1569), .ZN(n906) );
  AOI221_X1 U1198 ( .B1(B[23]), .B2(n1558), .C1(n1554), .C2(n1559), .A(n1570), 
        .ZN(n1569) );
  OAI22_X1 U1199 ( .A1(n1561), .A2(n1571), .B1(n1572), .B2(n1563), .ZN(n1570)
         );
  XNOR2_X1 U1200 ( .A(n1573), .B(n1553), .ZN(n904) );
  OAI22_X1 U1201 ( .A1(n1574), .A2(n1575), .B1(n1576), .B2(n1574), .ZN(n1573)
         );
  XNOR2_X1 U1202 ( .A(n1577), .B(n1553), .ZN(n903) );
  OAI222_X1 U1203 ( .A1(n1575), .A2(n1578), .B1(n1574), .B2(n1579), .C1(n1576), 
        .C2(n1580), .ZN(n1577) );
  INV_X1 U1204 ( .A(n1581), .ZN(n1579) );
  INV_X1 U1205 ( .A(n1582), .ZN(n1575) );
  XNOR2_X1 U1206 ( .A(n1552), .B(n1583), .ZN(n902) );
  AOI221_X1 U1207 ( .B1(B[2]), .B2(n1582), .C1(B[1]), .C2(n1581), .A(n1584), 
        .ZN(n1583) );
  OAI22_X1 U1208 ( .A1(n1576), .A2(n1585), .B1(n1574), .B2(n1586), .ZN(n1584)
         );
  XNOR2_X1 U1209 ( .A(n1552), .B(n1587), .ZN(n901) );
  AOI221_X1 U1210 ( .B1(B[3]), .B2(n1582), .C1(B[2]), .C2(n1581), .A(n1588), 
        .ZN(n1587) );
  OAI22_X1 U1211 ( .A1(n1576), .A2(n1589), .B1(n1578), .B2(n1586), .ZN(n1588)
         );
  XNOR2_X1 U1212 ( .A(n1552), .B(n1590), .ZN(n900) );
  AOI221_X1 U1213 ( .B1(B[4]), .B2(n1582), .C1(B[3]), .C2(n1581), .A(n1591), 
        .ZN(n1590) );
  OAI22_X1 U1214 ( .A1(n1576), .A2(n1592), .B1(n1593), .B2(n1586), .ZN(n1591)
         );
  XNOR2_X1 U1215 ( .A(n1552), .B(n1594), .ZN(n899) );
  AOI221_X1 U1216 ( .B1(B[5]), .B2(n1582), .C1(B[4]), .C2(n1581), .A(n1595), 
        .ZN(n1594) );
  OAI22_X1 U1217 ( .A1(n1576), .A2(n1596), .B1(n1586), .B2(n1597), .ZN(n1595)
         );
  XNOR2_X1 U1218 ( .A(n1552), .B(n1598), .ZN(n898) );
  AOI221_X1 U1219 ( .B1(B[6]), .B2(n1582), .C1(B[5]), .C2(n1581), .A(n1599), 
        .ZN(n1598) );
  OAI22_X1 U1220 ( .A1(n1576), .A2(n1600), .B1(n1586), .B2(n1601), .ZN(n1599)
         );
  XNOR2_X1 U1221 ( .A(n1552), .B(n1602), .ZN(n897) );
  AOI221_X1 U1222 ( .B1(B[7]), .B2(n1582), .C1(B[6]), .C2(n1581), .A(n1603), 
        .ZN(n1602) );
  OAI22_X1 U1223 ( .A1(n1576), .A2(n1604), .B1(n1586), .B2(n1605), .ZN(n1603)
         );
  XNOR2_X1 U1224 ( .A(n1552), .B(n1606), .ZN(n896) );
  AOI221_X1 U1225 ( .B1(B[8]), .B2(n1582), .C1(B[7]), .C2(n1581), .A(n1607), 
        .ZN(n1606) );
  OAI22_X1 U1226 ( .A1(n1576), .A2(n1608), .B1(n1586), .B2(n1609), .ZN(n1607)
         );
  XNOR2_X1 U1227 ( .A(n1552), .B(n1610), .ZN(n895) );
  AOI221_X1 U1228 ( .B1(B[9]), .B2(n1582), .C1(B[8]), .C2(n1581), .A(n1611), 
        .ZN(n1610) );
  OAI22_X1 U1229 ( .A1(n1576), .A2(n1612), .B1(n1586), .B2(n1613), .ZN(n1611)
         );
  XNOR2_X1 U1230 ( .A(n1552), .B(n1614), .ZN(n894) );
  AOI221_X1 U1231 ( .B1(B[10]), .B2(n1582), .C1(B[9]), .C2(n1581), .A(n1615), 
        .ZN(n1614) );
  OAI22_X1 U1232 ( .A1(n1576), .A2(n1616), .B1(n1586), .B2(n1617), .ZN(n1615)
         );
  XNOR2_X1 U1233 ( .A(n1552), .B(n1618), .ZN(n893) );
  AOI221_X1 U1234 ( .B1(B[11]), .B2(n1582), .C1(B[10]), .C2(n1581), .A(n1619), 
        .ZN(n1618) );
  OAI22_X1 U1235 ( .A1(n1576), .A2(n1620), .B1(n1586), .B2(n1621), .ZN(n1619)
         );
  XNOR2_X1 U1236 ( .A(n1552), .B(n1622), .ZN(n892) );
  AOI221_X1 U1237 ( .B1(B[12]), .B2(n1582), .C1(B[11]), .C2(n1581), .A(n1623), 
        .ZN(n1622) );
  OAI22_X1 U1238 ( .A1(n1576), .A2(n1624), .B1(n1586), .B2(n1625), .ZN(n1623)
         );
  XNOR2_X1 U1239 ( .A(n1552), .B(n1626), .ZN(n891) );
  AOI221_X1 U1240 ( .B1(B[13]), .B2(n1582), .C1(B[12]), .C2(n1581), .A(n1627), 
        .ZN(n1626) );
  OAI22_X1 U1241 ( .A1(n1576), .A2(n1628), .B1(n1586), .B2(n1629), .ZN(n1627)
         );
  XNOR2_X1 U1242 ( .A(n1552), .B(n1630), .ZN(n890) );
  AOI221_X1 U1243 ( .B1(B[14]), .B2(n1582), .C1(B[13]), .C2(n1581), .A(n1631), 
        .ZN(n1630) );
  OAI22_X1 U1244 ( .A1(n1576), .A2(n1632), .B1(n1586), .B2(n1633), .ZN(n1631)
         );
  XNOR2_X1 U1245 ( .A(n1552), .B(n1634), .ZN(n889) );
  AOI221_X1 U1246 ( .B1(B[15]), .B2(n1582), .C1(B[14]), .C2(n1581), .A(n1635), 
        .ZN(n1634) );
  OAI22_X1 U1247 ( .A1(n1576), .A2(n1636), .B1(n1586), .B2(n1637), .ZN(n1635)
         );
  XNOR2_X1 U1248 ( .A(n1552), .B(n1638), .ZN(n888) );
  AOI221_X1 U1249 ( .B1(B[16]), .B2(n1582), .C1(B[15]), .C2(n1581), .A(n1639), 
        .ZN(n1638) );
  OAI22_X1 U1250 ( .A1(n1576), .A2(n1640), .B1(n1586), .B2(n1641), .ZN(n1639)
         );
  XNOR2_X1 U1251 ( .A(n1552), .B(n1642), .ZN(n887) );
  AOI221_X1 U1252 ( .B1(B[17]), .B2(n1582), .C1(B[16]), .C2(n1581), .A(n1643), 
        .ZN(n1642) );
  OAI22_X1 U1253 ( .A1(n1576), .A2(n1644), .B1(n1586), .B2(n1645), .ZN(n1643)
         );
  XNOR2_X1 U1254 ( .A(n1552), .B(n1646), .ZN(n886) );
  AOI221_X1 U1255 ( .B1(B[18]), .B2(n1582), .C1(B[17]), .C2(n1581), .A(n1647), 
        .ZN(n1646) );
  OAI22_X1 U1256 ( .A1(n1576), .A2(n1648), .B1(n1586), .B2(n1649), .ZN(n1647)
         );
  XNOR2_X1 U1257 ( .A(n1552), .B(n1650), .ZN(n885) );
  AOI221_X1 U1258 ( .B1(B[19]), .B2(n1582), .C1(B[18]), .C2(n1581), .A(n1651), 
        .ZN(n1650) );
  OAI22_X1 U1259 ( .A1(n1576), .A2(n1652), .B1(n1586), .B2(n1653), .ZN(n1651)
         );
  XNOR2_X1 U1260 ( .A(A[5]), .B(n1654), .ZN(n884) );
  AOI221_X1 U1261 ( .B1(n1582), .B2(B[20]), .C1(B[19]), .C2(n1581), .A(n1655), 
        .ZN(n1654) );
  OAI22_X1 U1262 ( .A1(n1576), .A2(n1656), .B1(n1586), .B2(n1657), .ZN(n1655)
         );
  XNOR2_X1 U1263 ( .A(A[5]), .B(n1658), .ZN(n883) );
  AOI221_X1 U1264 ( .B1(n1582), .B2(B[21]), .C1(n1581), .C2(B[20]), .A(n1659), 
        .ZN(n1658) );
  OAI22_X1 U1265 ( .A1(n1576), .A2(n1660), .B1(n1586), .B2(n1661), .ZN(n1659)
         );
  XNOR2_X1 U1266 ( .A(A[5]), .B(n1662), .ZN(n882) );
  AOI221_X1 U1267 ( .B1(n1582), .B2(B[22]), .C1(n1581), .C2(B[21]), .A(n1663), 
        .ZN(n1662) );
  OAI22_X1 U1268 ( .A1(n1562), .A2(n1576), .B1(n1564), .B2(n1586), .ZN(n1663)
         );
  XNOR2_X1 U1269 ( .A(A[5]), .B(n1664), .ZN(n881) );
  AOI221_X1 U1270 ( .B1(n1582), .B2(B[23]), .C1(n1581), .C2(B[22]), .A(n1665), 
        .ZN(n1664) );
  OAI22_X1 U1271 ( .A1(n1567), .A2(n1576), .B1(n1568), .B2(n1586), .ZN(n1665)
         );
  XNOR2_X1 U1272 ( .A(A[5]), .B(n1666), .ZN(n880) );
  AOI221_X1 U1273 ( .B1(n1582), .B2(B[23]), .C1(n1581), .C2(n1554), .A(n1667), 
        .ZN(n1666) );
  OAI22_X1 U1274 ( .A1(n1571), .A2(n1576), .B1(n1572), .B2(n1586), .ZN(n1667)
         );
  XNOR2_X1 U1275 ( .A(n1552), .B(n1668), .ZN(n879) );
  OAI221_X1 U1276 ( .B1(n1556), .B2(n1586), .C1(n1556), .C2(n1576), .A(n1669), 
        .ZN(n1668) );
  OAI21_X1 U1277 ( .B1(n1582), .B2(n1581), .A(n1554), .ZN(n1669) );
  INV_X1 U1278 ( .A(n1673), .ZN(n1670) );
  XNOR2_X1 U1279 ( .A(A[3]), .B(A[4]), .ZN(n1671) );
  XNOR2_X1 U1280 ( .A(A[4]), .B(n1553), .ZN(n1672) );
  XOR2_X1 U1281 ( .A(A[3]), .B(n1674), .Z(n1673) );
  XNOR2_X1 U1282 ( .A(n1675), .B(n1551), .ZN(n878) );
  OAI22_X1 U1283 ( .A1(n1574), .A2(n1676), .B1(n1574), .B2(n1677), .ZN(n1675)
         );
  XNOR2_X1 U1284 ( .A(n1678), .B(n1551), .ZN(n877) );
  OAI222_X1 U1285 ( .A1(n1578), .A2(n1676), .B1(n1574), .B2(n1679), .C1(n1580), 
        .C2(n1677), .ZN(n1678) );
  INV_X1 U1286 ( .A(n1680), .ZN(n1679) );
  INV_X1 U1287 ( .A(n1681), .ZN(n1676) );
  XNOR2_X1 U1288 ( .A(n1550), .B(n1682), .ZN(n876) );
  AOI221_X1 U1289 ( .B1(n1681), .B2(B[2]), .C1(n1680), .C2(B[1]), .A(n1683), 
        .ZN(n1682) );
  OAI22_X1 U1290 ( .A1(n1585), .A2(n1677), .B1(n1574), .B2(n1684), .ZN(n1683)
         );
  XNOR2_X1 U1291 ( .A(n1550), .B(n1685), .ZN(n875) );
  AOI221_X1 U1292 ( .B1(n1681), .B2(B[3]), .C1(n1680), .C2(B[2]), .A(n1686), 
        .ZN(n1685) );
  OAI22_X1 U1293 ( .A1(n1589), .A2(n1677), .B1(n1578), .B2(n1684), .ZN(n1686)
         );
  XNOR2_X1 U1294 ( .A(n1550), .B(n1687), .ZN(n874) );
  AOI221_X1 U1295 ( .B1(n1681), .B2(B[4]), .C1(n1680), .C2(B[3]), .A(n1688), 
        .ZN(n1687) );
  OAI22_X1 U1296 ( .A1(n1592), .A2(n1677), .B1(n1593), .B2(n1684), .ZN(n1688)
         );
  XNOR2_X1 U1297 ( .A(n1550), .B(n1689), .ZN(n873) );
  AOI221_X1 U1298 ( .B1(n1681), .B2(B[5]), .C1(n1680), .C2(B[4]), .A(n1690), 
        .ZN(n1689) );
  OAI22_X1 U1299 ( .A1(n1596), .A2(n1677), .B1(n1597), .B2(n1684), .ZN(n1690)
         );
  XNOR2_X1 U1300 ( .A(n1550), .B(n1691), .ZN(n872) );
  AOI221_X1 U1301 ( .B1(n1681), .B2(B[6]), .C1(n1680), .C2(B[5]), .A(n1692), 
        .ZN(n1691) );
  OAI22_X1 U1302 ( .A1(n1600), .A2(n1677), .B1(n1601), .B2(n1684), .ZN(n1692)
         );
  XNOR2_X1 U1303 ( .A(n1550), .B(n1693), .ZN(n871) );
  AOI221_X1 U1304 ( .B1(n1681), .B2(B[7]), .C1(n1680), .C2(B[6]), .A(n1694), 
        .ZN(n1693) );
  OAI22_X1 U1305 ( .A1(n1604), .A2(n1677), .B1(n1605), .B2(n1684), .ZN(n1694)
         );
  XNOR2_X1 U1306 ( .A(n1550), .B(n1695), .ZN(n870) );
  AOI221_X1 U1307 ( .B1(n1681), .B2(B[8]), .C1(n1680), .C2(B[7]), .A(n1696), 
        .ZN(n1695) );
  OAI22_X1 U1308 ( .A1(n1608), .A2(n1677), .B1(n1609), .B2(n1684), .ZN(n1696)
         );
  XNOR2_X1 U1309 ( .A(n1550), .B(n1697), .ZN(n869) );
  AOI221_X1 U1310 ( .B1(n1681), .B2(B[9]), .C1(n1680), .C2(B[8]), .A(n1698), 
        .ZN(n1697) );
  OAI22_X1 U1311 ( .A1(n1612), .A2(n1677), .B1(n1613), .B2(n1684), .ZN(n1698)
         );
  XNOR2_X1 U1312 ( .A(n1550), .B(n1699), .ZN(n868) );
  AOI221_X1 U1313 ( .B1(n1681), .B2(B[10]), .C1(n1680), .C2(B[9]), .A(n1700), 
        .ZN(n1699) );
  OAI22_X1 U1314 ( .A1(n1616), .A2(n1677), .B1(n1617), .B2(n1684), .ZN(n1700)
         );
  XNOR2_X1 U1315 ( .A(n1550), .B(n1701), .ZN(n867) );
  AOI221_X1 U1316 ( .B1(n1681), .B2(B[11]), .C1(n1680), .C2(B[10]), .A(n1702), 
        .ZN(n1701) );
  OAI22_X1 U1317 ( .A1(n1620), .A2(n1677), .B1(n1621), .B2(n1684), .ZN(n1702)
         );
  XNOR2_X1 U1318 ( .A(n1550), .B(n1703), .ZN(n866) );
  AOI221_X1 U1319 ( .B1(n1681), .B2(B[12]), .C1(n1680), .C2(B[11]), .A(n1704), 
        .ZN(n1703) );
  OAI22_X1 U1320 ( .A1(n1624), .A2(n1677), .B1(n1625), .B2(n1684), .ZN(n1704)
         );
  XNOR2_X1 U1321 ( .A(n1550), .B(n1705), .ZN(n865) );
  AOI221_X1 U1322 ( .B1(n1681), .B2(B[13]), .C1(n1680), .C2(B[12]), .A(n1706), 
        .ZN(n1705) );
  OAI22_X1 U1323 ( .A1(n1628), .A2(n1677), .B1(n1629), .B2(n1684), .ZN(n1706)
         );
  XNOR2_X1 U1324 ( .A(n1550), .B(n1707), .ZN(n864) );
  AOI221_X1 U1325 ( .B1(n1681), .B2(B[14]), .C1(n1680), .C2(B[13]), .A(n1708), 
        .ZN(n1707) );
  OAI22_X1 U1326 ( .A1(n1632), .A2(n1677), .B1(n1633), .B2(n1684), .ZN(n1708)
         );
  XNOR2_X1 U1327 ( .A(n1550), .B(n1709), .ZN(n863) );
  AOI221_X1 U1328 ( .B1(n1681), .B2(B[15]), .C1(n1680), .C2(B[14]), .A(n1710), 
        .ZN(n1709) );
  OAI22_X1 U1329 ( .A1(n1636), .A2(n1677), .B1(n1637), .B2(n1684), .ZN(n1710)
         );
  XNOR2_X1 U1330 ( .A(n1550), .B(n1711), .ZN(n862) );
  AOI221_X1 U1331 ( .B1(n1681), .B2(B[16]), .C1(n1680), .C2(B[15]), .A(n1712), 
        .ZN(n1711) );
  OAI22_X1 U1332 ( .A1(n1640), .A2(n1677), .B1(n1641), .B2(n1684), .ZN(n1712)
         );
  XNOR2_X1 U1333 ( .A(n1550), .B(n1713), .ZN(n861) );
  AOI221_X1 U1334 ( .B1(n1681), .B2(B[17]), .C1(n1680), .C2(B[16]), .A(n1714), 
        .ZN(n1713) );
  OAI22_X1 U1335 ( .A1(n1644), .A2(n1677), .B1(n1645), .B2(n1684), .ZN(n1714)
         );
  XNOR2_X1 U1336 ( .A(n1550), .B(n1715), .ZN(n860) );
  AOI221_X1 U1337 ( .B1(n1681), .B2(B[18]), .C1(n1680), .C2(B[17]), .A(n1716), 
        .ZN(n1715) );
  OAI22_X1 U1338 ( .A1(n1648), .A2(n1677), .B1(n1649), .B2(n1684), .ZN(n1716)
         );
  XNOR2_X1 U1339 ( .A(n1550), .B(n1717), .ZN(n859) );
  AOI221_X1 U1340 ( .B1(n1681), .B2(B[19]), .C1(n1680), .C2(B[18]), .A(n1718), 
        .ZN(n1717) );
  OAI22_X1 U1341 ( .A1(n1652), .A2(n1677), .B1(n1653), .B2(n1684), .ZN(n1718)
         );
  XNOR2_X1 U1342 ( .A(A[8]), .B(n1719), .ZN(n858) );
  AOI221_X1 U1343 ( .B1(n1681), .B2(B[20]), .C1(n1680), .C2(B[19]), .A(n1720), 
        .ZN(n1719) );
  OAI22_X1 U1344 ( .A1(n1656), .A2(n1677), .B1(n1657), .B2(n1684), .ZN(n1720)
         );
  XNOR2_X1 U1345 ( .A(A[8]), .B(n1721), .ZN(n857) );
  AOI221_X1 U1346 ( .B1(n1681), .B2(B[21]), .C1(n1680), .C2(B[20]), .A(n1722), 
        .ZN(n1721) );
  OAI22_X1 U1347 ( .A1(n1660), .A2(n1677), .B1(n1661), .B2(n1684), .ZN(n1722)
         );
  XNOR2_X1 U1348 ( .A(A[8]), .B(n1723), .ZN(n856) );
  AOI221_X1 U1349 ( .B1(n1681), .B2(B[22]), .C1(n1680), .C2(B[21]), .A(n1724), 
        .ZN(n1723) );
  OAI22_X1 U1350 ( .A1(n1562), .A2(n1677), .B1(n1564), .B2(n1684), .ZN(n1724)
         );
  XNOR2_X1 U1351 ( .A(A[8]), .B(n1725), .ZN(n855) );
  AOI221_X1 U1352 ( .B1(n1681), .B2(B[23]), .C1(n1680), .C2(B[22]), .A(n1726), 
        .ZN(n1725) );
  OAI22_X1 U1353 ( .A1(n1567), .A2(n1677), .B1(n1568), .B2(n1684), .ZN(n1726)
         );
  XNOR2_X1 U1354 ( .A(A[8]), .B(n1727), .ZN(n854) );
  AOI221_X1 U1355 ( .B1(n1681), .B2(B[23]), .C1(n1680), .C2(n1554), .A(n1728), 
        .ZN(n1727) );
  OAI22_X1 U1356 ( .A1(n1571), .A2(n1677), .B1(n1572), .B2(n1684), .ZN(n1728)
         );
  XNOR2_X1 U1357 ( .A(n1550), .B(n1729), .ZN(n853) );
  OAI221_X1 U1358 ( .B1(n1555), .B2(n1684), .C1(n1556), .C2(n1677), .A(n1730), 
        .ZN(n1729) );
  OAI21_X1 U1359 ( .B1(n1681), .B2(n1680), .A(n1554), .ZN(n1730) );
  INV_X1 U1360 ( .A(n1734), .ZN(n1731) );
  XNOR2_X1 U1361 ( .A(A[6]), .B(A[7]), .ZN(n1732) );
  XNOR2_X1 U1362 ( .A(A[7]), .B(n1551), .ZN(n1733) );
  XOR2_X1 U1363 ( .A(A[6]), .B(n1553), .Z(n1734) );
  XNOR2_X1 U1364 ( .A(n1735), .B(n1549), .ZN(n852) );
  OAI22_X1 U1365 ( .A1(n1574), .A2(n1736), .B1(n1574), .B2(n1737), .ZN(n1735)
         );
  XNOR2_X1 U1366 ( .A(n1738), .B(n1549), .ZN(n851) );
  OAI222_X1 U1367 ( .A1(n1578), .A2(n1736), .B1(n1574), .B2(n1739), .C1(n1580), 
        .C2(n1737), .ZN(n1738) );
  INV_X1 U1368 ( .A(n1740), .ZN(n1739) );
  INV_X1 U1369 ( .A(n1741), .ZN(n1736) );
  XNOR2_X1 U1370 ( .A(n1548), .B(n1742), .ZN(n850) );
  AOI221_X1 U1371 ( .B1(n1741), .B2(B[2]), .C1(n1740), .C2(B[1]), .A(n1743), 
        .ZN(n1742) );
  OAI22_X1 U1372 ( .A1(n1585), .A2(n1737), .B1(n1574), .B2(n1744), .ZN(n1743)
         );
  XNOR2_X1 U1373 ( .A(n1548), .B(n1745), .ZN(n849) );
  AOI221_X1 U1374 ( .B1(n1741), .B2(B[3]), .C1(n1740), .C2(B[2]), .A(n1746), 
        .ZN(n1745) );
  OAI22_X1 U1375 ( .A1(n1589), .A2(n1737), .B1(n1578), .B2(n1744), .ZN(n1746)
         );
  XNOR2_X1 U1376 ( .A(n1548), .B(n1747), .ZN(n848) );
  AOI221_X1 U1377 ( .B1(n1741), .B2(B[4]), .C1(n1740), .C2(B[3]), .A(n1748), 
        .ZN(n1747) );
  OAI22_X1 U1378 ( .A1(n1592), .A2(n1737), .B1(n1593), .B2(n1744), .ZN(n1748)
         );
  XNOR2_X1 U1379 ( .A(n1548), .B(n1749), .ZN(n847) );
  AOI221_X1 U1380 ( .B1(n1741), .B2(B[5]), .C1(n1740), .C2(B[4]), .A(n1750), 
        .ZN(n1749) );
  OAI22_X1 U1381 ( .A1(n1596), .A2(n1737), .B1(n1597), .B2(n1744), .ZN(n1750)
         );
  XNOR2_X1 U1382 ( .A(n1548), .B(n1751), .ZN(n846) );
  AOI221_X1 U1383 ( .B1(n1741), .B2(B[6]), .C1(n1740), .C2(B[5]), .A(n1752), 
        .ZN(n1751) );
  OAI22_X1 U1384 ( .A1(n1600), .A2(n1737), .B1(n1601), .B2(n1744), .ZN(n1752)
         );
  XNOR2_X1 U1385 ( .A(n1548), .B(n1753), .ZN(n845) );
  AOI221_X1 U1386 ( .B1(n1741), .B2(B[7]), .C1(n1740), .C2(B[6]), .A(n1754), 
        .ZN(n1753) );
  OAI22_X1 U1387 ( .A1(n1604), .A2(n1737), .B1(n1605), .B2(n1744), .ZN(n1754)
         );
  XNOR2_X1 U1388 ( .A(n1548), .B(n1755), .ZN(n844) );
  AOI221_X1 U1389 ( .B1(n1741), .B2(B[8]), .C1(n1740), .C2(B[7]), .A(n1756), 
        .ZN(n1755) );
  OAI22_X1 U1390 ( .A1(n1608), .A2(n1737), .B1(n1609), .B2(n1744), .ZN(n1756)
         );
  XNOR2_X1 U1391 ( .A(n1548), .B(n1757), .ZN(n843) );
  AOI221_X1 U1392 ( .B1(n1741), .B2(B[9]), .C1(n1740), .C2(B[8]), .A(n1758), 
        .ZN(n1757) );
  OAI22_X1 U1393 ( .A1(n1612), .A2(n1737), .B1(n1613), .B2(n1744), .ZN(n1758)
         );
  XNOR2_X1 U1394 ( .A(n1548), .B(n1759), .ZN(n842) );
  AOI221_X1 U1395 ( .B1(n1741), .B2(B[10]), .C1(n1740), .C2(B[9]), .A(n1760), 
        .ZN(n1759) );
  OAI22_X1 U1396 ( .A1(n1616), .A2(n1737), .B1(n1617), .B2(n1744), .ZN(n1760)
         );
  XNOR2_X1 U1397 ( .A(n1548), .B(n1761), .ZN(n841) );
  AOI221_X1 U1398 ( .B1(n1741), .B2(B[11]), .C1(n1740), .C2(B[10]), .A(n1762), 
        .ZN(n1761) );
  OAI22_X1 U1399 ( .A1(n1620), .A2(n1737), .B1(n1621), .B2(n1744), .ZN(n1762)
         );
  XNOR2_X1 U1400 ( .A(n1548), .B(n1763), .ZN(n840) );
  AOI221_X1 U1401 ( .B1(n1741), .B2(B[12]), .C1(n1740), .C2(B[11]), .A(n1764), 
        .ZN(n1763) );
  OAI22_X1 U1402 ( .A1(n1624), .A2(n1737), .B1(n1625), .B2(n1744), .ZN(n1764)
         );
  XNOR2_X1 U1403 ( .A(n1548), .B(n1765), .ZN(n839) );
  AOI221_X1 U1404 ( .B1(n1741), .B2(B[13]), .C1(n1740), .C2(B[12]), .A(n1766), 
        .ZN(n1765) );
  OAI22_X1 U1405 ( .A1(n1628), .A2(n1737), .B1(n1629), .B2(n1744), .ZN(n1766)
         );
  XNOR2_X1 U1406 ( .A(n1548), .B(n1767), .ZN(n838) );
  AOI221_X1 U1407 ( .B1(n1741), .B2(B[14]), .C1(n1740), .C2(B[13]), .A(n1768), 
        .ZN(n1767) );
  OAI22_X1 U1408 ( .A1(n1632), .A2(n1737), .B1(n1633), .B2(n1744), .ZN(n1768)
         );
  XNOR2_X1 U1409 ( .A(n1548), .B(n1769), .ZN(n837) );
  AOI221_X1 U1410 ( .B1(n1741), .B2(B[15]), .C1(n1740), .C2(B[14]), .A(n1770), 
        .ZN(n1769) );
  OAI22_X1 U1411 ( .A1(n1636), .A2(n1737), .B1(n1637), .B2(n1744), .ZN(n1770)
         );
  XNOR2_X1 U1412 ( .A(n1548), .B(n1771), .ZN(n836) );
  AOI221_X1 U1413 ( .B1(n1741), .B2(B[16]), .C1(n1740), .C2(B[15]), .A(n1772), 
        .ZN(n1771) );
  OAI22_X1 U1414 ( .A1(n1640), .A2(n1737), .B1(n1641), .B2(n1744), .ZN(n1772)
         );
  XNOR2_X1 U1415 ( .A(n1548), .B(n1773), .ZN(n835) );
  AOI221_X1 U1416 ( .B1(n1741), .B2(B[17]), .C1(n1740), .C2(B[16]), .A(n1774), 
        .ZN(n1773) );
  OAI22_X1 U1417 ( .A1(n1644), .A2(n1737), .B1(n1645), .B2(n1744), .ZN(n1774)
         );
  XNOR2_X1 U1418 ( .A(n1548), .B(n1775), .ZN(n834) );
  AOI221_X1 U1419 ( .B1(n1741), .B2(B[18]), .C1(n1740), .C2(B[17]), .A(n1776), 
        .ZN(n1775) );
  OAI22_X1 U1420 ( .A1(n1648), .A2(n1737), .B1(n1649), .B2(n1744), .ZN(n1776)
         );
  XNOR2_X1 U1421 ( .A(n1548), .B(n1777), .ZN(n833) );
  AOI221_X1 U1422 ( .B1(n1741), .B2(B[19]), .C1(n1740), .C2(B[18]), .A(n1778), 
        .ZN(n1777) );
  OAI22_X1 U1423 ( .A1(n1652), .A2(n1737), .B1(n1653), .B2(n1744), .ZN(n1778)
         );
  XNOR2_X1 U1424 ( .A(n1548), .B(n1779), .ZN(n832) );
  AOI221_X1 U1425 ( .B1(n1741), .B2(B[20]), .C1(n1740), .C2(B[19]), .A(n1780), 
        .ZN(n1779) );
  OAI22_X1 U1426 ( .A1(n1656), .A2(n1737), .B1(n1657), .B2(n1744), .ZN(n1780)
         );
  XNOR2_X1 U1427 ( .A(A[11]), .B(n1781), .ZN(n831) );
  AOI221_X1 U1428 ( .B1(n1741), .B2(B[21]), .C1(n1740), .C2(B[20]), .A(n1782), 
        .ZN(n1781) );
  OAI22_X1 U1429 ( .A1(n1660), .A2(n1737), .B1(n1661), .B2(n1744), .ZN(n1782)
         );
  XNOR2_X1 U1430 ( .A(A[11]), .B(n1783), .ZN(n830) );
  AOI221_X1 U1431 ( .B1(n1741), .B2(B[22]), .C1(n1740), .C2(B[21]), .A(n1784), 
        .ZN(n1783) );
  OAI22_X1 U1432 ( .A1(n1562), .A2(n1737), .B1(n1564), .B2(n1744), .ZN(n1784)
         );
  XNOR2_X1 U1433 ( .A(A[11]), .B(n1785), .ZN(n829) );
  AOI221_X1 U1434 ( .B1(n1741), .B2(B[23]), .C1(n1740), .C2(B[22]), .A(n1786), 
        .ZN(n1785) );
  OAI22_X1 U1435 ( .A1(n1567), .A2(n1737), .B1(n1568), .B2(n1744), .ZN(n1786)
         );
  XNOR2_X1 U1436 ( .A(A[11]), .B(n1787), .ZN(n828) );
  AOI221_X1 U1437 ( .B1(n1741), .B2(B[23]), .C1(n1740), .C2(n1554), .A(n1788), 
        .ZN(n1787) );
  OAI22_X1 U1438 ( .A1(n1571), .A2(n1737), .B1(n1572), .B2(n1744), .ZN(n1788)
         );
  XNOR2_X1 U1439 ( .A(A[11]), .B(n1789), .ZN(n827) );
  OAI221_X1 U1440 ( .B1(n1556), .B2(n1744), .C1(n1556), .C2(n1737), .A(n1790), 
        .ZN(n1789) );
  OAI21_X1 U1441 ( .B1(n1741), .B2(n1740), .A(n1554), .ZN(n1790) );
  INV_X1 U1442 ( .A(n1794), .ZN(n1791) );
  XNOR2_X1 U1443 ( .A(A[10]), .B(A[9]), .ZN(n1792) );
  XNOR2_X1 U1444 ( .A(A[10]), .B(n1549), .ZN(n1793) );
  XOR2_X1 U1445 ( .A(A[9]), .B(n1551), .Z(n1794) );
  XNOR2_X1 U1446 ( .A(n1795), .B(n1547), .ZN(n826) );
  OAI22_X1 U1447 ( .A1(n1574), .A2(n1796), .B1(n1574), .B2(n1797), .ZN(n1795)
         );
  XNOR2_X1 U1448 ( .A(n1798), .B(n1547), .ZN(n825) );
  OAI222_X1 U1449 ( .A1(n1578), .A2(n1796), .B1(n1574), .B2(n1799), .C1(n1580), 
        .C2(n1797), .ZN(n1798) );
  INV_X1 U1450 ( .A(n1800), .ZN(n1799) );
  INV_X1 U1451 ( .A(n1801), .ZN(n1796) );
  XNOR2_X1 U1452 ( .A(n1546), .B(n1802), .ZN(n824) );
  AOI221_X1 U1453 ( .B1(n1801), .B2(B[2]), .C1(n1800), .C2(B[1]), .A(n1803), 
        .ZN(n1802) );
  OAI22_X1 U1454 ( .A1(n1585), .A2(n1797), .B1(n1574), .B2(n1804), .ZN(n1803)
         );
  XNOR2_X1 U1455 ( .A(n1546), .B(n1805), .ZN(n823) );
  AOI221_X1 U1456 ( .B1(n1801), .B2(B[3]), .C1(n1800), .C2(B[2]), .A(n1806), 
        .ZN(n1805) );
  OAI22_X1 U1457 ( .A1(n1589), .A2(n1797), .B1(n1578), .B2(n1804), .ZN(n1806)
         );
  XNOR2_X1 U1458 ( .A(n1546), .B(n1807), .ZN(n822) );
  AOI221_X1 U1459 ( .B1(n1801), .B2(B[4]), .C1(n1800), .C2(B[3]), .A(n1808), 
        .ZN(n1807) );
  OAI22_X1 U1460 ( .A1(n1592), .A2(n1797), .B1(n1593), .B2(n1804), .ZN(n1808)
         );
  XNOR2_X1 U1461 ( .A(n1546), .B(n1809), .ZN(n821) );
  AOI221_X1 U1462 ( .B1(n1801), .B2(B[5]), .C1(n1800), .C2(B[4]), .A(n1810), 
        .ZN(n1809) );
  OAI22_X1 U1463 ( .A1(n1596), .A2(n1797), .B1(n1597), .B2(n1804), .ZN(n1810)
         );
  XNOR2_X1 U1464 ( .A(n1546), .B(n1811), .ZN(n820) );
  AOI221_X1 U1465 ( .B1(n1801), .B2(B[6]), .C1(n1800), .C2(B[5]), .A(n1812), 
        .ZN(n1811) );
  OAI22_X1 U1466 ( .A1(n1600), .A2(n1797), .B1(n1601), .B2(n1804), .ZN(n1812)
         );
  XNOR2_X1 U1467 ( .A(n1546), .B(n1813), .ZN(n819) );
  AOI221_X1 U1468 ( .B1(n1801), .B2(B[7]), .C1(n1800), .C2(B[6]), .A(n1814), 
        .ZN(n1813) );
  OAI22_X1 U1469 ( .A1(n1604), .A2(n1797), .B1(n1605), .B2(n1804), .ZN(n1814)
         );
  XNOR2_X1 U1470 ( .A(n1546), .B(n1815), .ZN(n818) );
  AOI221_X1 U1471 ( .B1(n1801), .B2(B[8]), .C1(n1800), .C2(B[7]), .A(n1816), 
        .ZN(n1815) );
  OAI22_X1 U1472 ( .A1(n1608), .A2(n1797), .B1(n1609), .B2(n1804), .ZN(n1816)
         );
  XNOR2_X1 U1473 ( .A(n1546), .B(n1817), .ZN(n817) );
  AOI221_X1 U1474 ( .B1(n1801), .B2(B[9]), .C1(n1800), .C2(B[8]), .A(n1818), 
        .ZN(n1817) );
  OAI22_X1 U1475 ( .A1(n1612), .A2(n1797), .B1(n1613), .B2(n1804), .ZN(n1818)
         );
  XNOR2_X1 U1476 ( .A(n1546), .B(n1819), .ZN(n816) );
  AOI221_X1 U1477 ( .B1(n1801), .B2(B[10]), .C1(n1800), .C2(B[9]), .A(n1820), 
        .ZN(n1819) );
  OAI22_X1 U1478 ( .A1(n1616), .A2(n1797), .B1(n1617), .B2(n1804), .ZN(n1820)
         );
  XNOR2_X1 U1479 ( .A(n1546), .B(n1821), .ZN(n815) );
  AOI221_X1 U1480 ( .B1(n1801), .B2(B[11]), .C1(n1800), .C2(B[10]), .A(n1822), 
        .ZN(n1821) );
  OAI22_X1 U1481 ( .A1(n1620), .A2(n1797), .B1(n1621), .B2(n1804), .ZN(n1822)
         );
  XNOR2_X1 U1482 ( .A(n1546), .B(n1823), .ZN(n814) );
  AOI221_X1 U1483 ( .B1(n1801), .B2(B[12]), .C1(n1800), .C2(B[11]), .A(n1824), 
        .ZN(n1823) );
  OAI22_X1 U1484 ( .A1(n1624), .A2(n1797), .B1(n1625), .B2(n1804), .ZN(n1824)
         );
  XNOR2_X1 U1485 ( .A(n1546), .B(n1825), .ZN(n813) );
  AOI221_X1 U1486 ( .B1(n1801), .B2(B[13]), .C1(n1800), .C2(B[12]), .A(n1826), 
        .ZN(n1825) );
  OAI22_X1 U1487 ( .A1(n1628), .A2(n1797), .B1(n1629), .B2(n1804), .ZN(n1826)
         );
  XNOR2_X1 U1488 ( .A(n1546), .B(n1827), .ZN(n812) );
  AOI221_X1 U1489 ( .B1(n1801), .B2(B[14]), .C1(n1800), .C2(B[13]), .A(n1828), 
        .ZN(n1827) );
  OAI22_X1 U1490 ( .A1(n1632), .A2(n1797), .B1(n1633), .B2(n1804), .ZN(n1828)
         );
  XNOR2_X1 U1491 ( .A(n1546), .B(n1829), .ZN(n811) );
  AOI221_X1 U1492 ( .B1(n1801), .B2(B[15]), .C1(n1800), .C2(B[14]), .A(n1830), 
        .ZN(n1829) );
  OAI22_X1 U1493 ( .A1(n1636), .A2(n1797), .B1(n1637), .B2(n1804), .ZN(n1830)
         );
  XNOR2_X1 U1494 ( .A(n1546), .B(n1831), .ZN(n810) );
  AOI221_X1 U1495 ( .B1(n1801), .B2(B[16]), .C1(n1800), .C2(B[15]), .A(n1832), 
        .ZN(n1831) );
  OAI22_X1 U1496 ( .A1(n1640), .A2(n1797), .B1(n1641), .B2(n1804), .ZN(n1832)
         );
  XNOR2_X1 U1497 ( .A(n1546), .B(n1833), .ZN(n809) );
  AOI221_X1 U1498 ( .B1(n1801), .B2(B[17]), .C1(n1800), .C2(B[16]), .A(n1834), 
        .ZN(n1833) );
  OAI22_X1 U1499 ( .A1(n1644), .A2(n1797), .B1(n1645), .B2(n1804), .ZN(n1834)
         );
  XNOR2_X1 U1500 ( .A(n1546), .B(n1835), .ZN(n808) );
  AOI221_X1 U1501 ( .B1(n1801), .B2(B[18]), .C1(n1800), .C2(B[17]), .A(n1836), 
        .ZN(n1835) );
  OAI22_X1 U1502 ( .A1(n1648), .A2(n1797), .B1(n1649), .B2(n1804), .ZN(n1836)
         );
  XNOR2_X1 U1503 ( .A(n1546), .B(n1837), .ZN(n807) );
  AOI221_X1 U1504 ( .B1(n1801), .B2(B[19]), .C1(n1800), .C2(B[18]), .A(n1838), 
        .ZN(n1837) );
  OAI22_X1 U1505 ( .A1(n1652), .A2(n1797), .B1(n1653), .B2(n1804), .ZN(n1838)
         );
  XNOR2_X1 U1506 ( .A(n1546), .B(n1839), .ZN(n806) );
  AOI221_X1 U1507 ( .B1(n1801), .B2(B[20]), .C1(n1800), .C2(B[19]), .A(n1840), 
        .ZN(n1839) );
  OAI22_X1 U1508 ( .A1(n1656), .A2(n1797), .B1(n1657), .B2(n1804), .ZN(n1840)
         );
  XNOR2_X1 U1509 ( .A(A[14]), .B(n1841), .ZN(n805) );
  AOI221_X1 U1510 ( .B1(n1801), .B2(B[21]), .C1(n1800), .C2(B[20]), .A(n1842), 
        .ZN(n1841) );
  OAI22_X1 U1511 ( .A1(n1660), .A2(n1797), .B1(n1661), .B2(n1804), .ZN(n1842)
         );
  XNOR2_X1 U1512 ( .A(A[14]), .B(n1843), .ZN(n804) );
  AOI221_X1 U1513 ( .B1(n1801), .B2(B[22]), .C1(n1800), .C2(B[21]), .A(n1844), 
        .ZN(n1843) );
  OAI22_X1 U1514 ( .A1(n1562), .A2(n1797), .B1(n1564), .B2(n1804), .ZN(n1844)
         );
  XNOR2_X1 U1515 ( .A(A[14]), .B(n1845), .ZN(n803) );
  AOI221_X1 U1516 ( .B1(n1801), .B2(B[23]), .C1(n1800), .C2(B[22]), .A(n1846), 
        .ZN(n1845) );
  OAI22_X1 U1517 ( .A1(n1567), .A2(n1797), .B1(n1568), .B2(n1804), .ZN(n1846)
         );
  XNOR2_X1 U1518 ( .A(A[14]), .B(n1847), .ZN(n802) );
  AOI221_X1 U1519 ( .B1(n1801), .B2(B[23]), .C1(n1800), .C2(n1554), .A(n1848), 
        .ZN(n1847) );
  OAI22_X1 U1520 ( .A1(n1571), .A2(n1797), .B1(n1572), .B2(n1804), .ZN(n1848)
         );
  XNOR2_X1 U1521 ( .A(A[14]), .B(n1849), .ZN(n801) );
  OAI221_X1 U1522 ( .B1(n1556), .B2(n1804), .C1(n1556), .C2(n1797), .A(n1850), 
        .ZN(n1849) );
  OAI21_X1 U1523 ( .B1(n1801), .B2(n1800), .A(n1554), .ZN(n1850) );
  INV_X1 U1524 ( .A(n1854), .ZN(n1851) );
  XNOR2_X1 U1525 ( .A(A[12]), .B(A[13]), .ZN(n1852) );
  XNOR2_X1 U1526 ( .A(A[13]), .B(n1547), .ZN(n1853) );
  XOR2_X1 U1527 ( .A(A[12]), .B(n1549), .Z(n1854) );
  XNOR2_X1 U1528 ( .A(n1855), .B(n1545), .ZN(n800) );
  OAI22_X1 U1529 ( .A1(n1574), .A2(n1856), .B1(n1574), .B2(n1857), .ZN(n1855)
         );
  XNOR2_X1 U1530 ( .A(n1858), .B(n1545), .ZN(n799) );
  OAI222_X1 U1531 ( .A1(n1578), .A2(n1856), .B1(n1574), .B2(n1859), .C1(n1580), 
        .C2(n1857), .ZN(n1858) );
  INV_X1 U1532 ( .A(n1860), .ZN(n1859) );
  INV_X1 U1533 ( .A(n1861), .ZN(n1856) );
  XNOR2_X1 U1534 ( .A(n1544), .B(n1862), .ZN(n798) );
  AOI221_X1 U1535 ( .B1(n1861), .B2(B[2]), .C1(n1860), .C2(B[1]), .A(n1863), 
        .ZN(n1862) );
  OAI22_X1 U1536 ( .A1(n1585), .A2(n1857), .B1(n1574), .B2(n1864), .ZN(n1863)
         );
  XNOR2_X1 U1537 ( .A(n1544), .B(n1865), .ZN(n797) );
  AOI221_X1 U1538 ( .B1(n1861), .B2(B[3]), .C1(n1860), .C2(B[2]), .A(n1866), 
        .ZN(n1865) );
  OAI22_X1 U1539 ( .A1(n1589), .A2(n1857), .B1(n1578), .B2(n1864), .ZN(n1866)
         );
  XNOR2_X1 U1540 ( .A(n1544), .B(n1867), .ZN(n796) );
  AOI221_X1 U1541 ( .B1(n1861), .B2(B[4]), .C1(n1860), .C2(B[3]), .A(n1868), 
        .ZN(n1867) );
  OAI22_X1 U1542 ( .A1(n1592), .A2(n1857), .B1(n1593), .B2(n1864), .ZN(n1868)
         );
  XNOR2_X1 U1543 ( .A(n1544), .B(n1869), .ZN(n795) );
  AOI221_X1 U1544 ( .B1(n1861), .B2(B[5]), .C1(n1860), .C2(B[4]), .A(n1870), 
        .ZN(n1869) );
  OAI22_X1 U1545 ( .A1(n1596), .A2(n1857), .B1(n1597), .B2(n1864), .ZN(n1870)
         );
  XNOR2_X1 U1546 ( .A(n1544), .B(n1871), .ZN(n794) );
  AOI221_X1 U1547 ( .B1(n1861), .B2(B[6]), .C1(n1860), .C2(B[5]), .A(n1872), 
        .ZN(n1871) );
  OAI22_X1 U1548 ( .A1(n1600), .A2(n1857), .B1(n1601), .B2(n1864), .ZN(n1872)
         );
  XNOR2_X1 U1549 ( .A(n1544), .B(n1873), .ZN(n793) );
  AOI221_X1 U1550 ( .B1(n1861), .B2(B[7]), .C1(n1860), .C2(B[6]), .A(n1874), 
        .ZN(n1873) );
  OAI22_X1 U1551 ( .A1(n1604), .A2(n1857), .B1(n1605), .B2(n1864), .ZN(n1874)
         );
  XNOR2_X1 U1552 ( .A(n1544), .B(n1875), .ZN(n792) );
  AOI221_X1 U1553 ( .B1(n1861), .B2(B[8]), .C1(n1860), .C2(B[7]), .A(n1876), 
        .ZN(n1875) );
  OAI22_X1 U1554 ( .A1(n1608), .A2(n1857), .B1(n1609), .B2(n1864), .ZN(n1876)
         );
  XNOR2_X1 U1555 ( .A(n1544), .B(n1877), .ZN(n791) );
  AOI221_X1 U1556 ( .B1(n1861), .B2(B[9]), .C1(n1860), .C2(B[8]), .A(n1878), 
        .ZN(n1877) );
  OAI22_X1 U1557 ( .A1(n1612), .A2(n1857), .B1(n1613), .B2(n1864), .ZN(n1878)
         );
  XNOR2_X1 U1558 ( .A(n1544), .B(n1879), .ZN(n790) );
  AOI221_X1 U1559 ( .B1(n1861), .B2(B[10]), .C1(n1860), .C2(B[9]), .A(n1880), 
        .ZN(n1879) );
  OAI22_X1 U1560 ( .A1(n1616), .A2(n1857), .B1(n1617), .B2(n1864), .ZN(n1880)
         );
  XNOR2_X1 U1561 ( .A(n1544), .B(n1881), .ZN(n789) );
  AOI221_X1 U1562 ( .B1(n1861), .B2(B[11]), .C1(n1860), .C2(B[10]), .A(n1882), 
        .ZN(n1881) );
  OAI22_X1 U1563 ( .A1(n1620), .A2(n1857), .B1(n1621), .B2(n1864), .ZN(n1882)
         );
  XNOR2_X1 U1564 ( .A(n1544), .B(n1883), .ZN(n788) );
  AOI221_X1 U1565 ( .B1(n1861), .B2(B[12]), .C1(n1860), .C2(B[11]), .A(n1884), 
        .ZN(n1883) );
  OAI22_X1 U1566 ( .A1(n1624), .A2(n1857), .B1(n1625), .B2(n1864), .ZN(n1884)
         );
  XNOR2_X1 U1567 ( .A(n1544), .B(n1885), .ZN(n787) );
  AOI221_X1 U1568 ( .B1(n1861), .B2(B[13]), .C1(n1860), .C2(B[12]), .A(n1886), 
        .ZN(n1885) );
  OAI22_X1 U1569 ( .A1(n1628), .A2(n1857), .B1(n1629), .B2(n1864), .ZN(n1886)
         );
  XNOR2_X1 U1570 ( .A(n1544), .B(n1887), .ZN(n786) );
  AOI221_X1 U1571 ( .B1(n1861), .B2(B[14]), .C1(n1860), .C2(B[13]), .A(n1888), 
        .ZN(n1887) );
  OAI22_X1 U1572 ( .A1(n1632), .A2(n1857), .B1(n1633), .B2(n1864), .ZN(n1888)
         );
  XNOR2_X1 U1573 ( .A(n1544), .B(n1889), .ZN(n785) );
  AOI221_X1 U1574 ( .B1(n1861), .B2(B[15]), .C1(n1860), .C2(B[14]), .A(n1890), 
        .ZN(n1889) );
  OAI22_X1 U1575 ( .A1(n1636), .A2(n1857), .B1(n1637), .B2(n1864), .ZN(n1890)
         );
  XNOR2_X1 U1576 ( .A(n1544), .B(n1891), .ZN(n784) );
  AOI221_X1 U1577 ( .B1(n1861), .B2(B[16]), .C1(n1860), .C2(B[15]), .A(n1892), 
        .ZN(n1891) );
  OAI22_X1 U1578 ( .A1(n1640), .A2(n1857), .B1(n1641), .B2(n1864), .ZN(n1892)
         );
  XNOR2_X1 U1579 ( .A(n1544), .B(n1893), .ZN(n783) );
  AOI221_X1 U1580 ( .B1(n1861), .B2(B[17]), .C1(n1860), .C2(B[16]), .A(n1894), 
        .ZN(n1893) );
  OAI22_X1 U1581 ( .A1(n1644), .A2(n1857), .B1(n1645), .B2(n1864), .ZN(n1894)
         );
  XNOR2_X1 U1582 ( .A(n1544), .B(n1895), .ZN(n782) );
  AOI221_X1 U1583 ( .B1(n1861), .B2(B[18]), .C1(n1860), .C2(B[17]), .A(n1896), 
        .ZN(n1895) );
  OAI22_X1 U1584 ( .A1(n1648), .A2(n1857), .B1(n1649), .B2(n1864), .ZN(n1896)
         );
  XNOR2_X1 U1585 ( .A(n1544), .B(n1897), .ZN(n781) );
  AOI221_X1 U1586 ( .B1(n1861), .B2(B[19]), .C1(n1860), .C2(B[18]), .A(n1898), 
        .ZN(n1897) );
  OAI22_X1 U1587 ( .A1(n1652), .A2(n1857), .B1(n1653), .B2(n1864), .ZN(n1898)
         );
  XNOR2_X1 U1588 ( .A(n1544), .B(n1899), .ZN(n780) );
  AOI221_X1 U1589 ( .B1(n1861), .B2(B[20]), .C1(n1860), .C2(B[19]), .A(n1900), 
        .ZN(n1899) );
  OAI22_X1 U1590 ( .A1(n1656), .A2(n1857), .B1(n1657), .B2(n1864), .ZN(n1900)
         );
  XNOR2_X1 U1591 ( .A(A[17]), .B(n1901), .ZN(n779) );
  AOI221_X1 U1592 ( .B1(n1861), .B2(B[21]), .C1(n1860), .C2(B[20]), .A(n1902), 
        .ZN(n1901) );
  OAI22_X1 U1593 ( .A1(n1660), .A2(n1857), .B1(n1661), .B2(n1864), .ZN(n1902)
         );
  XNOR2_X1 U1594 ( .A(A[17]), .B(n1903), .ZN(n778) );
  AOI221_X1 U1595 ( .B1(n1861), .B2(B[22]), .C1(n1860), .C2(B[21]), .A(n1904), 
        .ZN(n1903) );
  OAI22_X1 U1596 ( .A1(n1562), .A2(n1857), .B1(n1564), .B2(n1864), .ZN(n1904)
         );
  XNOR2_X1 U1597 ( .A(A[17]), .B(n1905), .ZN(n777) );
  AOI221_X1 U1598 ( .B1(n1861), .B2(B[23]), .C1(n1860), .C2(B[22]), .A(n1906), 
        .ZN(n1905) );
  OAI22_X1 U1599 ( .A1(n1567), .A2(n1857), .B1(n1568), .B2(n1864), .ZN(n1906)
         );
  XNOR2_X1 U1600 ( .A(A[17]), .B(n1907), .ZN(n776) );
  AOI221_X1 U1601 ( .B1(n1861), .B2(B[23]), .C1(n1860), .C2(n1554), .A(n1908), 
        .ZN(n1907) );
  OAI22_X1 U1602 ( .A1(n1571), .A2(n1857), .B1(n1572), .B2(n1864), .ZN(n1908)
         );
  XNOR2_X1 U1603 ( .A(A[17]), .B(n1909), .ZN(n775) );
  OAI221_X1 U1604 ( .B1(n1556), .B2(n1864), .C1(n1556), .C2(n1857), .A(n1910), 
        .ZN(n1909) );
  OAI21_X1 U1605 ( .B1(n1861), .B2(n1860), .A(n1554), .ZN(n1910) );
  INV_X1 U1606 ( .A(n1914), .ZN(n1911) );
  XNOR2_X1 U1607 ( .A(A[15]), .B(A[16]), .ZN(n1912) );
  XNOR2_X1 U1608 ( .A(A[16]), .B(n1545), .ZN(n1913) );
  XOR2_X1 U1609 ( .A(A[15]), .B(n1547), .Z(n1914) );
  XNOR2_X1 U1610 ( .A(n1915), .B(n1543), .ZN(n774) );
  OAI22_X1 U1611 ( .A1(n1574), .A2(n1916), .B1(n1574), .B2(n1917), .ZN(n1915)
         );
  XNOR2_X1 U1612 ( .A(n1918), .B(n1543), .ZN(n773) );
  OAI222_X1 U1613 ( .A1(n1578), .A2(n1916), .B1(n1574), .B2(n1919), .C1(n1580), 
        .C2(n1917), .ZN(n1918) );
  INV_X1 U1614 ( .A(n1920), .ZN(n1919) );
  INV_X1 U1615 ( .A(n1921), .ZN(n1916) );
  XNOR2_X1 U1616 ( .A(n1542), .B(n1922), .ZN(n772) );
  AOI221_X1 U1617 ( .B1(n1921), .B2(B[2]), .C1(n1920), .C2(B[1]), .A(n1923), 
        .ZN(n1922) );
  OAI22_X1 U1618 ( .A1(n1585), .A2(n1917), .B1(n1574), .B2(n1924), .ZN(n1923)
         );
  XNOR2_X1 U1619 ( .A(n1542), .B(n1925), .ZN(n771) );
  AOI221_X1 U1620 ( .B1(n1921), .B2(B[3]), .C1(n1920), .C2(B[2]), .A(n1926), 
        .ZN(n1925) );
  OAI22_X1 U1621 ( .A1(n1589), .A2(n1917), .B1(n1578), .B2(n1924), .ZN(n1926)
         );
  XNOR2_X1 U1622 ( .A(n1542), .B(n1927), .ZN(n770) );
  AOI221_X1 U1623 ( .B1(n1921), .B2(B[4]), .C1(n1920), .C2(B[3]), .A(n1928), 
        .ZN(n1927) );
  OAI22_X1 U1624 ( .A1(n1592), .A2(n1917), .B1(n1593), .B2(n1924), .ZN(n1928)
         );
  XNOR2_X1 U1625 ( .A(n1542), .B(n1929), .ZN(n769) );
  AOI221_X1 U1626 ( .B1(n1921), .B2(B[5]), .C1(n1920), .C2(B[4]), .A(n1930), 
        .ZN(n1929) );
  OAI22_X1 U1627 ( .A1(n1596), .A2(n1917), .B1(n1597), .B2(n1924), .ZN(n1930)
         );
  XNOR2_X1 U1628 ( .A(n1542), .B(n1931), .ZN(n768) );
  AOI221_X1 U1629 ( .B1(n1921), .B2(B[6]), .C1(n1920), .C2(B[5]), .A(n1932), 
        .ZN(n1931) );
  OAI22_X1 U1630 ( .A1(n1600), .A2(n1917), .B1(n1601), .B2(n1924), .ZN(n1932)
         );
  XNOR2_X1 U1631 ( .A(n1542), .B(n1933), .ZN(n767) );
  AOI221_X1 U1632 ( .B1(n1921), .B2(B[7]), .C1(n1920), .C2(B[6]), .A(n1934), 
        .ZN(n1933) );
  OAI22_X1 U1633 ( .A1(n1604), .A2(n1917), .B1(n1605), .B2(n1924), .ZN(n1934)
         );
  XNOR2_X1 U1634 ( .A(n1542), .B(n1935), .ZN(n766) );
  AOI221_X1 U1635 ( .B1(n1921), .B2(B[8]), .C1(n1920), .C2(B[7]), .A(n1936), 
        .ZN(n1935) );
  OAI22_X1 U1636 ( .A1(n1608), .A2(n1917), .B1(n1609), .B2(n1924), .ZN(n1936)
         );
  XNOR2_X1 U1637 ( .A(n1542), .B(n1937), .ZN(n765) );
  AOI221_X1 U1638 ( .B1(n1921), .B2(B[9]), .C1(n1920), .C2(B[8]), .A(n1938), 
        .ZN(n1937) );
  OAI22_X1 U1639 ( .A1(n1612), .A2(n1917), .B1(n1613), .B2(n1924), .ZN(n1938)
         );
  XNOR2_X1 U1640 ( .A(n1542), .B(n1939), .ZN(n764) );
  AOI221_X1 U1641 ( .B1(n1921), .B2(B[10]), .C1(n1920), .C2(B[9]), .A(n1940), 
        .ZN(n1939) );
  OAI22_X1 U1642 ( .A1(n1616), .A2(n1917), .B1(n1617), .B2(n1924), .ZN(n1940)
         );
  XNOR2_X1 U1643 ( .A(n1542), .B(n1941), .ZN(n763) );
  AOI221_X1 U1644 ( .B1(n1921), .B2(B[11]), .C1(n1920), .C2(B[10]), .A(n1942), 
        .ZN(n1941) );
  OAI22_X1 U1645 ( .A1(n1620), .A2(n1917), .B1(n1621), .B2(n1924), .ZN(n1942)
         );
  XNOR2_X1 U1646 ( .A(n1542), .B(n1943), .ZN(n762) );
  AOI221_X1 U1647 ( .B1(n1921), .B2(B[12]), .C1(n1920), .C2(B[11]), .A(n1944), 
        .ZN(n1943) );
  OAI22_X1 U1648 ( .A1(n1624), .A2(n1917), .B1(n1625), .B2(n1924), .ZN(n1944)
         );
  XNOR2_X1 U1649 ( .A(n1542), .B(n1945), .ZN(n761) );
  AOI221_X1 U1650 ( .B1(n1921), .B2(B[13]), .C1(n1920), .C2(B[12]), .A(n1946), 
        .ZN(n1945) );
  OAI22_X1 U1651 ( .A1(n1628), .A2(n1917), .B1(n1629), .B2(n1924), .ZN(n1946)
         );
  XNOR2_X1 U1652 ( .A(n1542), .B(n1947), .ZN(n760) );
  AOI221_X1 U1653 ( .B1(n1921), .B2(B[14]), .C1(n1920), .C2(B[13]), .A(n1948), 
        .ZN(n1947) );
  OAI22_X1 U1654 ( .A1(n1632), .A2(n1917), .B1(n1633), .B2(n1924), .ZN(n1948)
         );
  XNOR2_X1 U1655 ( .A(n1542), .B(n1949), .ZN(n759) );
  AOI221_X1 U1656 ( .B1(n1921), .B2(B[15]), .C1(n1920), .C2(B[14]), .A(n1950), 
        .ZN(n1949) );
  OAI22_X1 U1657 ( .A1(n1636), .A2(n1917), .B1(n1637), .B2(n1924), .ZN(n1950)
         );
  XNOR2_X1 U1658 ( .A(n1542), .B(n1951), .ZN(n758) );
  AOI221_X1 U1659 ( .B1(n1921), .B2(B[16]), .C1(n1920), .C2(B[15]), .A(n1952), 
        .ZN(n1951) );
  OAI22_X1 U1660 ( .A1(n1640), .A2(n1917), .B1(n1641), .B2(n1924), .ZN(n1952)
         );
  XNOR2_X1 U1661 ( .A(n1542), .B(n1953), .ZN(n757) );
  AOI221_X1 U1662 ( .B1(n1921), .B2(B[17]), .C1(n1920), .C2(B[16]), .A(n1954), 
        .ZN(n1953) );
  OAI22_X1 U1663 ( .A1(n1644), .A2(n1917), .B1(n1645), .B2(n1924), .ZN(n1954)
         );
  XNOR2_X1 U1664 ( .A(n1542), .B(n1955), .ZN(n756) );
  AOI221_X1 U1665 ( .B1(n1921), .B2(B[18]), .C1(n1920), .C2(B[17]), .A(n1956), 
        .ZN(n1955) );
  OAI22_X1 U1666 ( .A1(n1648), .A2(n1917), .B1(n1649), .B2(n1924), .ZN(n1956)
         );
  XNOR2_X1 U1667 ( .A(n1542), .B(n1957), .ZN(n755) );
  AOI221_X1 U1668 ( .B1(n1921), .B2(B[19]), .C1(n1920), .C2(B[18]), .A(n1958), 
        .ZN(n1957) );
  OAI22_X1 U1669 ( .A1(n1652), .A2(n1917), .B1(n1653), .B2(n1924), .ZN(n1958)
         );
  XNOR2_X1 U1670 ( .A(n1542), .B(n1959), .ZN(n754) );
  AOI221_X1 U1671 ( .B1(n1921), .B2(B[20]), .C1(n1920), .C2(B[19]), .A(n1960), 
        .ZN(n1959) );
  OAI22_X1 U1672 ( .A1(n1656), .A2(n1917), .B1(n1657), .B2(n1924), .ZN(n1960)
         );
  XNOR2_X1 U1673 ( .A(A[20]), .B(n1961), .ZN(n753) );
  AOI221_X1 U1674 ( .B1(n1921), .B2(B[21]), .C1(n1920), .C2(B[20]), .A(n1962), 
        .ZN(n1961) );
  OAI22_X1 U1675 ( .A1(n1660), .A2(n1917), .B1(n1661), .B2(n1924), .ZN(n1962)
         );
  XNOR2_X1 U1676 ( .A(A[20]), .B(n1963), .ZN(n752) );
  AOI221_X1 U1677 ( .B1(n1921), .B2(B[22]), .C1(n1920), .C2(B[21]), .A(n1964), 
        .ZN(n1963) );
  OAI22_X1 U1678 ( .A1(n1562), .A2(n1917), .B1(n1564), .B2(n1924), .ZN(n1964)
         );
  XNOR2_X1 U1679 ( .A(A[20]), .B(n1965), .ZN(n751) );
  AOI221_X1 U1680 ( .B1(n1921), .B2(n1554), .C1(n1920), .C2(B[22]), .A(n1966), 
        .ZN(n1965) );
  OAI22_X1 U1681 ( .A1(n1567), .A2(n1917), .B1(n1568), .B2(n1924), .ZN(n1966)
         );
  XNOR2_X1 U1682 ( .A(A[20]), .B(n1967), .ZN(n750) );
  AOI221_X1 U1683 ( .B1(n1921), .B2(B[23]), .C1(n1920), .C2(n1554), .A(n1968), 
        .ZN(n1967) );
  OAI22_X1 U1684 ( .A1(n1571), .A2(n1917), .B1(n1572), .B2(n1924), .ZN(n1968)
         );
  XNOR2_X1 U1685 ( .A(A[20]), .B(n1969), .ZN(n749) );
  OAI221_X1 U1686 ( .B1(n1556), .B2(n1924), .C1(n1556), .C2(n1917), .A(n1970), 
        .ZN(n1969) );
  OAI21_X1 U1687 ( .B1(n1921), .B2(n1920), .A(n1554), .ZN(n1970) );
  INV_X1 U1688 ( .A(n1974), .ZN(n1971) );
  XNOR2_X1 U1689 ( .A(A[18]), .B(A[19]), .ZN(n1972) );
  XNOR2_X1 U1690 ( .A(A[19]), .B(n1543), .ZN(n1973) );
  XOR2_X1 U1691 ( .A(A[18]), .B(n1545), .Z(n1974) );
  XNOR2_X1 U1692 ( .A(n1975), .B(n1541), .ZN(n748) );
  OAI22_X1 U1693 ( .A1(n1574), .A2(n1535), .B1(n1574), .B2(n1976), .ZN(n1975)
         );
  XNOR2_X1 U1694 ( .A(n1977), .B(n1541), .ZN(n747) );
  OAI222_X1 U1695 ( .A1(n1578), .A2(n1535), .B1(n1574), .B2(n1534), .C1(n1580), 
        .C2(n1976), .ZN(n1977) );
  INV_X1 U1696 ( .A(n1397), .ZN(n1580) );
  XNOR2_X1 U1697 ( .A(n1540), .B(n1978), .ZN(n746) );
  AOI221_X1 U1698 ( .B1(n1537), .B2(B[2]), .C1(n1536), .C2(B[1]), .A(n1979), 
        .ZN(n1978) );
  OAI22_X1 U1699 ( .A1(n1585), .A2(n1976), .B1(n1574), .B2(n1538), .ZN(n1979)
         );
  INV_X1 U1700 ( .A(n1396), .ZN(n1585) );
  XNOR2_X1 U1701 ( .A(n1540), .B(n1981), .ZN(n745) );
  AOI221_X1 U1702 ( .B1(n1537), .B2(B[3]), .C1(n1536), .C2(B[2]), .A(n1982), 
        .ZN(n1981) );
  OAI22_X1 U1703 ( .A1(n1589), .A2(n1976), .B1(n1578), .B2(n1539), .ZN(n1982)
         );
  XNOR2_X1 U1704 ( .A(n1540), .B(n1983), .ZN(n744) );
  AOI221_X1 U1705 ( .B1(n1537), .B2(B[4]), .C1(n1536), .C2(B[3]), .A(n1984), 
        .ZN(n1983) );
  OAI22_X1 U1706 ( .A1(n1592), .A2(n1976), .B1(n1593), .B2(n1539), .ZN(n1984)
         );
  XNOR2_X1 U1707 ( .A(n1540), .B(n1985), .ZN(n743) );
  AOI221_X1 U1708 ( .B1(n1537), .B2(B[5]), .C1(n1536), .C2(B[4]), .A(n1986), 
        .ZN(n1985) );
  OAI22_X1 U1709 ( .A1(n1596), .A2(n1976), .B1(n1597), .B2(n1539), .ZN(n1986)
         );
  XNOR2_X1 U1710 ( .A(n1540), .B(n1987), .ZN(n742) );
  AOI221_X1 U1711 ( .B1(n1537), .B2(B[6]), .C1(n1536), .C2(B[5]), .A(n1988), 
        .ZN(n1987) );
  OAI22_X1 U1712 ( .A1(n1600), .A2(n1976), .B1(n1601), .B2(n1539), .ZN(n1988)
         );
  XNOR2_X1 U1713 ( .A(n1540), .B(n1989), .ZN(n741) );
  AOI221_X1 U1714 ( .B1(n1537), .B2(B[7]), .C1(n1536), .C2(B[6]), .A(n1990), 
        .ZN(n1989) );
  OAI22_X1 U1715 ( .A1(n1604), .A2(n1976), .B1(n1605), .B2(n1539), .ZN(n1990)
         );
  XNOR2_X1 U1716 ( .A(n1540), .B(n1991), .ZN(n740) );
  AOI221_X1 U1717 ( .B1(n1537), .B2(B[9]), .C1(n1536), .C2(B[8]), .A(n1992), 
        .ZN(n1991) );
  OAI22_X1 U1718 ( .A1(n1612), .A2(n1976), .B1(n1613), .B2(n1539), .ZN(n1992)
         );
  XNOR2_X1 U1719 ( .A(n1540), .B(n1993), .ZN(n739) );
  AOI221_X1 U1720 ( .B1(n1537), .B2(B[10]), .C1(n1536), .C2(B[9]), .A(n1994), 
        .ZN(n1993) );
  OAI22_X1 U1721 ( .A1(n1616), .A2(n1976), .B1(n1617), .B2(n1539), .ZN(n1994)
         );
  XNOR2_X1 U1722 ( .A(n1540), .B(n1995), .ZN(n738) );
  AOI221_X1 U1723 ( .B1(n1537), .B2(B[12]), .C1(n1536), .C2(B[11]), .A(n1996), 
        .ZN(n1995) );
  OAI22_X1 U1724 ( .A1(n1624), .A2(n1976), .B1(n1625), .B2(n1539), .ZN(n1996)
         );
  XNOR2_X1 U1725 ( .A(n1540), .B(n1997), .ZN(n737) );
  AOI221_X1 U1726 ( .B1(n1537), .B2(B[13]), .C1(n1536), .C2(B[12]), .A(n1998), 
        .ZN(n1997) );
  OAI22_X1 U1727 ( .A1(n1628), .A2(n1976), .B1(n1629), .B2(n1539), .ZN(n1998)
         );
  XNOR2_X1 U1728 ( .A(n1540), .B(n1999), .ZN(n736) );
  AOI221_X1 U1729 ( .B1(n1537), .B2(B[14]), .C1(n1536), .C2(B[13]), .A(n2000), 
        .ZN(n1999) );
  OAI22_X1 U1730 ( .A1(n1632), .A2(n1976), .B1(n1633), .B2(n1539), .ZN(n2000)
         );
  XNOR2_X1 U1731 ( .A(n1540), .B(n2001), .ZN(n735) );
  AOI221_X1 U1732 ( .B1(n1537), .B2(B[15]), .C1(n1536), .C2(B[14]), .A(n2002), 
        .ZN(n2001) );
  OAI22_X1 U1733 ( .A1(n1636), .A2(n1976), .B1(n1637), .B2(n1539), .ZN(n2002)
         );
  XNOR2_X1 U1734 ( .A(n1540), .B(n2003), .ZN(n734) );
  AOI221_X1 U1735 ( .B1(n1537), .B2(B[16]), .C1(n1536), .C2(B[15]), .A(n2004), 
        .ZN(n2003) );
  OAI22_X1 U1736 ( .A1(n1640), .A2(n1976), .B1(n1641), .B2(n1538), .ZN(n2004)
         );
  XNOR2_X1 U1737 ( .A(n1540), .B(n2005), .ZN(n733) );
  AOI221_X1 U1738 ( .B1(n1537), .B2(B[18]), .C1(n1536), .C2(B[17]), .A(n2006), 
        .ZN(n2005) );
  OAI22_X1 U1739 ( .A1(n1648), .A2(n1976), .B1(n1649), .B2(n1538), .ZN(n2006)
         );
  XNOR2_X1 U1740 ( .A(n1540), .B(n2007), .ZN(n732) );
  AOI221_X1 U1741 ( .B1(n1537), .B2(B[19]), .C1(n1536), .C2(B[18]), .A(n2008), 
        .ZN(n2007) );
  OAI22_X1 U1742 ( .A1(n1652), .A2(n1976), .B1(n1653), .B2(n1538), .ZN(n2008)
         );
  XNOR2_X1 U1743 ( .A(n1540), .B(n2009), .ZN(n731) );
  AOI221_X1 U1744 ( .B1(n1537), .B2(B[20]), .C1(n1536), .C2(B[19]), .A(n2010), 
        .ZN(n2009) );
  OAI22_X1 U1745 ( .A1(n1656), .A2(n1976), .B1(n1657), .B2(n1538), .ZN(n2010)
         );
  XNOR2_X1 U1746 ( .A(A[23]), .B(n2011), .ZN(n730) );
  AOI221_X1 U1747 ( .B1(n1537), .B2(B[21]), .C1(n1536), .C2(B[20]), .A(n2012), 
        .ZN(n2011) );
  OAI22_X1 U1748 ( .A1(n1660), .A2(n1976), .B1(n1661), .B2(n1538), .ZN(n2012)
         );
  XNOR2_X1 U1749 ( .A(A[23]), .B(n2013), .ZN(n729) );
  AOI221_X1 U1750 ( .B1(n1537), .B2(B[22]), .C1(n1536), .C2(B[21]), .A(n2014), 
        .ZN(n2013) );
  OAI22_X1 U1751 ( .A1(n1562), .A2(n1976), .B1(n1564), .B2(n1538), .ZN(n2014)
         );
  INV_X1 U1752 ( .A(B[20]), .ZN(n1564) );
  INV_X1 U1753 ( .A(n1376), .ZN(n1562) );
  XNOR2_X1 U1754 ( .A(n519), .B(n2015), .ZN(n506) );
  INV_X1 U1755 ( .A(n493), .ZN(n479) );
  NOR2_X1 U1756 ( .A1(n2015), .A2(n519), .ZN(n493) );
  XOR2_X1 U1757 ( .A(n2016), .B(n1674), .Z(n2015) );
  OAI221_X1 U1758 ( .B1(n1563), .B2(n1556), .C1(n1561), .C2(n1556), .A(n2017), 
        .ZN(n2016) );
  OAI21_X1 U1759 ( .B1(n1558), .B2(n1559), .A(n1554), .ZN(n2017) );
  INV_X1 U1760 ( .A(n454), .ZN(n442) );
  XOR2_X1 U1761 ( .A(n1540), .B(n2018), .Z(n454) );
  AOI221_X1 U1762 ( .B1(n1537), .B2(B[8]), .C1(n1536), .C2(B[7]), .A(n2019), 
        .ZN(n2018) );
  OAI22_X1 U1763 ( .A1(n1608), .A2(n1976), .B1(n1609), .B2(n1538), .ZN(n2019)
         );
  INV_X1 U1764 ( .A(n421), .ZN(n411) );
  XOR2_X1 U1765 ( .A(n1540), .B(n2020), .Z(n421) );
  AOI221_X1 U1766 ( .B1(n1537), .B2(B[11]), .C1(n1536), .C2(B[10]), .A(n2021), 
        .ZN(n2020) );
  OAI22_X1 U1767 ( .A1(n1620), .A2(n1976), .B1(n1621), .B2(n1538), .ZN(n2021)
         );
  INV_X1 U1768 ( .A(n387), .ZN(n395) );
  INV_X1 U1769 ( .A(n374), .ZN(n368) );
  XOR2_X1 U1770 ( .A(n1540), .B(n2022), .Z(n374) );
  AOI221_X1 U1771 ( .B1(n1537), .B2(B[17]), .C1(n1536), .C2(B[16]), .A(n2023), 
        .ZN(n2022) );
  OAI22_X1 U1772 ( .A1(n1644), .A2(n1976), .B1(n1645), .B2(n1538), .ZN(n2023)
         );
  INV_X1 U1773 ( .A(n356), .ZN(n360) );
  INV_X1 U1774 ( .A(n2024), .ZN(n351) );
  OAI222_X1 U1775 ( .A1(n2025), .A2(n2026), .B1(n2025), .B2(n2027), .C1(n2027), 
        .C2(n2026), .ZN(n326) );
  INV_X1 U1776 ( .A(n550), .ZN(n2027) );
  XNOR2_X1 U1777 ( .A(n1674), .B(n2028), .ZN(n2026) );
  AOI221_X1 U1778 ( .B1(B[21]), .B2(n1558), .C1(B[20]), .C2(n1559), .A(n2029), 
        .ZN(n2028) );
  OAI22_X1 U1779 ( .A1(n1561), .A2(n1660), .B1(n1563), .B2(n1661), .ZN(n2029)
         );
  INV_X1 U1780 ( .A(B[19]), .ZN(n1661) );
  INV_X1 U1781 ( .A(n1377), .ZN(n1660) );
  AOI222_X1 U1782 ( .A1(n2030), .A2(n2031), .B1(n2030), .B2(n564), .C1(n564), 
        .C2(n2031), .ZN(n2025) );
  XNOR2_X1 U1783 ( .A(A[2]), .B(n2032), .ZN(n2031) );
  AOI221_X1 U1784 ( .B1(B[20]), .B2(n1558), .C1(B[19]), .C2(n1559), .A(n2033), 
        .ZN(n2032) );
  OAI22_X1 U1785 ( .A1(n1561), .A2(n1656), .B1(n1563), .B2(n1657), .ZN(n2033)
         );
  INV_X1 U1786 ( .A(B[18]), .ZN(n1657) );
  INV_X1 U1787 ( .A(n1378), .ZN(n1656) );
  INV_X1 U1788 ( .A(n2034), .ZN(n2030) );
  AOI222_X1 U1789 ( .A1(n2035), .A2(n2036), .B1(n2035), .B2(n576), .C1(n576), 
        .C2(n2036), .ZN(n2034) );
  XNOR2_X1 U1790 ( .A(A[2]), .B(n2037), .ZN(n2036) );
  AOI221_X1 U1791 ( .B1(B[19]), .B2(n1558), .C1(B[18]), .C2(n1559), .A(n2038), 
        .ZN(n2037) );
  OAI22_X1 U1792 ( .A1(n1561), .A2(n1652), .B1(n1563), .B2(n1653), .ZN(n2038)
         );
  INV_X1 U1793 ( .A(B[17]), .ZN(n1653) );
  INV_X1 U1794 ( .A(n1379), .ZN(n1652) );
  OAI222_X1 U1795 ( .A1(n2039), .A2(n2040), .B1(n2039), .B2(n2041), .C1(n2041), 
        .C2(n2040), .ZN(n2035) );
  INV_X1 U1796 ( .A(n588), .ZN(n2041) );
  XNOR2_X1 U1797 ( .A(n1674), .B(n2042), .ZN(n2040) );
  AOI221_X1 U1798 ( .B1(B[18]), .B2(n1558), .C1(B[17]), .C2(n1559), .A(n2043), 
        .ZN(n2042) );
  OAI22_X1 U1799 ( .A1(n1561), .A2(n1648), .B1(n1563), .B2(n1649), .ZN(n2043)
         );
  INV_X1 U1800 ( .A(B[16]), .ZN(n1649) );
  INV_X1 U1801 ( .A(n1380), .ZN(n1648) );
  AOI222_X1 U1802 ( .A1(n2044), .A2(n2045), .B1(n2044), .B2(n600), .C1(n600), 
        .C2(n2045), .ZN(n2039) );
  XNOR2_X1 U1803 ( .A(A[2]), .B(n2046), .ZN(n2045) );
  AOI221_X1 U1804 ( .B1(B[17]), .B2(n1558), .C1(B[16]), .C2(n1559), .A(n2047), 
        .ZN(n2046) );
  OAI22_X1 U1805 ( .A1(n1561), .A2(n1644), .B1(n1563), .B2(n1645), .ZN(n2047)
         );
  INV_X1 U1806 ( .A(B[15]), .ZN(n1645) );
  INV_X1 U1807 ( .A(n1381), .ZN(n1644) );
  OAI222_X1 U1808 ( .A1(n2048), .A2(n2049), .B1(n2048), .B2(n2050), .C1(n2050), 
        .C2(n2049), .ZN(n2044) );
  INV_X1 U1809 ( .A(n610), .ZN(n2050) );
  XNOR2_X1 U1810 ( .A(n1674), .B(n2051), .ZN(n2049) );
  AOI221_X1 U1811 ( .B1(B[16]), .B2(n1558), .C1(B[15]), .C2(n1559), .A(n2052), 
        .ZN(n2051) );
  OAI22_X1 U1812 ( .A1(n1561), .A2(n1640), .B1(n1563), .B2(n1641), .ZN(n2052)
         );
  INV_X1 U1813 ( .A(B[14]), .ZN(n1641) );
  INV_X1 U1814 ( .A(n1382), .ZN(n1640) );
  AOI222_X1 U1815 ( .A1(n2053), .A2(n2054), .B1(n2053), .B2(n620), .C1(n620), 
        .C2(n2054), .ZN(n2048) );
  XNOR2_X1 U1816 ( .A(A[2]), .B(n2055), .ZN(n2054) );
  AOI221_X1 U1817 ( .B1(B[15]), .B2(n1558), .C1(B[14]), .C2(n1559), .A(n2056), 
        .ZN(n2055) );
  OAI22_X1 U1818 ( .A1(n1561), .A2(n1636), .B1(n1563), .B2(n1637), .ZN(n2056)
         );
  INV_X1 U1819 ( .A(B[13]), .ZN(n1637) );
  INV_X1 U1820 ( .A(n1383), .ZN(n1636) );
  OAI222_X1 U1821 ( .A1(n2057), .A2(n2058), .B1(n2057), .B2(n2059), .C1(n2059), 
        .C2(n2058), .ZN(n2053) );
  INV_X1 U1822 ( .A(n630), .ZN(n2059) );
  XNOR2_X1 U1823 ( .A(n1674), .B(n2060), .ZN(n2058) );
  AOI221_X1 U1824 ( .B1(B[14]), .B2(n1558), .C1(B[13]), .C2(n1559), .A(n2061), 
        .ZN(n2060) );
  OAI22_X1 U1825 ( .A1(n1561), .A2(n1632), .B1(n1563), .B2(n1633), .ZN(n2061)
         );
  INV_X1 U1826 ( .A(B[12]), .ZN(n1633) );
  INV_X1 U1827 ( .A(n1384), .ZN(n1632) );
  AOI222_X1 U1828 ( .A1(n2062), .A2(n2063), .B1(n2062), .B2(n638), .C1(n638), 
        .C2(n2063), .ZN(n2057) );
  XNOR2_X1 U1829 ( .A(A[2]), .B(n2064), .ZN(n2063) );
  AOI221_X1 U1830 ( .B1(B[13]), .B2(n1558), .C1(B[12]), .C2(n1559), .A(n2065), 
        .ZN(n2064) );
  OAI22_X1 U1831 ( .A1(n1561), .A2(n1628), .B1(n1563), .B2(n1629), .ZN(n2065)
         );
  INV_X1 U1832 ( .A(B[11]), .ZN(n1629) );
  INV_X1 U1833 ( .A(n1385), .ZN(n1628) );
  OAI222_X1 U1834 ( .A1(n2066), .A2(n2067), .B1(n2066), .B2(n2068), .C1(n2068), 
        .C2(n2067), .ZN(n2062) );
  INV_X1 U1835 ( .A(n646), .ZN(n2068) );
  XNOR2_X1 U1836 ( .A(n1674), .B(n2069), .ZN(n2067) );
  AOI221_X1 U1837 ( .B1(B[12]), .B2(n1558), .C1(B[11]), .C2(n1559), .A(n2070), 
        .ZN(n2069) );
  OAI22_X1 U1838 ( .A1(n1561), .A2(n1624), .B1(n1563), .B2(n1625), .ZN(n2070)
         );
  INV_X1 U1839 ( .A(B[10]), .ZN(n1625) );
  INV_X1 U1840 ( .A(n1386), .ZN(n1624) );
  AOI222_X1 U1841 ( .A1(n2071), .A2(n2072), .B1(n2071), .B2(n654), .C1(n654), 
        .C2(n2072), .ZN(n2066) );
  XNOR2_X1 U1842 ( .A(A[2]), .B(n2073), .ZN(n2072) );
  AOI221_X1 U1843 ( .B1(B[11]), .B2(n1558), .C1(B[10]), .C2(n1559), .A(n2074), 
        .ZN(n2073) );
  OAI22_X1 U1844 ( .A1(n1561), .A2(n1620), .B1(n1563), .B2(n1621), .ZN(n2074)
         );
  INV_X1 U1845 ( .A(B[9]), .ZN(n1621) );
  INV_X1 U1846 ( .A(n1387), .ZN(n1620) );
  OAI222_X1 U1847 ( .A1(n2075), .A2(n2076), .B1(n2075), .B2(n2077), .C1(n2077), 
        .C2(n2076), .ZN(n2071) );
  INV_X1 U1848 ( .A(n660), .ZN(n2077) );
  XNOR2_X1 U1849 ( .A(n1674), .B(n2078), .ZN(n2076) );
  AOI221_X1 U1850 ( .B1(B[10]), .B2(n1558), .C1(B[9]), .C2(n1559), .A(n2079), 
        .ZN(n2078) );
  OAI22_X1 U1851 ( .A1(n1561), .A2(n1616), .B1(n1563), .B2(n1617), .ZN(n2079)
         );
  INV_X1 U1852 ( .A(B[8]), .ZN(n1617) );
  INV_X1 U1853 ( .A(n1388), .ZN(n1616) );
  AOI222_X1 U1854 ( .A1(n2080), .A2(n2081), .B1(n2080), .B2(n666), .C1(n666), 
        .C2(n2081), .ZN(n2075) );
  XNOR2_X1 U1855 ( .A(A[2]), .B(n2082), .ZN(n2081) );
  AOI221_X1 U1856 ( .B1(B[9]), .B2(n1558), .C1(B[8]), .C2(n1559), .A(n2083), 
        .ZN(n2082) );
  OAI22_X1 U1857 ( .A1(n1561), .A2(n1612), .B1(n1563), .B2(n1613), .ZN(n2083)
         );
  INV_X1 U1858 ( .A(B[7]), .ZN(n1613) );
  INV_X1 U1859 ( .A(n1389), .ZN(n1612) );
  OAI222_X1 U1860 ( .A1(n2084), .A2(n2085), .B1(n2084), .B2(n2086), .C1(n2086), 
        .C2(n2085), .ZN(n2080) );
  INV_X1 U1861 ( .A(n672), .ZN(n2086) );
  XNOR2_X1 U1862 ( .A(n1674), .B(n2087), .ZN(n2085) );
  AOI221_X1 U1863 ( .B1(B[8]), .B2(n1558), .C1(B[7]), .C2(n1559), .A(n2088), 
        .ZN(n2087) );
  OAI22_X1 U1864 ( .A1(n1561), .A2(n1608), .B1(n1563), .B2(n1609), .ZN(n2088)
         );
  INV_X1 U1865 ( .A(B[6]), .ZN(n1609) );
  INV_X1 U1866 ( .A(n1390), .ZN(n1608) );
  AOI222_X1 U1867 ( .A1(n2089), .A2(n2090), .B1(n2089), .B2(n676), .C1(n676), 
        .C2(n2090), .ZN(n2084) );
  XNOR2_X1 U1868 ( .A(A[2]), .B(n2091), .ZN(n2090) );
  AOI221_X1 U1869 ( .B1(B[7]), .B2(n1558), .C1(B[6]), .C2(n1559), .A(n2092), 
        .ZN(n2091) );
  OAI22_X1 U1870 ( .A1(n1561), .A2(n1604), .B1(n1563), .B2(n1605), .ZN(n2092)
         );
  INV_X1 U1871 ( .A(B[5]), .ZN(n1605) );
  INV_X1 U1872 ( .A(n1391), .ZN(n1604) );
  OAI222_X1 U1873 ( .A1(n2093), .A2(n2094), .B1(n2093), .B2(n2095), .C1(n2095), 
        .C2(n2094), .ZN(n2089) );
  INV_X1 U1874 ( .A(n680), .ZN(n2095) );
  XNOR2_X1 U1875 ( .A(n1674), .B(n2096), .ZN(n2094) );
  AOI221_X1 U1876 ( .B1(B[6]), .B2(n1558), .C1(B[5]), .C2(n1559), .A(n2097), 
        .ZN(n2096) );
  OAI22_X1 U1877 ( .A1(n1561), .A2(n1600), .B1(n1563), .B2(n1601), .ZN(n2097)
         );
  INV_X1 U1878 ( .A(B[4]), .ZN(n1601) );
  INV_X1 U1879 ( .A(n1392), .ZN(n1600) );
  AOI222_X1 U1880 ( .A1(n2098), .A2(n2099), .B1(n2098), .B2(n684), .C1(n684), 
        .C2(n2099), .ZN(n2093) );
  XNOR2_X1 U1881 ( .A(A[2]), .B(n2100), .ZN(n2099) );
  AOI221_X1 U1882 ( .B1(B[5]), .B2(n1558), .C1(B[4]), .C2(n1559), .A(n2101), 
        .ZN(n2100) );
  OAI22_X1 U1883 ( .A1(n1561), .A2(n1596), .B1(n1563), .B2(n1597), .ZN(n2101)
         );
  INV_X1 U1884 ( .A(B[3]), .ZN(n1597) );
  INV_X1 U1885 ( .A(n1393), .ZN(n1596) );
  OAI222_X1 U1886 ( .A1(n2102), .A2(n2103), .B1(n2102), .B2(n2104), .C1(n2104), 
        .C2(n2103), .ZN(n2098) );
  INV_X1 U1887 ( .A(n686), .ZN(n2104) );
  XNOR2_X1 U1888 ( .A(n1674), .B(n2105), .ZN(n2103) );
  AOI221_X1 U1889 ( .B1(B[4]), .B2(n1558), .C1(B[3]), .C2(n1559), .A(n2106), 
        .ZN(n2105) );
  OAI22_X1 U1890 ( .A1(n1561), .A2(n1592), .B1(n1563), .B2(n1593), .ZN(n2106)
         );
  INV_X1 U1891 ( .A(B[2]), .ZN(n1593) );
  INV_X1 U1892 ( .A(n1394), .ZN(n1592) );
  AOI222_X1 U1893 ( .A1(n2107), .A2(n2108), .B1(n2107), .B2(n688), .C1(n688), 
        .C2(n2108), .ZN(n2102) );
  XNOR2_X1 U1894 ( .A(A[2]), .B(n2109), .ZN(n2108) );
  AOI221_X1 U1895 ( .B1(B[3]), .B2(n1558), .C1(B[2]), .C2(n1559), .A(n2110), 
        .ZN(n2109) );
  OAI22_X1 U1896 ( .A1(n1561), .A2(n1589), .B1(n1563), .B2(n1578), .ZN(n2110)
         );
  INV_X1 U1897 ( .A(B[1]), .ZN(n1578) );
  INV_X1 U1898 ( .A(n1395), .ZN(n1589) );
  AND2_X1 U1899 ( .A1(n2114), .A2(n2115), .ZN(n2107) );
  AOI211_X1 U1900 ( .C1(B[1]), .C2(n1558), .A(n2116), .B(B[0]), .ZN(n2115) );
  INV_X1 U1901 ( .A(n2117), .ZN(n2116) );
  AOI22_X1 U1902 ( .A1(n1558), .A2(B[2]), .B1(n2118), .B2(n1397), .ZN(n2117)
         );
  INV_X1 U1903 ( .A(A[0]), .ZN(n2112) );
  AOI221_X1 U1904 ( .B1(B[1]), .B2(n1559), .C1(n1396), .C2(n2118), .A(n1674), 
        .ZN(n2114) );
  INV_X1 U1905 ( .A(n1561), .ZN(n2118) );
  XNOR2_X1 U1906 ( .A(A[1]), .B(n1674), .ZN(n2111) );
  INV_X1 U1907 ( .A(A[2]), .ZN(n1674) );
  INV_X1 U1908 ( .A(A[1]), .ZN(n2113) );
  AOI21_X1 U1909 ( .B1(n2119), .B2(n2120), .A(n2121), .ZN(PRODUCT[47]) );
  OAI22_X1 U1910 ( .A1(n2122), .A2(n2123), .B1(n2122), .B2(n2124), .ZN(n2121)
         );
  INV_X1 U1911 ( .A(n2120), .ZN(n2124) );
  AOI222_X1 U1912 ( .A1(n2024), .A2(n303), .B1(n2123), .B2(n303), .C1(n2024), 
        .C2(n2123), .ZN(n2122) );
  XOR2_X1 U1913 ( .A(n1541), .B(n2125), .Z(n2024) );
  AOI221_X1 U1914 ( .B1(n1537), .B2(B[23]), .C1(n1536), .C2(B[22]), .A(n2126), 
        .ZN(n2125) );
  OAI22_X1 U1915 ( .A1(n1567), .A2(n1976), .B1(n1568), .B2(n1538), .ZN(n2126)
         );
  INV_X1 U1916 ( .A(B[21]), .ZN(n1568) );
  INV_X1 U1917 ( .A(n1375), .ZN(n1567) );
  XOR2_X1 U1918 ( .A(n2127), .B(n1541), .Z(n2120) );
  OAI221_X1 U1919 ( .B1(n1556), .B2(n1539), .C1(n1556), .C2(n1976), .A(n2128), 
        .ZN(n2127) );
  OAI21_X1 U1920 ( .B1(n1537), .B2(n1536), .A(n1554), .ZN(n2128) );
  INV_X1 U1921 ( .A(n2123), .ZN(n2119) );
  XOR2_X1 U1922 ( .A(A[23]), .B(n2129), .Z(n2123) );
  AOI221_X1 U1923 ( .B1(n1537), .B2(n1554), .C1(n1536), .C2(n1554), .A(n2130), 
        .ZN(n2129) );
  OAI22_X1 U1924 ( .A1(n1571), .A2(n1976), .B1(n1572), .B2(n1538), .ZN(n2130)
         );
  NAND3_X1 U1925 ( .A1(n2131), .A2(n2132), .A3(n2133), .ZN(n1980) );
  INV_X1 U1926 ( .A(B[22]), .ZN(n1572) );
  INV_X1 U1927 ( .A(n1374), .ZN(n1571) );
  XNOR2_X1 U1928 ( .A(A[21]), .B(A[22]), .ZN(n2133) );
  INV_X1 U1929 ( .A(n2131), .ZN(n2134) );
  XOR2_X1 U1930 ( .A(A[21]), .B(n1543), .Z(n2131) );
  XNOR2_X1 U1931 ( .A(A[22]), .B(n1541), .ZN(n2132) );
endmodule


module iir_filter_DW02_mult_2 ( A, B, PRODUCT, TC );
  input [23:0] A;
  input [23:0] B;
  output [47:0] PRODUCT;
  input TC;
  wire   n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n351, n352, n353, n354, n355, n356, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n906, n907, n908, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134;

  FA_X1 U182 ( .A(n351), .B(n352), .CI(n304), .CO(n303), .S(PRODUCT[44]) );
  FA_X1 U183 ( .A(n353), .B(n354), .CI(n305), .CO(n304), .S(PRODUCT[43]) );
  FA_X1 U184 ( .A(n355), .B(n358), .CI(n306), .CO(n305), .S(PRODUCT[42]) );
  FA_X1 U185 ( .A(n359), .B(n361), .CI(n307), .CO(n306), .S(PRODUCT[41]) );
  FA_X1 U186 ( .A(n362), .B(n364), .CI(n308), .CO(n307), .S(PRODUCT[40]) );
  FA_X1 U187 ( .A(n365), .B(n370), .CI(n309), .CO(n308), .S(PRODUCT[39]) );
  FA_X1 U188 ( .A(n371), .B(n375), .CI(n310), .CO(n309), .S(PRODUCT[38]) );
  FA_X1 U189 ( .A(n376), .B(n381), .CI(n311), .CO(n310), .S(PRODUCT[37]) );
  FA_X1 U190 ( .A(n382), .B(n389), .CI(n312), .CO(n311), .S(PRODUCT[36]) );
  FA_X1 U191 ( .A(n390), .B(n396), .CI(n313), .CO(n312), .S(PRODUCT[35]) );
  FA_X1 U192 ( .A(n397), .B(n403), .CI(n314), .CO(n313), .S(PRODUCT[34]) );
  FA_X1 U193 ( .A(n404), .B(n413), .CI(n315), .CO(n314), .S(PRODUCT[33]) );
  FA_X1 U194 ( .A(n414), .B(n422), .CI(n316), .CO(n315), .S(PRODUCT[32]) );
  FA_X1 U195 ( .A(n423), .B(n432), .CI(n317), .CO(n316), .S(PRODUCT[31]) );
  FA_X1 U196 ( .A(n433), .B(n444), .CI(n318), .CO(n317), .S(PRODUCT[30]) );
  FA_X1 U197 ( .A(n445), .B(n455), .CI(n319), .CO(n318), .S(PRODUCT[29]) );
  FA_X1 U198 ( .A(n456), .B(n467), .CI(n320), .CO(n319), .S(PRODUCT[28]) );
  FA_X1 U199 ( .A(n468), .B(n481), .CI(n321), .CO(n320), .S(PRODUCT[27]) );
  FA_X1 U200 ( .A(n482), .B(n494), .CI(n322), .CO(n321), .S(PRODUCT[26]) );
  FA_X1 U201 ( .A(n495), .B(n507), .CI(n323), .CO(n322), .S(PRODUCT[25]) );
  FA_X1 U202 ( .A(n508), .B(n906), .CI(n324), .CO(n323), .S(PRODUCT[24]) );
  FA_X1 U203 ( .A(n907), .B(n522), .CI(n325), .CO(n324), .S(PRODUCT[23]) );
  FA_X1 U204 ( .A(n908), .B(n536), .CI(n326), .CO(n325), .S(PRODUCT[22]) );
  FA_X1 U235 ( .A(n356), .B(n749), .CI(n729), .CO(n352), .S(n353) );
  FA_X1 U236 ( .A(n730), .B(n360), .CI(n750), .CO(n354), .S(n355) );
  FA_X1 U238 ( .A(n360), .B(n731), .CI(n751), .CO(n358), .S(n359) );
  FA_X1 U240 ( .A(n752), .B(n363), .CI(n366), .CO(n361), .S(n362) );
  FA_X1 U241 ( .A(n368), .B(n775), .CI(n732), .CO(n356), .S(n363) );
  FA_X1 U242 ( .A(n776), .B(n753), .CI(n367), .CO(n364), .S(n365) );
  FA_X1 U243 ( .A(n733), .B(n374), .CI(n372), .CO(n366), .S(n367) );
  FA_X1 U245 ( .A(n373), .B(n377), .CI(n777), .CO(n370), .S(n371) );
  FA_X1 U246 ( .A(n374), .B(n379), .CI(n754), .CO(n372), .S(n373) );
  FA_X1 U248 ( .A(n778), .B(n378), .CI(n383), .CO(n375), .S(n376) );
  FA_X1 U249 ( .A(n385), .B(n380), .CI(n755), .CO(n377), .S(n378) );
  FA_X1 U250 ( .A(n387), .B(n801), .CI(n734), .CO(n379), .S(n380) );
  FA_X1 U251 ( .A(n802), .B(n779), .CI(n384), .CO(n381), .S(n382) );
  FA_X1 U252 ( .A(n386), .B(n393), .CI(n391), .CO(n383), .S(n384) );
  FA_X1 U253 ( .A(n735), .B(n395), .CI(n756), .CO(n385), .S(n386) );
  FA_X1 U255 ( .A(n392), .B(n398), .CI(n803), .CO(n389), .S(n390) );
  FA_X1 U256 ( .A(n394), .B(n400), .CI(n780), .CO(n391), .S(n392) );
  FA_X1 U257 ( .A(n395), .B(n736), .CI(n757), .CO(n393), .S(n394) );
  FA_X1 U259 ( .A(n804), .B(n399), .CI(n405), .CO(n396), .S(n397) );
  FA_X1 U260 ( .A(n407), .B(n401), .CI(n781), .CO(n398), .S(n399) );
  FA_X1 U261 ( .A(n758), .B(n402), .CI(n409), .CO(n400), .S(n401) );
  FA_X1 U262 ( .A(n411), .B(n827), .CI(n737), .CO(n387), .S(n402) );
  FA_X1 U263 ( .A(n828), .B(n805), .CI(n406), .CO(n403), .S(n404) );
  FA_X1 U264 ( .A(n408), .B(n417), .CI(n415), .CO(n405), .S(n406) );
  FA_X1 U265 ( .A(n410), .B(n759), .CI(n782), .CO(n407), .S(n408) );
  FA_X1 U266 ( .A(n738), .B(n421), .CI(n419), .CO(n409), .S(n410) );
  FA_X1 U268 ( .A(n416), .B(n424), .CI(n829), .CO(n413), .S(n414) );
  FA_X1 U269 ( .A(n418), .B(n426), .CI(n806), .CO(n415), .S(n416) );
  FA_X1 U270 ( .A(n420), .B(n428), .CI(n783), .CO(n417), .S(n418) );
  FA_X1 U271 ( .A(n421), .B(n430), .CI(n760), .CO(n419), .S(n420) );
  FA_X1 U273 ( .A(n830), .B(n425), .CI(n434), .CO(n422), .S(n423) );
  FA_X1 U274 ( .A(n436), .B(n427), .CI(n807), .CO(n424), .S(n425) );
  FA_X1 U275 ( .A(n784), .B(n429), .CI(n438), .CO(n426), .S(n427) );
  FA_X1 U276 ( .A(n440), .B(n431), .CI(n761), .CO(n428), .S(n429) );
  FA_X1 U277 ( .A(n442), .B(n853), .CI(n739), .CO(n430), .S(n431) );
  FA_X1 U278 ( .A(n854), .B(n831), .CI(n435), .CO(n432), .S(n433) );
  FA_X1 U279 ( .A(n437), .B(n448), .CI(n446), .CO(n434), .S(n435) );
  FA_X1 U280 ( .A(n439), .B(n785), .CI(n808), .CO(n436), .S(n437) );
  FA_X1 U281 ( .A(n441), .B(n452), .CI(n450), .CO(n438), .S(n439) );
  FA_X1 U282 ( .A(n740), .B(n454), .CI(n762), .CO(n440), .S(n441) );
  FA_X1 U284 ( .A(n447), .B(n457), .CI(n855), .CO(n444), .S(n445) );
  FA_X1 U285 ( .A(n449), .B(n459), .CI(n832), .CO(n446), .S(n447) );
  FA_X1 U286 ( .A(n451), .B(n461), .CI(n809), .CO(n448), .S(n449) );
  FA_X1 U287 ( .A(n453), .B(n463), .CI(n786), .CO(n450), .S(n451) );
  FA_X1 U288 ( .A(n454), .B(n465), .CI(n763), .CO(n452), .S(n453) );
  FA_X1 U290 ( .A(n856), .B(n458), .CI(n469), .CO(n455), .S(n456) );
  FA_X1 U291 ( .A(n471), .B(n460), .CI(n833), .CO(n457), .S(n458) );
  FA_X1 U292 ( .A(n810), .B(n462), .CI(n473), .CO(n459), .S(n460) );
  FA_X1 U293 ( .A(n475), .B(n464), .CI(n787), .CO(n461), .S(n462) );
  FA_X1 U294 ( .A(n764), .B(n466), .CI(n477), .CO(n463), .S(n464) );
  FA_X1 U295 ( .A(n479), .B(n879), .CI(n741), .CO(n465), .S(n466) );
  FA_X1 U296 ( .A(n880), .B(n857), .CI(n470), .CO(n467), .S(n468) );
  FA_X1 U297 ( .A(n472), .B(n485), .CI(n483), .CO(n469), .S(n470) );
  FA_X1 U298 ( .A(n474), .B(n811), .CI(n834), .CO(n471), .S(n472) );
  FA_X1 U299 ( .A(n476), .B(n489), .CI(n487), .CO(n473), .S(n474) );
  FA_X1 U300 ( .A(n478), .B(n765), .CI(n788), .CO(n475), .S(n476) );
  FA_X1 U301 ( .A(n742), .B(n493), .CI(n491), .CO(n477), .S(n478) );
  FA_X1 U303 ( .A(n484), .B(n858), .CI(n881), .CO(n481), .S(n482) );
  FA_X1 U304 ( .A(n486), .B(n498), .CI(n496), .CO(n483), .S(n484) );
  FA_X1 U305 ( .A(n488), .B(n812), .CI(n835), .CO(n485), .S(n486) );
  FA_X1 U306 ( .A(n490), .B(n502), .CI(n500), .CO(n487), .S(n488) );
  FA_X1 U307 ( .A(n492), .B(n504), .CI(n789), .CO(n489), .S(n490) );
  FA_X1 U308 ( .A(n743), .B(n493), .CI(n766), .CO(n491), .S(n492) );
  FA_X1 U310 ( .A(n497), .B(n509), .CI(n882), .CO(n494), .S(n495) );
  FA_X1 U311 ( .A(n499), .B(n511), .CI(n859), .CO(n496), .S(n497) );
  FA_X1 U312 ( .A(n501), .B(n513), .CI(n836), .CO(n498), .S(n499) );
  FA_X1 U313 ( .A(n503), .B(n515), .CI(n813), .CO(n500), .S(n501) );
  FA_X1 U314 ( .A(n505), .B(n517), .CI(n790), .CO(n502), .S(n503) );
  FA_X1 U315 ( .A(n506), .B(n744), .CI(n767), .CO(n504), .S(n505) );
  FA_X1 U318 ( .A(n883), .B(n510), .CI(n521), .CO(n507), .S(n508) );
  FA_X1 U319 ( .A(n860), .B(n512), .CI(n523), .CO(n509), .S(n510) );
  FA_X1 U320 ( .A(n837), .B(n514), .CI(n525), .CO(n511), .S(n512) );
  FA_X1 U321 ( .A(n814), .B(n516), .CI(n527), .CO(n513), .S(n514) );
  FA_X1 U322 ( .A(n791), .B(n518), .CI(n529), .CO(n515), .S(n516) );
  FA_X1 U323 ( .A(n768), .B(n520), .CI(n531), .CO(n517), .S(n518) );
  HA_X1 U324 ( .A(n533), .B(n745), .CO(n519), .S(n520) );
  FA_X1 U325 ( .A(n884), .B(n524), .CI(n535), .CO(n521), .S(n522) );
  FA_X1 U326 ( .A(n861), .B(n526), .CI(n537), .CO(n523), .S(n524) );
  FA_X1 U327 ( .A(n838), .B(n528), .CI(n539), .CO(n525), .S(n526) );
  FA_X1 U328 ( .A(n815), .B(n530), .CI(n541), .CO(n527), .S(n528) );
  FA_X1 U329 ( .A(n792), .B(n532), .CI(n543), .CO(n529), .S(n530) );
  FA_X1 U330 ( .A(n769), .B(n534), .CI(n545), .CO(n531), .S(n532) );
  HA_X1 U331 ( .A(n547), .B(n746), .CO(n533), .S(n534) );
  FA_X1 U332 ( .A(n885), .B(n538), .CI(n549), .CO(n535), .S(n536) );
  FA_X1 U333 ( .A(n862), .B(n540), .CI(n551), .CO(n537), .S(n538) );
  FA_X1 U334 ( .A(n839), .B(n542), .CI(n553), .CO(n539), .S(n540) );
  FA_X1 U335 ( .A(n816), .B(n544), .CI(n555), .CO(n541), .S(n542) );
  FA_X1 U336 ( .A(n793), .B(n546), .CI(n557), .CO(n543), .S(n544) );
  FA_X1 U337 ( .A(n770), .B(n548), .CI(n559), .CO(n545), .S(n546) );
  HA_X1 U338 ( .A(n561), .B(n747), .CO(n547), .S(n548) );
  FA_X1 U339 ( .A(n886), .B(n552), .CI(n563), .CO(n549), .S(n550) );
  FA_X1 U340 ( .A(n863), .B(n554), .CI(n565), .CO(n551), .S(n552) );
  FA_X1 U341 ( .A(n840), .B(n556), .CI(n567), .CO(n553), .S(n554) );
  FA_X1 U342 ( .A(n817), .B(n558), .CI(n569), .CO(n555), .S(n556) );
  FA_X1 U343 ( .A(n794), .B(n560), .CI(n571), .CO(n557), .S(n558) );
  FA_X1 U344 ( .A(n771), .B(n562), .CI(n573), .CO(n559), .S(n560) );
  HA_X1 U345 ( .A(n748), .B(n1540), .CO(n561), .S(n562) );
  FA_X1 U346 ( .A(n887), .B(n566), .CI(n575), .CO(n563), .S(n564) );
  FA_X1 U347 ( .A(n864), .B(n568), .CI(n577), .CO(n565), .S(n566) );
  FA_X1 U348 ( .A(n841), .B(n570), .CI(n579), .CO(n567), .S(n568) );
  FA_X1 U349 ( .A(n818), .B(n572), .CI(n581), .CO(n569), .S(n570) );
  FA_X1 U350 ( .A(n795), .B(n574), .CI(n583), .CO(n571), .S(n572) );
  HA_X1 U351 ( .A(n585), .B(n772), .CO(n573), .S(n574) );
  FA_X1 U352 ( .A(n888), .B(n578), .CI(n587), .CO(n575), .S(n576) );
  FA_X1 U353 ( .A(n865), .B(n580), .CI(n589), .CO(n577), .S(n578) );
  FA_X1 U354 ( .A(n842), .B(n582), .CI(n591), .CO(n579), .S(n580) );
  FA_X1 U355 ( .A(n819), .B(n584), .CI(n593), .CO(n581), .S(n582) );
  FA_X1 U356 ( .A(n796), .B(n586), .CI(n595), .CO(n583), .S(n584) );
  HA_X1 U357 ( .A(n597), .B(n773), .CO(n585), .S(n586) );
  FA_X1 U358 ( .A(n889), .B(n590), .CI(n599), .CO(n587), .S(n588) );
  FA_X1 U359 ( .A(n866), .B(n592), .CI(n601), .CO(n589), .S(n590) );
  FA_X1 U360 ( .A(n843), .B(n594), .CI(n603), .CO(n591), .S(n592) );
  FA_X1 U361 ( .A(n820), .B(n596), .CI(n605), .CO(n593), .S(n594) );
  FA_X1 U362 ( .A(n797), .B(n598), .CI(n607), .CO(n595), .S(n596) );
  HA_X1 U363 ( .A(n774), .B(n1542), .CO(n597), .S(n598) );
  FA_X1 U364 ( .A(n890), .B(n602), .CI(n609), .CO(n599), .S(n600) );
  FA_X1 U365 ( .A(n867), .B(n604), .CI(n611), .CO(n601), .S(n602) );
  FA_X1 U366 ( .A(n844), .B(n606), .CI(n613), .CO(n603), .S(n604) );
  FA_X1 U367 ( .A(n821), .B(n608), .CI(n615), .CO(n605), .S(n606) );
  HA_X1 U368 ( .A(n617), .B(n798), .CO(n607), .S(n608) );
  FA_X1 U369 ( .A(n891), .B(n612), .CI(n619), .CO(n609), .S(n610) );
  FA_X1 U370 ( .A(n868), .B(n614), .CI(n621), .CO(n611), .S(n612) );
  FA_X1 U371 ( .A(n845), .B(n616), .CI(n623), .CO(n613), .S(n614) );
  FA_X1 U372 ( .A(n822), .B(n618), .CI(n625), .CO(n615), .S(n616) );
  HA_X1 U373 ( .A(n627), .B(n799), .CO(n617), .S(n618) );
  FA_X1 U374 ( .A(n892), .B(n622), .CI(n629), .CO(n619), .S(n620) );
  FA_X1 U375 ( .A(n869), .B(n624), .CI(n631), .CO(n621), .S(n622) );
  FA_X1 U376 ( .A(n846), .B(n626), .CI(n633), .CO(n623), .S(n624) );
  FA_X1 U377 ( .A(n823), .B(n628), .CI(n635), .CO(n625), .S(n626) );
  HA_X1 U378 ( .A(n800), .B(n1544), .CO(n627), .S(n628) );
  FA_X1 U379 ( .A(n893), .B(n632), .CI(n637), .CO(n629), .S(n630) );
  FA_X1 U380 ( .A(n870), .B(n634), .CI(n639), .CO(n631), .S(n632) );
  FA_X1 U381 ( .A(n847), .B(n636), .CI(n641), .CO(n633), .S(n634) );
  HA_X1 U382 ( .A(n643), .B(n824), .CO(n635), .S(n636) );
  FA_X1 U383 ( .A(n894), .B(n640), .CI(n645), .CO(n637), .S(n638) );
  FA_X1 U384 ( .A(n871), .B(n642), .CI(n647), .CO(n639), .S(n640) );
  FA_X1 U385 ( .A(n848), .B(n644), .CI(n649), .CO(n641), .S(n642) );
  HA_X1 U386 ( .A(n651), .B(n825), .CO(n643), .S(n644) );
  FA_X1 U387 ( .A(n895), .B(n648), .CI(n653), .CO(n645), .S(n646) );
  FA_X1 U388 ( .A(n872), .B(n650), .CI(n655), .CO(n647), .S(n648) );
  FA_X1 U389 ( .A(n849), .B(n652), .CI(n657), .CO(n649), .S(n650) );
  HA_X1 U390 ( .A(n826), .B(n1546), .CO(n651), .S(n652) );
  FA_X1 U391 ( .A(n896), .B(n656), .CI(n659), .CO(n653), .S(n654) );
  FA_X1 U392 ( .A(n873), .B(n658), .CI(n661), .CO(n655), .S(n656) );
  HA_X1 U393 ( .A(n663), .B(n850), .CO(n657), .S(n658) );
  FA_X1 U394 ( .A(n897), .B(n662), .CI(n665), .CO(n659), .S(n660) );
  FA_X1 U395 ( .A(n874), .B(n664), .CI(n667), .CO(n661), .S(n662) );
  HA_X1 U396 ( .A(n669), .B(n851), .CO(n663), .S(n664) );
  FA_X1 U397 ( .A(n898), .B(n668), .CI(n671), .CO(n665), .S(n666) );
  FA_X1 U398 ( .A(n875), .B(n670), .CI(n673), .CO(n667), .S(n668) );
  HA_X1 U399 ( .A(n852), .B(n1548), .CO(n669), .S(n670) );
  FA_X1 U400 ( .A(n899), .B(n674), .CI(n675), .CO(n671), .S(n672) );
  HA_X1 U401 ( .A(n677), .B(n876), .CO(n673), .S(n674) );
  FA_X1 U402 ( .A(n900), .B(n678), .CI(n679), .CO(n675), .S(n676) );
  HA_X1 U403 ( .A(n681), .B(n877), .CO(n677), .S(n678) );
  FA_X1 U404 ( .A(n901), .B(n682), .CI(n683), .CO(n679), .S(n680) );
  HA_X1 U405 ( .A(n878), .B(n1550), .CO(n681), .S(n682) );
  HA_X1 U406 ( .A(n685), .B(n902), .CO(n683), .S(n684) );
  HA_X1 U407 ( .A(n687), .B(n903), .CO(n685), .S(n686) );
  HA_X1 U408 ( .A(n904), .B(n1552), .CO(n687), .S(n688) );
  FA_X1 U1112 ( .A(B[22]), .B(n1554), .CI(n706), .CO(n1374), .S(n1375) );
  FA_X1 U1113 ( .A(B[21]), .B(B[22]), .CI(n707), .CO(n706), .S(n1376) );
  FA_X1 U1114 ( .A(B[20]), .B(B[21]), .CI(n708), .CO(n707), .S(n1377) );
  FA_X1 U1115 ( .A(B[19]), .B(B[20]), .CI(n709), .CO(n708), .S(n1378) );
  FA_X1 U1116 ( .A(B[18]), .B(B[19]), .CI(n710), .CO(n709), .S(n1379) );
  FA_X1 U1117 ( .A(B[17]), .B(B[18]), .CI(n711), .CO(n710), .S(n1380) );
  FA_X1 U1118 ( .A(B[16]), .B(B[17]), .CI(n712), .CO(n711), .S(n1381) );
  FA_X1 U1119 ( .A(B[15]), .B(B[16]), .CI(n713), .CO(n712), .S(n1382) );
  FA_X1 U1120 ( .A(B[14]), .B(B[15]), .CI(n714), .CO(n713), .S(n1383) );
  FA_X1 U1121 ( .A(B[13]), .B(B[14]), .CI(n715), .CO(n714), .S(n1384) );
  FA_X1 U1122 ( .A(B[12]), .B(B[13]), .CI(n716), .CO(n715), .S(n1385) );
  FA_X1 U1123 ( .A(B[11]), .B(B[12]), .CI(n717), .CO(n716), .S(n1386) );
  FA_X1 U1124 ( .A(B[10]), .B(B[11]), .CI(n718), .CO(n717), .S(n1387) );
  FA_X1 U1125 ( .A(B[9]), .B(B[10]), .CI(n719), .CO(n718), .S(n1388) );
  FA_X1 U1126 ( .A(B[8]), .B(B[9]), .CI(n720), .CO(n719), .S(n1389) );
  FA_X1 U1127 ( .A(B[7]), .B(B[8]), .CI(n721), .CO(n720), .S(n1390) );
  FA_X1 U1128 ( .A(B[6]), .B(B[7]), .CI(n722), .CO(n721), .S(n1391) );
  FA_X1 U1129 ( .A(B[5]), .B(B[6]), .CI(n723), .CO(n722), .S(n1392) );
  FA_X1 U1130 ( .A(B[4]), .B(B[5]), .CI(n724), .CO(n723), .S(n1393) );
  FA_X1 U1131 ( .A(B[3]), .B(B[4]), .CI(n725), .CO(n724), .S(n1394) );
  FA_X1 U1132 ( .A(B[2]), .B(B[3]), .CI(n726), .CO(n725), .S(n1395) );
  FA_X1 U1133 ( .A(B[1]), .B(B[2]), .CI(n727), .CO(n726), .S(n1396) );
  HA_X1 U1134 ( .A(B[0]), .B(B[1]), .CO(n727), .S(n1397) );
  OR2_X1 U1138 ( .A1(n2134), .A2(n2133), .ZN(n1534) );
  INV_X1 U1139 ( .A(n1534), .ZN(n1536) );
  INV_X1 U1140 ( .A(n1535), .ZN(n1537) );
  BUF_X1 U1141 ( .A(n1980), .Z(n1538) );
  BUF_X1 U1142 ( .A(n1980), .Z(n1539) );
  NAND3_X1 U1143 ( .A1(n1673), .A2(n1672), .A3(n1671), .ZN(n1586) );
  NAND3_X1 U1144 ( .A1(n1854), .A2(n1853), .A3(n1852), .ZN(n1804) );
  NAND3_X1 U1145 ( .A1(n1794), .A2(n1793), .A3(n1792), .ZN(n1744) );
  NAND3_X1 U1146 ( .A1(n1734), .A2(n1733), .A3(n1732), .ZN(n1684) );
  NAND3_X1 U1147 ( .A1(n2111), .A2(n2112), .A3(n2113), .ZN(n1563) );
  NAND2_X1 U1148 ( .A1(n1911), .A2(n1913), .ZN(n1857) );
  NAND2_X1 U1149 ( .A1(n1851), .A2(n1853), .ZN(n1797) );
  NAND2_X1 U1150 ( .A1(n1791), .A2(n1793), .ZN(n1737) );
  NAND2_X1 U1151 ( .A1(n1731), .A2(n1733), .ZN(n1677) );
  INV_X1 U1152 ( .A(n1553), .ZN(n1552) );
  INV_X1 U1153 ( .A(n1549), .ZN(n1548) );
  INV_X1 U1154 ( .A(n1551), .ZN(n1550) );
  NAND3_X1 U1155 ( .A1(n1914), .A2(n1913), .A3(n1912), .ZN(n1864) );
  NAND3_X1 U1156 ( .A1(n1974), .A2(n1973), .A3(n1972), .ZN(n1924) );
  NAND2_X1 U1157 ( .A1(n2134), .A2(n2132), .ZN(n1976) );
  NAND2_X1 U1158 ( .A1(n1971), .A2(n1973), .ZN(n1917) );
  INV_X1 U1159 ( .A(n1541), .ZN(n1540) );
  INV_X1 U1160 ( .A(n1543), .ZN(n1542) );
  INV_X1 U1161 ( .A(n1545), .ZN(n1544) );
  INV_X1 U1162 ( .A(n1547), .ZN(n1546) );
  INV_X1 U1163 ( .A(n1555), .ZN(n1554) );
  OR2_X1 U1164 ( .A1(n2132), .A2(n2131), .ZN(n1535) );
  NAND2_X1 U1165 ( .A1(A[0]), .A2(n2111), .ZN(n1561) );
  INV_X2 U1166 ( .A(B[0]), .ZN(n1574) );
  INV_X1 U1167 ( .A(A[5]), .ZN(n1553) );
  INV_X1 U1168 ( .A(A[11]), .ZN(n1549) );
  INV_X1 U1169 ( .A(A[8]), .ZN(n1551) );
  INV_X1 U1170 ( .A(A[17]), .ZN(n1545) );
  INV_X1 U1171 ( .A(A[14]), .ZN(n1547) );
  INV_X1 U1172 ( .A(A[23]), .ZN(n1541) );
  INV_X1 U1173 ( .A(A[20]), .ZN(n1543) );
  NOR2_X4 U1174 ( .A1(n1670), .A2(n1671), .ZN(n1581) );
  NOR2_X4 U1175 ( .A1(n1672), .A2(n1673), .ZN(n1582) );
  NAND2_X2 U1176 ( .A1(n1670), .A2(n1672), .ZN(n1576) );
  NOR2_X4 U1177 ( .A1(n1731), .A2(n1732), .ZN(n1680) );
  NOR2_X4 U1178 ( .A1(n1733), .A2(n1734), .ZN(n1681) );
  NOR2_X4 U1179 ( .A1(n1791), .A2(n1792), .ZN(n1740) );
  NOR2_X4 U1180 ( .A1(n1793), .A2(n1794), .ZN(n1741) );
  NOR2_X4 U1181 ( .A1(n1851), .A2(n1852), .ZN(n1800) );
  NOR2_X4 U1182 ( .A1(n1853), .A2(n1854), .ZN(n1801) );
  NOR2_X4 U1183 ( .A1(n1911), .A2(n1912), .ZN(n1860) );
  NOR2_X4 U1184 ( .A1(n1913), .A2(n1914), .ZN(n1861) );
  NOR2_X4 U1185 ( .A1(n1971), .A2(n1972), .ZN(n1920) );
  NOR2_X4 U1186 ( .A1(n1973), .A2(n1974), .ZN(n1921) );
  NOR2_X4 U1187 ( .A1(n2112), .A2(n2111), .ZN(n1558) );
  NOR2_X4 U1188 ( .A1(n2113), .A2(A[0]), .ZN(n1559) );
  INV_X1 U1189 ( .A(B[23]), .ZN(n1555) );
  INV_X1 U1190 ( .A(B[23]), .ZN(n1556) );
  XNOR2_X1 U1191 ( .A(A[2]), .B(n1557), .ZN(n908) );
  AOI221_X1 U1192 ( .B1(B[22]), .B2(n1558), .C1(B[21]), .C2(n1559), .A(n1560), 
        .ZN(n1557) );
  OAI22_X1 U1193 ( .A1(n1561), .A2(n1562), .B1(n1563), .B2(n1564), .ZN(n1560)
         );
  XNOR2_X1 U1194 ( .A(A[2]), .B(n1565), .ZN(n907) );
  AOI221_X1 U1195 ( .B1(B[23]), .B2(n1558), .C1(n1559), .C2(B[22]), .A(n1566), 
        .ZN(n1565) );
  OAI22_X1 U1196 ( .A1(n1561), .A2(n1567), .B1(n1568), .B2(n1563), .ZN(n1566)
         );
  XNOR2_X1 U1197 ( .A(A[2]), .B(n1569), .ZN(n906) );
  AOI221_X1 U1198 ( .B1(B[23]), .B2(n1558), .C1(n1554), .C2(n1559), .A(n1570), 
        .ZN(n1569) );
  OAI22_X1 U1199 ( .A1(n1561), .A2(n1571), .B1(n1572), .B2(n1563), .ZN(n1570)
         );
  XNOR2_X1 U1200 ( .A(n1573), .B(n1553), .ZN(n904) );
  OAI22_X1 U1201 ( .A1(n1574), .A2(n1575), .B1(n1576), .B2(n1574), .ZN(n1573)
         );
  XNOR2_X1 U1202 ( .A(n1577), .B(n1553), .ZN(n903) );
  OAI222_X1 U1203 ( .A1(n1575), .A2(n1578), .B1(n1574), .B2(n1579), .C1(n1576), 
        .C2(n1580), .ZN(n1577) );
  INV_X1 U1204 ( .A(n1581), .ZN(n1579) );
  INV_X1 U1205 ( .A(n1582), .ZN(n1575) );
  XNOR2_X1 U1206 ( .A(n1552), .B(n1583), .ZN(n902) );
  AOI221_X1 U1207 ( .B1(B[2]), .B2(n1582), .C1(B[1]), .C2(n1581), .A(n1584), 
        .ZN(n1583) );
  OAI22_X1 U1208 ( .A1(n1576), .A2(n1585), .B1(n1574), .B2(n1586), .ZN(n1584)
         );
  XNOR2_X1 U1209 ( .A(n1552), .B(n1587), .ZN(n901) );
  AOI221_X1 U1210 ( .B1(B[3]), .B2(n1582), .C1(B[2]), .C2(n1581), .A(n1588), 
        .ZN(n1587) );
  OAI22_X1 U1211 ( .A1(n1576), .A2(n1589), .B1(n1578), .B2(n1586), .ZN(n1588)
         );
  XNOR2_X1 U1212 ( .A(n1552), .B(n1590), .ZN(n900) );
  AOI221_X1 U1213 ( .B1(B[4]), .B2(n1582), .C1(B[3]), .C2(n1581), .A(n1591), 
        .ZN(n1590) );
  OAI22_X1 U1214 ( .A1(n1576), .A2(n1592), .B1(n1593), .B2(n1586), .ZN(n1591)
         );
  XNOR2_X1 U1215 ( .A(n1552), .B(n1594), .ZN(n899) );
  AOI221_X1 U1216 ( .B1(B[5]), .B2(n1582), .C1(B[4]), .C2(n1581), .A(n1595), 
        .ZN(n1594) );
  OAI22_X1 U1217 ( .A1(n1576), .A2(n1596), .B1(n1586), .B2(n1597), .ZN(n1595)
         );
  XNOR2_X1 U1218 ( .A(n1552), .B(n1598), .ZN(n898) );
  AOI221_X1 U1219 ( .B1(B[6]), .B2(n1582), .C1(B[5]), .C2(n1581), .A(n1599), 
        .ZN(n1598) );
  OAI22_X1 U1220 ( .A1(n1576), .A2(n1600), .B1(n1586), .B2(n1601), .ZN(n1599)
         );
  XNOR2_X1 U1221 ( .A(n1552), .B(n1602), .ZN(n897) );
  AOI221_X1 U1222 ( .B1(B[7]), .B2(n1582), .C1(B[6]), .C2(n1581), .A(n1603), 
        .ZN(n1602) );
  OAI22_X1 U1223 ( .A1(n1576), .A2(n1604), .B1(n1586), .B2(n1605), .ZN(n1603)
         );
  XNOR2_X1 U1224 ( .A(n1552), .B(n1606), .ZN(n896) );
  AOI221_X1 U1225 ( .B1(B[8]), .B2(n1582), .C1(B[7]), .C2(n1581), .A(n1607), 
        .ZN(n1606) );
  OAI22_X1 U1226 ( .A1(n1576), .A2(n1608), .B1(n1586), .B2(n1609), .ZN(n1607)
         );
  XNOR2_X1 U1227 ( .A(n1552), .B(n1610), .ZN(n895) );
  AOI221_X1 U1228 ( .B1(B[9]), .B2(n1582), .C1(B[8]), .C2(n1581), .A(n1611), 
        .ZN(n1610) );
  OAI22_X1 U1229 ( .A1(n1576), .A2(n1612), .B1(n1586), .B2(n1613), .ZN(n1611)
         );
  XNOR2_X1 U1230 ( .A(n1552), .B(n1614), .ZN(n894) );
  AOI221_X1 U1231 ( .B1(B[10]), .B2(n1582), .C1(B[9]), .C2(n1581), .A(n1615), 
        .ZN(n1614) );
  OAI22_X1 U1232 ( .A1(n1576), .A2(n1616), .B1(n1586), .B2(n1617), .ZN(n1615)
         );
  XNOR2_X1 U1233 ( .A(n1552), .B(n1618), .ZN(n893) );
  AOI221_X1 U1234 ( .B1(B[11]), .B2(n1582), .C1(B[10]), .C2(n1581), .A(n1619), 
        .ZN(n1618) );
  OAI22_X1 U1235 ( .A1(n1576), .A2(n1620), .B1(n1586), .B2(n1621), .ZN(n1619)
         );
  XNOR2_X1 U1236 ( .A(n1552), .B(n1622), .ZN(n892) );
  AOI221_X1 U1237 ( .B1(B[12]), .B2(n1582), .C1(B[11]), .C2(n1581), .A(n1623), 
        .ZN(n1622) );
  OAI22_X1 U1238 ( .A1(n1576), .A2(n1624), .B1(n1586), .B2(n1625), .ZN(n1623)
         );
  XNOR2_X1 U1239 ( .A(n1552), .B(n1626), .ZN(n891) );
  AOI221_X1 U1240 ( .B1(B[13]), .B2(n1582), .C1(B[12]), .C2(n1581), .A(n1627), 
        .ZN(n1626) );
  OAI22_X1 U1241 ( .A1(n1576), .A2(n1628), .B1(n1586), .B2(n1629), .ZN(n1627)
         );
  XNOR2_X1 U1242 ( .A(n1552), .B(n1630), .ZN(n890) );
  AOI221_X1 U1243 ( .B1(B[14]), .B2(n1582), .C1(B[13]), .C2(n1581), .A(n1631), 
        .ZN(n1630) );
  OAI22_X1 U1244 ( .A1(n1576), .A2(n1632), .B1(n1586), .B2(n1633), .ZN(n1631)
         );
  XNOR2_X1 U1245 ( .A(n1552), .B(n1634), .ZN(n889) );
  AOI221_X1 U1246 ( .B1(B[15]), .B2(n1582), .C1(B[14]), .C2(n1581), .A(n1635), 
        .ZN(n1634) );
  OAI22_X1 U1247 ( .A1(n1576), .A2(n1636), .B1(n1586), .B2(n1637), .ZN(n1635)
         );
  XNOR2_X1 U1248 ( .A(n1552), .B(n1638), .ZN(n888) );
  AOI221_X1 U1249 ( .B1(B[16]), .B2(n1582), .C1(B[15]), .C2(n1581), .A(n1639), 
        .ZN(n1638) );
  OAI22_X1 U1250 ( .A1(n1576), .A2(n1640), .B1(n1586), .B2(n1641), .ZN(n1639)
         );
  XNOR2_X1 U1251 ( .A(n1552), .B(n1642), .ZN(n887) );
  AOI221_X1 U1252 ( .B1(B[17]), .B2(n1582), .C1(B[16]), .C2(n1581), .A(n1643), 
        .ZN(n1642) );
  OAI22_X1 U1253 ( .A1(n1576), .A2(n1644), .B1(n1586), .B2(n1645), .ZN(n1643)
         );
  XNOR2_X1 U1254 ( .A(n1552), .B(n1646), .ZN(n886) );
  AOI221_X1 U1255 ( .B1(B[18]), .B2(n1582), .C1(B[17]), .C2(n1581), .A(n1647), 
        .ZN(n1646) );
  OAI22_X1 U1256 ( .A1(n1576), .A2(n1648), .B1(n1586), .B2(n1649), .ZN(n1647)
         );
  XNOR2_X1 U1257 ( .A(n1552), .B(n1650), .ZN(n885) );
  AOI221_X1 U1258 ( .B1(B[19]), .B2(n1582), .C1(B[18]), .C2(n1581), .A(n1651), 
        .ZN(n1650) );
  OAI22_X1 U1259 ( .A1(n1576), .A2(n1652), .B1(n1586), .B2(n1653), .ZN(n1651)
         );
  XNOR2_X1 U1260 ( .A(A[5]), .B(n1654), .ZN(n884) );
  AOI221_X1 U1261 ( .B1(n1582), .B2(B[20]), .C1(B[19]), .C2(n1581), .A(n1655), 
        .ZN(n1654) );
  OAI22_X1 U1262 ( .A1(n1576), .A2(n1656), .B1(n1586), .B2(n1657), .ZN(n1655)
         );
  XNOR2_X1 U1263 ( .A(A[5]), .B(n1658), .ZN(n883) );
  AOI221_X1 U1264 ( .B1(n1582), .B2(B[21]), .C1(n1581), .C2(B[20]), .A(n1659), 
        .ZN(n1658) );
  OAI22_X1 U1265 ( .A1(n1576), .A2(n1660), .B1(n1586), .B2(n1661), .ZN(n1659)
         );
  XNOR2_X1 U1266 ( .A(A[5]), .B(n1662), .ZN(n882) );
  AOI221_X1 U1267 ( .B1(n1582), .B2(B[22]), .C1(n1581), .C2(B[21]), .A(n1663), 
        .ZN(n1662) );
  OAI22_X1 U1268 ( .A1(n1562), .A2(n1576), .B1(n1564), .B2(n1586), .ZN(n1663)
         );
  XNOR2_X1 U1269 ( .A(A[5]), .B(n1664), .ZN(n881) );
  AOI221_X1 U1270 ( .B1(n1582), .B2(B[23]), .C1(n1581), .C2(B[22]), .A(n1665), 
        .ZN(n1664) );
  OAI22_X1 U1271 ( .A1(n1567), .A2(n1576), .B1(n1568), .B2(n1586), .ZN(n1665)
         );
  XNOR2_X1 U1272 ( .A(A[5]), .B(n1666), .ZN(n880) );
  AOI221_X1 U1273 ( .B1(n1582), .B2(B[23]), .C1(n1581), .C2(n1554), .A(n1667), 
        .ZN(n1666) );
  OAI22_X1 U1274 ( .A1(n1571), .A2(n1576), .B1(n1572), .B2(n1586), .ZN(n1667)
         );
  XNOR2_X1 U1275 ( .A(n1552), .B(n1668), .ZN(n879) );
  OAI221_X1 U1276 ( .B1(n1556), .B2(n1586), .C1(n1556), .C2(n1576), .A(n1669), 
        .ZN(n1668) );
  OAI21_X1 U1277 ( .B1(n1582), .B2(n1581), .A(n1554), .ZN(n1669) );
  INV_X1 U1278 ( .A(n1673), .ZN(n1670) );
  XNOR2_X1 U1279 ( .A(A[3]), .B(A[4]), .ZN(n1671) );
  XNOR2_X1 U1280 ( .A(A[4]), .B(n1553), .ZN(n1672) );
  XOR2_X1 U1281 ( .A(A[3]), .B(n1674), .Z(n1673) );
  XNOR2_X1 U1282 ( .A(n1675), .B(n1551), .ZN(n878) );
  OAI22_X1 U1283 ( .A1(n1574), .A2(n1676), .B1(n1574), .B2(n1677), .ZN(n1675)
         );
  XNOR2_X1 U1284 ( .A(n1678), .B(n1551), .ZN(n877) );
  OAI222_X1 U1285 ( .A1(n1578), .A2(n1676), .B1(n1574), .B2(n1679), .C1(n1580), 
        .C2(n1677), .ZN(n1678) );
  INV_X1 U1286 ( .A(n1680), .ZN(n1679) );
  INV_X1 U1287 ( .A(n1681), .ZN(n1676) );
  XNOR2_X1 U1288 ( .A(n1550), .B(n1682), .ZN(n876) );
  AOI221_X1 U1289 ( .B1(n1681), .B2(B[2]), .C1(n1680), .C2(B[1]), .A(n1683), 
        .ZN(n1682) );
  OAI22_X1 U1290 ( .A1(n1585), .A2(n1677), .B1(n1574), .B2(n1684), .ZN(n1683)
         );
  XNOR2_X1 U1291 ( .A(n1550), .B(n1685), .ZN(n875) );
  AOI221_X1 U1292 ( .B1(n1681), .B2(B[3]), .C1(n1680), .C2(B[2]), .A(n1686), 
        .ZN(n1685) );
  OAI22_X1 U1293 ( .A1(n1589), .A2(n1677), .B1(n1578), .B2(n1684), .ZN(n1686)
         );
  XNOR2_X1 U1294 ( .A(n1550), .B(n1687), .ZN(n874) );
  AOI221_X1 U1295 ( .B1(n1681), .B2(B[4]), .C1(n1680), .C2(B[3]), .A(n1688), 
        .ZN(n1687) );
  OAI22_X1 U1296 ( .A1(n1592), .A2(n1677), .B1(n1593), .B2(n1684), .ZN(n1688)
         );
  XNOR2_X1 U1297 ( .A(n1550), .B(n1689), .ZN(n873) );
  AOI221_X1 U1298 ( .B1(n1681), .B2(B[5]), .C1(n1680), .C2(B[4]), .A(n1690), 
        .ZN(n1689) );
  OAI22_X1 U1299 ( .A1(n1596), .A2(n1677), .B1(n1597), .B2(n1684), .ZN(n1690)
         );
  XNOR2_X1 U1300 ( .A(n1550), .B(n1691), .ZN(n872) );
  AOI221_X1 U1301 ( .B1(n1681), .B2(B[6]), .C1(n1680), .C2(B[5]), .A(n1692), 
        .ZN(n1691) );
  OAI22_X1 U1302 ( .A1(n1600), .A2(n1677), .B1(n1601), .B2(n1684), .ZN(n1692)
         );
  XNOR2_X1 U1303 ( .A(n1550), .B(n1693), .ZN(n871) );
  AOI221_X1 U1304 ( .B1(n1681), .B2(B[7]), .C1(n1680), .C2(B[6]), .A(n1694), 
        .ZN(n1693) );
  OAI22_X1 U1305 ( .A1(n1604), .A2(n1677), .B1(n1605), .B2(n1684), .ZN(n1694)
         );
  XNOR2_X1 U1306 ( .A(n1550), .B(n1695), .ZN(n870) );
  AOI221_X1 U1307 ( .B1(n1681), .B2(B[8]), .C1(n1680), .C2(B[7]), .A(n1696), 
        .ZN(n1695) );
  OAI22_X1 U1308 ( .A1(n1608), .A2(n1677), .B1(n1609), .B2(n1684), .ZN(n1696)
         );
  XNOR2_X1 U1309 ( .A(n1550), .B(n1697), .ZN(n869) );
  AOI221_X1 U1310 ( .B1(n1681), .B2(B[9]), .C1(n1680), .C2(B[8]), .A(n1698), 
        .ZN(n1697) );
  OAI22_X1 U1311 ( .A1(n1612), .A2(n1677), .B1(n1613), .B2(n1684), .ZN(n1698)
         );
  XNOR2_X1 U1312 ( .A(n1550), .B(n1699), .ZN(n868) );
  AOI221_X1 U1313 ( .B1(n1681), .B2(B[10]), .C1(n1680), .C2(B[9]), .A(n1700), 
        .ZN(n1699) );
  OAI22_X1 U1314 ( .A1(n1616), .A2(n1677), .B1(n1617), .B2(n1684), .ZN(n1700)
         );
  XNOR2_X1 U1315 ( .A(n1550), .B(n1701), .ZN(n867) );
  AOI221_X1 U1316 ( .B1(n1681), .B2(B[11]), .C1(n1680), .C2(B[10]), .A(n1702), 
        .ZN(n1701) );
  OAI22_X1 U1317 ( .A1(n1620), .A2(n1677), .B1(n1621), .B2(n1684), .ZN(n1702)
         );
  XNOR2_X1 U1318 ( .A(n1550), .B(n1703), .ZN(n866) );
  AOI221_X1 U1319 ( .B1(n1681), .B2(B[12]), .C1(n1680), .C2(B[11]), .A(n1704), 
        .ZN(n1703) );
  OAI22_X1 U1320 ( .A1(n1624), .A2(n1677), .B1(n1625), .B2(n1684), .ZN(n1704)
         );
  XNOR2_X1 U1321 ( .A(n1550), .B(n1705), .ZN(n865) );
  AOI221_X1 U1322 ( .B1(n1681), .B2(B[13]), .C1(n1680), .C2(B[12]), .A(n1706), 
        .ZN(n1705) );
  OAI22_X1 U1323 ( .A1(n1628), .A2(n1677), .B1(n1629), .B2(n1684), .ZN(n1706)
         );
  XNOR2_X1 U1324 ( .A(n1550), .B(n1707), .ZN(n864) );
  AOI221_X1 U1325 ( .B1(n1681), .B2(B[14]), .C1(n1680), .C2(B[13]), .A(n1708), 
        .ZN(n1707) );
  OAI22_X1 U1326 ( .A1(n1632), .A2(n1677), .B1(n1633), .B2(n1684), .ZN(n1708)
         );
  XNOR2_X1 U1327 ( .A(n1550), .B(n1709), .ZN(n863) );
  AOI221_X1 U1328 ( .B1(n1681), .B2(B[15]), .C1(n1680), .C2(B[14]), .A(n1710), 
        .ZN(n1709) );
  OAI22_X1 U1329 ( .A1(n1636), .A2(n1677), .B1(n1637), .B2(n1684), .ZN(n1710)
         );
  XNOR2_X1 U1330 ( .A(n1550), .B(n1711), .ZN(n862) );
  AOI221_X1 U1331 ( .B1(n1681), .B2(B[16]), .C1(n1680), .C2(B[15]), .A(n1712), 
        .ZN(n1711) );
  OAI22_X1 U1332 ( .A1(n1640), .A2(n1677), .B1(n1641), .B2(n1684), .ZN(n1712)
         );
  XNOR2_X1 U1333 ( .A(n1550), .B(n1713), .ZN(n861) );
  AOI221_X1 U1334 ( .B1(n1681), .B2(B[17]), .C1(n1680), .C2(B[16]), .A(n1714), 
        .ZN(n1713) );
  OAI22_X1 U1335 ( .A1(n1644), .A2(n1677), .B1(n1645), .B2(n1684), .ZN(n1714)
         );
  XNOR2_X1 U1336 ( .A(n1550), .B(n1715), .ZN(n860) );
  AOI221_X1 U1337 ( .B1(n1681), .B2(B[18]), .C1(n1680), .C2(B[17]), .A(n1716), 
        .ZN(n1715) );
  OAI22_X1 U1338 ( .A1(n1648), .A2(n1677), .B1(n1649), .B2(n1684), .ZN(n1716)
         );
  XNOR2_X1 U1339 ( .A(n1550), .B(n1717), .ZN(n859) );
  AOI221_X1 U1340 ( .B1(n1681), .B2(B[19]), .C1(n1680), .C2(B[18]), .A(n1718), 
        .ZN(n1717) );
  OAI22_X1 U1341 ( .A1(n1652), .A2(n1677), .B1(n1653), .B2(n1684), .ZN(n1718)
         );
  XNOR2_X1 U1342 ( .A(A[8]), .B(n1719), .ZN(n858) );
  AOI221_X1 U1343 ( .B1(n1681), .B2(B[20]), .C1(n1680), .C2(B[19]), .A(n1720), 
        .ZN(n1719) );
  OAI22_X1 U1344 ( .A1(n1656), .A2(n1677), .B1(n1657), .B2(n1684), .ZN(n1720)
         );
  XNOR2_X1 U1345 ( .A(A[8]), .B(n1721), .ZN(n857) );
  AOI221_X1 U1346 ( .B1(n1681), .B2(B[21]), .C1(n1680), .C2(B[20]), .A(n1722), 
        .ZN(n1721) );
  OAI22_X1 U1347 ( .A1(n1660), .A2(n1677), .B1(n1661), .B2(n1684), .ZN(n1722)
         );
  XNOR2_X1 U1348 ( .A(A[8]), .B(n1723), .ZN(n856) );
  AOI221_X1 U1349 ( .B1(n1681), .B2(B[22]), .C1(n1680), .C2(B[21]), .A(n1724), 
        .ZN(n1723) );
  OAI22_X1 U1350 ( .A1(n1562), .A2(n1677), .B1(n1564), .B2(n1684), .ZN(n1724)
         );
  XNOR2_X1 U1351 ( .A(A[8]), .B(n1725), .ZN(n855) );
  AOI221_X1 U1352 ( .B1(n1681), .B2(B[23]), .C1(n1680), .C2(B[22]), .A(n1726), 
        .ZN(n1725) );
  OAI22_X1 U1353 ( .A1(n1567), .A2(n1677), .B1(n1568), .B2(n1684), .ZN(n1726)
         );
  XNOR2_X1 U1354 ( .A(A[8]), .B(n1727), .ZN(n854) );
  AOI221_X1 U1355 ( .B1(n1681), .B2(B[23]), .C1(n1680), .C2(n1554), .A(n1728), 
        .ZN(n1727) );
  OAI22_X1 U1356 ( .A1(n1571), .A2(n1677), .B1(n1572), .B2(n1684), .ZN(n1728)
         );
  XNOR2_X1 U1357 ( .A(n1550), .B(n1729), .ZN(n853) );
  OAI221_X1 U1358 ( .B1(n1555), .B2(n1684), .C1(n1556), .C2(n1677), .A(n1730), 
        .ZN(n1729) );
  OAI21_X1 U1359 ( .B1(n1681), .B2(n1680), .A(n1554), .ZN(n1730) );
  INV_X1 U1360 ( .A(n1734), .ZN(n1731) );
  XNOR2_X1 U1361 ( .A(A[6]), .B(A[7]), .ZN(n1732) );
  XNOR2_X1 U1362 ( .A(A[7]), .B(n1551), .ZN(n1733) );
  XOR2_X1 U1363 ( .A(A[6]), .B(n1553), .Z(n1734) );
  XNOR2_X1 U1364 ( .A(n1735), .B(n1549), .ZN(n852) );
  OAI22_X1 U1365 ( .A1(n1574), .A2(n1736), .B1(n1574), .B2(n1737), .ZN(n1735)
         );
  XNOR2_X1 U1366 ( .A(n1738), .B(n1549), .ZN(n851) );
  OAI222_X1 U1367 ( .A1(n1578), .A2(n1736), .B1(n1574), .B2(n1739), .C1(n1580), 
        .C2(n1737), .ZN(n1738) );
  INV_X1 U1368 ( .A(n1740), .ZN(n1739) );
  INV_X1 U1369 ( .A(n1741), .ZN(n1736) );
  XNOR2_X1 U1370 ( .A(n1548), .B(n1742), .ZN(n850) );
  AOI221_X1 U1371 ( .B1(n1741), .B2(B[2]), .C1(n1740), .C2(B[1]), .A(n1743), 
        .ZN(n1742) );
  OAI22_X1 U1372 ( .A1(n1585), .A2(n1737), .B1(n1574), .B2(n1744), .ZN(n1743)
         );
  XNOR2_X1 U1373 ( .A(n1548), .B(n1745), .ZN(n849) );
  AOI221_X1 U1374 ( .B1(n1741), .B2(B[3]), .C1(n1740), .C2(B[2]), .A(n1746), 
        .ZN(n1745) );
  OAI22_X1 U1375 ( .A1(n1589), .A2(n1737), .B1(n1578), .B2(n1744), .ZN(n1746)
         );
  XNOR2_X1 U1376 ( .A(n1548), .B(n1747), .ZN(n848) );
  AOI221_X1 U1377 ( .B1(n1741), .B2(B[4]), .C1(n1740), .C2(B[3]), .A(n1748), 
        .ZN(n1747) );
  OAI22_X1 U1378 ( .A1(n1592), .A2(n1737), .B1(n1593), .B2(n1744), .ZN(n1748)
         );
  XNOR2_X1 U1379 ( .A(n1548), .B(n1749), .ZN(n847) );
  AOI221_X1 U1380 ( .B1(n1741), .B2(B[5]), .C1(n1740), .C2(B[4]), .A(n1750), 
        .ZN(n1749) );
  OAI22_X1 U1381 ( .A1(n1596), .A2(n1737), .B1(n1597), .B2(n1744), .ZN(n1750)
         );
  XNOR2_X1 U1382 ( .A(n1548), .B(n1751), .ZN(n846) );
  AOI221_X1 U1383 ( .B1(n1741), .B2(B[6]), .C1(n1740), .C2(B[5]), .A(n1752), 
        .ZN(n1751) );
  OAI22_X1 U1384 ( .A1(n1600), .A2(n1737), .B1(n1601), .B2(n1744), .ZN(n1752)
         );
  XNOR2_X1 U1385 ( .A(n1548), .B(n1753), .ZN(n845) );
  AOI221_X1 U1386 ( .B1(n1741), .B2(B[7]), .C1(n1740), .C2(B[6]), .A(n1754), 
        .ZN(n1753) );
  OAI22_X1 U1387 ( .A1(n1604), .A2(n1737), .B1(n1605), .B2(n1744), .ZN(n1754)
         );
  XNOR2_X1 U1388 ( .A(n1548), .B(n1755), .ZN(n844) );
  AOI221_X1 U1389 ( .B1(n1741), .B2(B[8]), .C1(n1740), .C2(B[7]), .A(n1756), 
        .ZN(n1755) );
  OAI22_X1 U1390 ( .A1(n1608), .A2(n1737), .B1(n1609), .B2(n1744), .ZN(n1756)
         );
  XNOR2_X1 U1391 ( .A(n1548), .B(n1757), .ZN(n843) );
  AOI221_X1 U1392 ( .B1(n1741), .B2(B[9]), .C1(n1740), .C2(B[8]), .A(n1758), 
        .ZN(n1757) );
  OAI22_X1 U1393 ( .A1(n1612), .A2(n1737), .B1(n1613), .B2(n1744), .ZN(n1758)
         );
  XNOR2_X1 U1394 ( .A(n1548), .B(n1759), .ZN(n842) );
  AOI221_X1 U1395 ( .B1(n1741), .B2(B[10]), .C1(n1740), .C2(B[9]), .A(n1760), 
        .ZN(n1759) );
  OAI22_X1 U1396 ( .A1(n1616), .A2(n1737), .B1(n1617), .B2(n1744), .ZN(n1760)
         );
  XNOR2_X1 U1397 ( .A(n1548), .B(n1761), .ZN(n841) );
  AOI221_X1 U1398 ( .B1(n1741), .B2(B[11]), .C1(n1740), .C2(B[10]), .A(n1762), 
        .ZN(n1761) );
  OAI22_X1 U1399 ( .A1(n1620), .A2(n1737), .B1(n1621), .B2(n1744), .ZN(n1762)
         );
  XNOR2_X1 U1400 ( .A(n1548), .B(n1763), .ZN(n840) );
  AOI221_X1 U1401 ( .B1(n1741), .B2(B[12]), .C1(n1740), .C2(B[11]), .A(n1764), 
        .ZN(n1763) );
  OAI22_X1 U1402 ( .A1(n1624), .A2(n1737), .B1(n1625), .B2(n1744), .ZN(n1764)
         );
  XNOR2_X1 U1403 ( .A(n1548), .B(n1765), .ZN(n839) );
  AOI221_X1 U1404 ( .B1(n1741), .B2(B[13]), .C1(n1740), .C2(B[12]), .A(n1766), 
        .ZN(n1765) );
  OAI22_X1 U1405 ( .A1(n1628), .A2(n1737), .B1(n1629), .B2(n1744), .ZN(n1766)
         );
  XNOR2_X1 U1406 ( .A(n1548), .B(n1767), .ZN(n838) );
  AOI221_X1 U1407 ( .B1(n1741), .B2(B[14]), .C1(n1740), .C2(B[13]), .A(n1768), 
        .ZN(n1767) );
  OAI22_X1 U1408 ( .A1(n1632), .A2(n1737), .B1(n1633), .B2(n1744), .ZN(n1768)
         );
  XNOR2_X1 U1409 ( .A(n1548), .B(n1769), .ZN(n837) );
  AOI221_X1 U1410 ( .B1(n1741), .B2(B[15]), .C1(n1740), .C2(B[14]), .A(n1770), 
        .ZN(n1769) );
  OAI22_X1 U1411 ( .A1(n1636), .A2(n1737), .B1(n1637), .B2(n1744), .ZN(n1770)
         );
  XNOR2_X1 U1412 ( .A(n1548), .B(n1771), .ZN(n836) );
  AOI221_X1 U1413 ( .B1(n1741), .B2(B[16]), .C1(n1740), .C2(B[15]), .A(n1772), 
        .ZN(n1771) );
  OAI22_X1 U1414 ( .A1(n1640), .A2(n1737), .B1(n1641), .B2(n1744), .ZN(n1772)
         );
  XNOR2_X1 U1415 ( .A(n1548), .B(n1773), .ZN(n835) );
  AOI221_X1 U1416 ( .B1(n1741), .B2(B[17]), .C1(n1740), .C2(B[16]), .A(n1774), 
        .ZN(n1773) );
  OAI22_X1 U1417 ( .A1(n1644), .A2(n1737), .B1(n1645), .B2(n1744), .ZN(n1774)
         );
  XNOR2_X1 U1418 ( .A(n1548), .B(n1775), .ZN(n834) );
  AOI221_X1 U1419 ( .B1(n1741), .B2(B[18]), .C1(n1740), .C2(B[17]), .A(n1776), 
        .ZN(n1775) );
  OAI22_X1 U1420 ( .A1(n1648), .A2(n1737), .B1(n1649), .B2(n1744), .ZN(n1776)
         );
  XNOR2_X1 U1421 ( .A(n1548), .B(n1777), .ZN(n833) );
  AOI221_X1 U1422 ( .B1(n1741), .B2(B[19]), .C1(n1740), .C2(B[18]), .A(n1778), 
        .ZN(n1777) );
  OAI22_X1 U1423 ( .A1(n1652), .A2(n1737), .B1(n1653), .B2(n1744), .ZN(n1778)
         );
  XNOR2_X1 U1424 ( .A(n1548), .B(n1779), .ZN(n832) );
  AOI221_X1 U1425 ( .B1(n1741), .B2(B[20]), .C1(n1740), .C2(B[19]), .A(n1780), 
        .ZN(n1779) );
  OAI22_X1 U1426 ( .A1(n1656), .A2(n1737), .B1(n1657), .B2(n1744), .ZN(n1780)
         );
  XNOR2_X1 U1427 ( .A(A[11]), .B(n1781), .ZN(n831) );
  AOI221_X1 U1428 ( .B1(n1741), .B2(B[21]), .C1(n1740), .C2(B[20]), .A(n1782), 
        .ZN(n1781) );
  OAI22_X1 U1429 ( .A1(n1660), .A2(n1737), .B1(n1661), .B2(n1744), .ZN(n1782)
         );
  XNOR2_X1 U1430 ( .A(A[11]), .B(n1783), .ZN(n830) );
  AOI221_X1 U1431 ( .B1(n1741), .B2(B[22]), .C1(n1740), .C2(B[21]), .A(n1784), 
        .ZN(n1783) );
  OAI22_X1 U1432 ( .A1(n1562), .A2(n1737), .B1(n1564), .B2(n1744), .ZN(n1784)
         );
  XNOR2_X1 U1433 ( .A(A[11]), .B(n1785), .ZN(n829) );
  AOI221_X1 U1434 ( .B1(n1741), .B2(B[23]), .C1(n1740), .C2(B[22]), .A(n1786), 
        .ZN(n1785) );
  OAI22_X1 U1435 ( .A1(n1567), .A2(n1737), .B1(n1568), .B2(n1744), .ZN(n1786)
         );
  XNOR2_X1 U1436 ( .A(A[11]), .B(n1787), .ZN(n828) );
  AOI221_X1 U1437 ( .B1(n1741), .B2(B[23]), .C1(n1740), .C2(n1554), .A(n1788), 
        .ZN(n1787) );
  OAI22_X1 U1438 ( .A1(n1571), .A2(n1737), .B1(n1572), .B2(n1744), .ZN(n1788)
         );
  XNOR2_X1 U1439 ( .A(A[11]), .B(n1789), .ZN(n827) );
  OAI221_X1 U1440 ( .B1(n1556), .B2(n1744), .C1(n1556), .C2(n1737), .A(n1790), 
        .ZN(n1789) );
  OAI21_X1 U1441 ( .B1(n1741), .B2(n1740), .A(n1554), .ZN(n1790) );
  INV_X1 U1442 ( .A(n1794), .ZN(n1791) );
  XNOR2_X1 U1443 ( .A(A[10]), .B(A[9]), .ZN(n1792) );
  XNOR2_X1 U1444 ( .A(A[10]), .B(n1549), .ZN(n1793) );
  XOR2_X1 U1445 ( .A(A[9]), .B(n1551), .Z(n1794) );
  XNOR2_X1 U1446 ( .A(n1795), .B(n1547), .ZN(n826) );
  OAI22_X1 U1447 ( .A1(n1574), .A2(n1796), .B1(n1574), .B2(n1797), .ZN(n1795)
         );
  XNOR2_X1 U1448 ( .A(n1798), .B(n1547), .ZN(n825) );
  OAI222_X1 U1449 ( .A1(n1578), .A2(n1796), .B1(n1574), .B2(n1799), .C1(n1580), 
        .C2(n1797), .ZN(n1798) );
  INV_X1 U1450 ( .A(n1800), .ZN(n1799) );
  INV_X1 U1451 ( .A(n1801), .ZN(n1796) );
  XNOR2_X1 U1452 ( .A(n1546), .B(n1802), .ZN(n824) );
  AOI221_X1 U1453 ( .B1(n1801), .B2(B[2]), .C1(n1800), .C2(B[1]), .A(n1803), 
        .ZN(n1802) );
  OAI22_X1 U1454 ( .A1(n1585), .A2(n1797), .B1(n1574), .B2(n1804), .ZN(n1803)
         );
  XNOR2_X1 U1455 ( .A(n1546), .B(n1805), .ZN(n823) );
  AOI221_X1 U1456 ( .B1(n1801), .B2(B[3]), .C1(n1800), .C2(B[2]), .A(n1806), 
        .ZN(n1805) );
  OAI22_X1 U1457 ( .A1(n1589), .A2(n1797), .B1(n1578), .B2(n1804), .ZN(n1806)
         );
  XNOR2_X1 U1458 ( .A(n1546), .B(n1807), .ZN(n822) );
  AOI221_X1 U1459 ( .B1(n1801), .B2(B[4]), .C1(n1800), .C2(B[3]), .A(n1808), 
        .ZN(n1807) );
  OAI22_X1 U1460 ( .A1(n1592), .A2(n1797), .B1(n1593), .B2(n1804), .ZN(n1808)
         );
  XNOR2_X1 U1461 ( .A(n1546), .B(n1809), .ZN(n821) );
  AOI221_X1 U1462 ( .B1(n1801), .B2(B[5]), .C1(n1800), .C2(B[4]), .A(n1810), 
        .ZN(n1809) );
  OAI22_X1 U1463 ( .A1(n1596), .A2(n1797), .B1(n1597), .B2(n1804), .ZN(n1810)
         );
  XNOR2_X1 U1464 ( .A(n1546), .B(n1811), .ZN(n820) );
  AOI221_X1 U1465 ( .B1(n1801), .B2(B[6]), .C1(n1800), .C2(B[5]), .A(n1812), 
        .ZN(n1811) );
  OAI22_X1 U1466 ( .A1(n1600), .A2(n1797), .B1(n1601), .B2(n1804), .ZN(n1812)
         );
  XNOR2_X1 U1467 ( .A(n1546), .B(n1813), .ZN(n819) );
  AOI221_X1 U1468 ( .B1(n1801), .B2(B[7]), .C1(n1800), .C2(B[6]), .A(n1814), 
        .ZN(n1813) );
  OAI22_X1 U1469 ( .A1(n1604), .A2(n1797), .B1(n1605), .B2(n1804), .ZN(n1814)
         );
  XNOR2_X1 U1470 ( .A(n1546), .B(n1815), .ZN(n818) );
  AOI221_X1 U1471 ( .B1(n1801), .B2(B[8]), .C1(n1800), .C2(B[7]), .A(n1816), 
        .ZN(n1815) );
  OAI22_X1 U1472 ( .A1(n1608), .A2(n1797), .B1(n1609), .B2(n1804), .ZN(n1816)
         );
  XNOR2_X1 U1473 ( .A(n1546), .B(n1817), .ZN(n817) );
  AOI221_X1 U1474 ( .B1(n1801), .B2(B[9]), .C1(n1800), .C2(B[8]), .A(n1818), 
        .ZN(n1817) );
  OAI22_X1 U1475 ( .A1(n1612), .A2(n1797), .B1(n1613), .B2(n1804), .ZN(n1818)
         );
  XNOR2_X1 U1476 ( .A(n1546), .B(n1819), .ZN(n816) );
  AOI221_X1 U1477 ( .B1(n1801), .B2(B[10]), .C1(n1800), .C2(B[9]), .A(n1820), 
        .ZN(n1819) );
  OAI22_X1 U1478 ( .A1(n1616), .A2(n1797), .B1(n1617), .B2(n1804), .ZN(n1820)
         );
  XNOR2_X1 U1479 ( .A(n1546), .B(n1821), .ZN(n815) );
  AOI221_X1 U1480 ( .B1(n1801), .B2(B[11]), .C1(n1800), .C2(B[10]), .A(n1822), 
        .ZN(n1821) );
  OAI22_X1 U1481 ( .A1(n1620), .A2(n1797), .B1(n1621), .B2(n1804), .ZN(n1822)
         );
  XNOR2_X1 U1482 ( .A(n1546), .B(n1823), .ZN(n814) );
  AOI221_X1 U1483 ( .B1(n1801), .B2(B[12]), .C1(n1800), .C2(B[11]), .A(n1824), 
        .ZN(n1823) );
  OAI22_X1 U1484 ( .A1(n1624), .A2(n1797), .B1(n1625), .B2(n1804), .ZN(n1824)
         );
  XNOR2_X1 U1485 ( .A(n1546), .B(n1825), .ZN(n813) );
  AOI221_X1 U1486 ( .B1(n1801), .B2(B[13]), .C1(n1800), .C2(B[12]), .A(n1826), 
        .ZN(n1825) );
  OAI22_X1 U1487 ( .A1(n1628), .A2(n1797), .B1(n1629), .B2(n1804), .ZN(n1826)
         );
  XNOR2_X1 U1488 ( .A(n1546), .B(n1827), .ZN(n812) );
  AOI221_X1 U1489 ( .B1(n1801), .B2(B[14]), .C1(n1800), .C2(B[13]), .A(n1828), 
        .ZN(n1827) );
  OAI22_X1 U1490 ( .A1(n1632), .A2(n1797), .B1(n1633), .B2(n1804), .ZN(n1828)
         );
  XNOR2_X1 U1491 ( .A(n1546), .B(n1829), .ZN(n811) );
  AOI221_X1 U1492 ( .B1(n1801), .B2(B[15]), .C1(n1800), .C2(B[14]), .A(n1830), 
        .ZN(n1829) );
  OAI22_X1 U1493 ( .A1(n1636), .A2(n1797), .B1(n1637), .B2(n1804), .ZN(n1830)
         );
  XNOR2_X1 U1494 ( .A(n1546), .B(n1831), .ZN(n810) );
  AOI221_X1 U1495 ( .B1(n1801), .B2(B[16]), .C1(n1800), .C2(B[15]), .A(n1832), 
        .ZN(n1831) );
  OAI22_X1 U1496 ( .A1(n1640), .A2(n1797), .B1(n1641), .B2(n1804), .ZN(n1832)
         );
  XNOR2_X1 U1497 ( .A(n1546), .B(n1833), .ZN(n809) );
  AOI221_X1 U1498 ( .B1(n1801), .B2(B[17]), .C1(n1800), .C2(B[16]), .A(n1834), 
        .ZN(n1833) );
  OAI22_X1 U1499 ( .A1(n1644), .A2(n1797), .B1(n1645), .B2(n1804), .ZN(n1834)
         );
  XNOR2_X1 U1500 ( .A(n1546), .B(n1835), .ZN(n808) );
  AOI221_X1 U1501 ( .B1(n1801), .B2(B[18]), .C1(n1800), .C2(B[17]), .A(n1836), 
        .ZN(n1835) );
  OAI22_X1 U1502 ( .A1(n1648), .A2(n1797), .B1(n1649), .B2(n1804), .ZN(n1836)
         );
  XNOR2_X1 U1503 ( .A(n1546), .B(n1837), .ZN(n807) );
  AOI221_X1 U1504 ( .B1(n1801), .B2(B[19]), .C1(n1800), .C2(B[18]), .A(n1838), 
        .ZN(n1837) );
  OAI22_X1 U1505 ( .A1(n1652), .A2(n1797), .B1(n1653), .B2(n1804), .ZN(n1838)
         );
  XNOR2_X1 U1506 ( .A(n1546), .B(n1839), .ZN(n806) );
  AOI221_X1 U1507 ( .B1(n1801), .B2(B[20]), .C1(n1800), .C2(B[19]), .A(n1840), 
        .ZN(n1839) );
  OAI22_X1 U1508 ( .A1(n1656), .A2(n1797), .B1(n1657), .B2(n1804), .ZN(n1840)
         );
  XNOR2_X1 U1509 ( .A(A[14]), .B(n1841), .ZN(n805) );
  AOI221_X1 U1510 ( .B1(n1801), .B2(B[21]), .C1(n1800), .C2(B[20]), .A(n1842), 
        .ZN(n1841) );
  OAI22_X1 U1511 ( .A1(n1660), .A2(n1797), .B1(n1661), .B2(n1804), .ZN(n1842)
         );
  XNOR2_X1 U1512 ( .A(A[14]), .B(n1843), .ZN(n804) );
  AOI221_X1 U1513 ( .B1(n1801), .B2(B[22]), .C1(n1800), .C2(B[21]), .A(n1844), 
        .ZN(n1843) );
  OAI22_X1 U1514 ( .A1(n1562), .A2(n1797), .B1(n1564), .B2(n1804), .ZN(n1844)
         );
  XNOR2_X1 U1515 ( .A(A[14]), .B(n1845), .ZN(n803) );
  AOI221_X1 U1516 ( .B1(n1801), .B2(B[23]), .C1(n1800), .C2(B[22]), .A(n1846), 
        .ZN(n1845) );
  OAI22_X1 U1517 ( .A1(n1567), .A2(n1797), .B1(n1568), .B2(n1804), .ZN(n1846)
         );
  XNOR2_X1 U1518 ( .A(A[14]), .B(n1847), .ZN(n802) );
  AOI221_X1 U1519 ( .B1(n1801), .B2(B[23]), .C1(n1800), .C2(n1554), .A(n1848), 
        .ZN(n1847) );
  OAI22_X1 U1520 ( .A1(n1571), .A2(n1797), .B1(n1572), .B2(n1804), .ZN(n1848)
         );
  XNOR2_X1 U1521 ( .A(A[14]), .B(n1849), .ZN(n801) );
  OAI221_X1 U1522 ( .B1(n1556), .B2(n1804), .C1(n1556), .C2(n1797), .A(n1850), 
        .ZN(n1849) );
  OAI21_X1 U1523 ( .B1(n1801), .B2(n1800), .A(n1554), .ZN(n1850) );
  INV_X1 U1524 ( .A(n1854), .ZN(n1851) );
  XNOR2_X1 U1525 ( .A(A[12]), .B(A[13]), .ZN(n1852) );
  XNOR2_X1 U1526 ( .A(A[13]), .B(n1547), .ZN(n1853) );
  XOR2_X1 U1527 ( .A(A[12]), .B(n1549), .Z(n1854) );
  XNOR2_X1 U1528 ( .A(n1855), .B(n1545), .ZN(n800) );
  OAI22_X1 U1529 ( .A1(n1574), .A2(n1856), .B1(n1574), .B2(n1857), .ZN(n1855)
         );
  XNOR2_X1 U1530 ( .A(n1858), .B(n1545), .ZN(n799) );
  OAI222_X1 U1531 ( .A1(n1578), .A2(n1856), .B1(n1574), .B2(n1859), .C1(n1580), 
        .C2(n1857), .ZN(n1858) );
  INV_X1 U1532 ( .A(n1860), .ZN(n1859) );
  INV_X1 U1533 ( .A(n1861), .ZN(n1856) );
  XNOR2_X1 U1534 ( .A(n1544), .B(n1862), .ZN(n798) );
  AOI221_X1 U1535 ( .B1(n1861), .B2(B[2]), .C1(n1860), .C2(B[1]), .A(n1863), 
        .ZN(n1862) );
  OAI22_X1 U1536 ( .A1(n1585), .A2(n1857), .B1(n1574), .B2(n1864), .ZN(n1863)
         );
  XNOR2_X1 U1537 ( .A(n1544), .B(n1865), .ZN(n797) );
  AOI221_X1 U1538 ( .B1(n1861), .B2(B[3]), .C1(n1860), .C2(B[2]), .A(n1866), 
        .ZN(n1865) );
  OAI22_X1 U1539 ( .A1(n1589), .A2(n1857), .B1(n1578), .B2(n1864), .ZN(n1866)
         );
  XNOR2_X1 U1540 ( .A(n1544), .B(n1867), .ZN(n796) );
  AOI221_X1 U1541 ( .B1(n1861), .B2(B[4]), .C1(n1860), .C2(B[3]), .A(n1868), 
        .ZN(n1867) );
  OAI22_X1 U1542 ( .A1(n1592), .A2(n1857), .B1(n1593), .B2(n1864), .ZN(n1868)
         );
  XNOR2_X1 U1543 ( .A(n1544), .B(n1869), .ZN(n795) );
  AOI221_X1 U1544 ( .B1(n1861), .B2(B[5]), .C1(n1860), .C2(B[4]), .A(n1870), 
        .ZN(n1869) );
  OAI22_X1 U1545 ( .A1(n1596), .A2(n1857), .B1(n1597), .B2(n1864), .ZN(n1870)
         );
  XNOR2_X1 U1546 ( .A(n1544), .B(n1871), .ZN(n794) );
  AOI221_X1 U1547 ( .B1(n1861), .B2(B[6]), .C1(n1860), .C2(B[5]), .A(n1872), 
        .ZN(n1871) );
  OAI22_X1 U1548 ( .A1(n1600), .A2(n1857), .B1(n1601), .B2(n1864), .ZN(n1872)
         );
  XNOR2_X1 U1549 ( .A(n1544), .B(n1873), .ZN(n793) );
  AOI221_X1 U1550 ( .B1(n1861), .B2(B[7]), .C1(n1860), .C2(B[6]), .A(n1874), 
        .ZN(n1873) );
  OAI22_X1 U1551 ( .A1(n1604), .A2(n1857), .B1(n1605), .B2(n1864), .ZN(n1874)
         );
  XNOR2_X1 U1552 ( .A(n1544), .B(n1875), .ZN(n792) );
  AOI221_X1 U1553 ( .B1(n1861), .B2(B[8]), .C1(n1860), .C2(B[7]), .A(n1876), 
        .ZN(n1875) );
  OAI22_X1 U1554 ( .A1(n1608), .A2(n1857), .B1(n1609), .B2(n1864), .ZN(n1876)
         );
  XNOR2_X1 U1555 ( .A(n1544), .B(n1877), .ZN(n791) );
  AOI221_X1 U1556 ( .B1(n1861), .B2(B[9]), .C1(n1860), .C2(B[8]), .A(n1878), 
        .ZN(n1877) );
  OAI22_X1 U1557 ( .A1(n1612), .A2(n1857), .B1(n1613), .B2(n1864), .ZN(n1878)
         );
  XNOR2_X1 U1558 ( .A(n1544), .B(n1879), .ZN(n790) );
  AOI221_X1 U1559 ( .B1(n1861), .B2(B[10]), .C1(n1860), .C2(B[9]), .A(n1880), 
        .ZN(n1879) );
  OAI22_X1 U1560 ( .A1(n1616), .A2(n1857), .B1(n1617), .B2(n1864), .ZN(n1880)
         );
  XNOR2_X1 U1561 ( .A(n1544), .B(n1881), .ZN(n789) );
  AOI221_X1 U1562 ( .B1(n1861), .B2(B[11]), .C1(n1860), .C2(B[10]), .A(n1882), 
        .ZN(n1881) );
  OAI22_X1 U1563 ( .A1(n1620), .A2(n1857), .B1(n1621), .B2(n1864), .ZN(n1882)
         );
  XNOR2_X1 U1564 ( .A(n1544), .B(n1883), .ZN(n788) );
  AOI221_X1 U1565 ( .B1(n1861), .B2(B[12]), .C1(n1860), .C2(B[11]), .A(n1884), 
        .ZN(n1883) );
  OAI22_X1 U1566 ( .A1(n1624), .A2(n1857), .B1(n1625), .B2(n1864), .ZN(n1884)
         );
  XNOR2_X1 U1567 ( .A(n1544), .B(n1885), .ZN(n787) );
  AOI221_X1 U1568 ( .B1(n1861), .B2(B[13]), .C1(n1860), .C2(B[12]), .A(n1886), 
        .ZN(n1885) );
  OAI22_X1 U1569 ( .A1(n1628), .A2(n1857), .B1(n1629), .B2(n1864), .ZN(n1886)
         );
  XNOR2_X1 U1570 ( .A(n1544), .B(n1887), .ZN(n786) );
  AOI221_X1 U1571 ( .B1(n1861), .B2(B[14]), .C1(n1860), .C2(B[13]), .A(n1888), 
        .ZN(n1887) );
  OAI22_X1 U1572 ( .A1(n1632), .A2(n1857), .B1(n1633), .B2(n1864), .ZN(n1888)
         );
  XNOR2_X1 U1573 ( .A(n1544), .B(n1889), .ZN(n785) );
  AOI221_X1 U1574 ( .B1(n1861), .B2(B[15]), .C1(n1860), .C2(B[14]), .A(n1890), 
        .ZN(n1889) );
  OAI22_X1 U1575 ( .A1(n1636), .A2(n1857), .B1(n1637), .B2(n1864), .ZN(n1890)
         );
  XNOR2_X1 U1576 ( .A(n1544), .B(n1891), .ZN(n784) );
  AOI221_X1 U1577 ( .B1(n1861), .B2(B[16]), .C1(n1860), .C2(B[15]), .A(n1892), 
        .ZN(n1891) );
  OAI22_X1 U1578 ( .A1(n1640), .A2(n1857), .B1(n1641), .B2(n1864), .ZN(n1892)
         );
  XNOR2_X1 U1579 ( .A(n1544), .B(n1893), .ZN(n783) );
  AOI221_X1 U1580 ( .B1(n1861), .B2(B[17]), .C1(n1860), .C2(B[16]), .A(n1894), 
        .ZN(n1893) );
  OAI22_X1 U1581 ( .A1(n1644), .A2(n1857), .B1(n1645), .B2(n1864), .ZN(n1894)
         );
  XNOR2_X1 U1582 ( .A(n1544), .B(n1895), .ZN(n782) );
  AOI221_X1 U1583 ( .B1(n1861), .B2(B[18]), .C1(n1860), .C2(B[17]), .A(n1896), 
        .ZN(n1895) );
  OAI22_X1 U1584 ( .A1(n1648), .A2(n1857), .B1(n1649), .B2(n1864), .ZN(n1896)
         );
  XNOR2_X1 U1585 ( .A(n1544), .B(n1897), .ZN(n781) );
  AOI221_X1 U1586 ( .B1(n1861), .B2(B[19]), .C1(n1860), .C2(B[18]), .A(n1898), 
        .ZN(n1897) );
  OAI22_X1 U1587 ( .A1(n1652), .A2(n1857), .B1(n1653), .B2(n1864), .ZN(n1898)
         );
  XNOR2_X1 U1588 ( .A(n1544), .B(n1899), .ZN(n780) );
  AOI221_X1 U1589 ( .B1(n1861), .B2(B[20]), .C1(n1860), .C2(B[19]), .A(n1900), 
        .ZN(n1899) );
  OAI22_X1 U1590 ( .A1(n1656), .A2(n1857), .B1(n1657), .B2(n1864), .ZN(n1900)
         );
  XNOR2_X1 U1591 ( .A(A[17]), .B(n1901), .ZN(n779) );
  AOI221_X1 U1592 ( .B1(n1861), .B2(B[21]), .C1(n1860), .C2(B[20]), .A(n1902), 
        .ZN(n1901) );
  OAI22_X1 U1593 ( .A1(n1660), .A2(n1857), .B1(n1661), .B2(n1864), .ZN(n1902)
         );
  XNOR2_X1 U1594 ( .A(A[17]), .B(n1903), .ZN(n778) );
  AOI221_X1 U1595 ( .B1(n1861), .B2(B[22]), .C1(n1860), .C2(B[21]), .A(n1904), 
        .ZN(n1903) );
  OAI22_X1 U1596 ( .A1(n1562), .A2(n1857), .B1(n1564), .B2(n1864), .ZN(n1904)
         );
  XNOR2_X1 U1597 ( .A(A[17]), .B(n1905), .ZN(n777) );
  AOI221_X1 U1598 ( .B1(n1861), .B2(B[23]), .C1(n1860), .C2(B[22]), .A(n1906), 
        .ZN(n1905) );
  OAI22_X1 U1599 ( .A1(n1567), .A2(n1857), .B1(n1568), .B2(n1864), .ZN(n1906)
         );
  XNOR2_X1 U1600 ( .A(A[17]), .B(n1907), .ZN(n776) );
  AOI221_X1 U1601 ( .B1(n1861), .B2(B[23]), .C1(n1860), .C2(n1554), .A(n1908), 
        .ZN(n1907) );
  OAI22_X1 U1602 ( .A1(n1571), .A2(n1857), .B1(n1572), .B2(n1864), .ZN(n1908)
         );
  XNOR2_X1 U1603 ( .A(A[17]), .B(n1909), .ZN(n775) );
  OAI221_X1 U1604 ( .B1(n1556), .B2(n1864), .C1(n1556), .C2(n1857), .A(n1910), 
        .ZN(n1909) );
  OAI21_X1 U1605 ( .B1(n1861), .B2(n1860), .A(n1554), .ZN(n1910) );
  INV_X1 U1606 ( .A(n1914), .ZN(n1911) );
  XNOR2_X1 U1607 ( .A(A[15]), .B(A[16]), .ZN(n1912) );
  XNOR2_X1 U1608 ( .A(A[16]), .B(n1545), .ZN(n1913) );
  XOR2_X1 U1609 ( .A(A[15]), .B(n1547), .Z(n1914) );
  XNOR2_X1 U1610 ( .A(n1915), .B(n1543), .ZN(n774) );
  OAI22_X1 U1611 ( .A1(n1574), .A2(n1916), .B1(n1574), .B2(n1917), .ZN(n1915)
         );
  XNOR2_X1 U1612 ( .A(n1918), .B(n1543), .ZN(n773) );
  OAI222_X1 U1613 ( .A1(n1578), .A2(n1916), .B1(n1574), .B2(n1919), .C1(n1580), 
        .C2(n1917), .ZN(n1918) );
  INV_X1 U1614 ( .A(n1920), .ZN(n1919) );
  INV_X1 U1615 ( .A(n1921), .ZN(n1916) );
  XNOR2_X1 U1616 ( .A(n1542), .B(n1922), .ZN(n772) );
  AOI221_X1 U1617 ( .B1(n1921), .B2(B[2]), .C1(n1920), .C2(B[1]), .A(n1923), 
        .ZN(n1922) );
  OAI22_X1 U1618 ( .A1(n1585), .A2(n1917), .B1(n1574), .B2(n1924), .ZN(n1923)
         );
  XNOR2_X1 U1619 ( .A(n1542), .B(n1925), .ZN(n771) );
  AOI221_X1 U1620 ( .B1(n1921), .B2(B[3]), .C1(n1920), .C2(B[2]), .A(n1926), 
        .ZN(n1925) );
  OAI22_X1 U1621 ( .A1(n1589), .A2(n1917), .B1(n1578), .B2(n1924), .ZN(n1926)
         );
  XNOR2_X1 U1622 ( .A(n1542), .B(n1927), .ZN(n770) );
  AOI221_X1 U1623 ( .B1(n1921), .B2(B[4]), .C1(n1920), .C2(B[3]), .A(n1928), 
        .ZN(n1927) );
  OAI22_X1 U1624 ( .A1(n1592), .A2(n1917), .B1(n1593), .B2(n1924), .ZN(n1928)
         );
  XNOR2_X1 U1625 ( .A(n1542), .B(n1929), .ZN(n769) );
  AOI221_X1 U1626 ( .B1(n1921), .B2(B[5]), .C1(n1920), .C2(B[4]), .A(n1930), 
        .ZN(n1929) );
  OAI22_X1 U1627 ( .A1(n1596), .A2(n1917), .B1(n1597), .B2(n1924), .ZN(n1930)
         );
  XNOR2_X1 U1628 ( .A(n1542), .B(n1931), .ZN(n768) );
  AOI221_X1 U1629 ( .B1(n1921), .B2(B[6]), .C1(n1920), .C2(B[5]), .A(n1932), 
        .ZN(n1931) );
  OAI22_X1 U1630 ( .A1(n1600), .A2(n1917), .B1(n1601), .B2(n1924), .ZN(n1932)
         );
  XNOR2_X1 U1631 ( .A(n1542), .B(n1933), .ZN(n767) );
  AOI221_X1 U1632 ( .B1(n1921), .B2(B[7]), .C1(n1920), .C2(B[6]), .A(n1934), 
        .ZN(n1933) );
  OAI22_X1 U1633 ( .A1(n1604), .A2(n1917), .B1(n1605), .B2(n1924), .ZN(n1934)
         );
  XNOR2_X1 U1634 ( .A(n1542), .B(n1935), .ZN(n766) );
  AOI221_X1 U1635 ( .B1(n1921), .B2(B[8]), .C1(n1920), .C2(B[7]), .A(n1936), 
        .ZN(n1935) );
  OAI22_X1 U1636 ( .A1(n1608), .A2(n1917), .B1(n1609), .B2(n1924), .ZN(n1936)
         );
  XNOR2_X1 U1637 ( .A(n1542), .B(n1937), .ZN(n765) );
  AOI221_X1 U1638 ( .B1(n1921), .B2(B[9]), .C1(n1920), .C2(B[8]), .A(n1938), 
        .ZN(n1937) );
  OAI22_X1 U1639 ( .A1(n1612), .A2(n1917), .B1(n1613), .B2(n1924), .ZN(n1938)
         );
  XNOR2_X1 U1640 ( .A(n1542), .B(n1939), .ZN(n764) );
  AOI221_X1 U1641 ( .B1(n1921), .B2(B[10]), .C1(n1920), .C2(B[9]), .A(n1940), 
        .ZN(n1939) );
  OAI22_X1 U1642 ( .A1(n1616), .A2(n1917), .B1(n1617), .B2(n1924), .ZN(n1940)
         );
  XNOR2_X1 U1643 ( .A(n1542), .B(n1941), .ZN(n763) );
  AOI221_X1 U1644 ( .B1(n1921), .B2(B[11]), .C1(n1920), .C2(B[10]), .A(n1942), 
        .ZN(n1941) );
  OAI22_X1 U1645 ( .A1(n1620), .A2(n1917), .B1(n1621), .B2(n1924), .ZN(n1942)
         );
  XNOR2_X1 U1646 ( .A(n1542), .B(n1943), .ZN(n762) );
  AOI221_X1 U1647 ( .B1(n1921), .B2(B[12]), .C1(n1920), .C2(B[11]), .A(n1944), 
        .ZN(n1943) );
  OAI22_X1 U1648 ( .A1(n1624), .A2(n1917), .B1(n1625), .B2(n1924), .ZN(n1944)
         );
  XNOR2_X1 U1649 ( .A(n1542), .B(n1945), .ZN(n761) );
  AOI221_X1 U1650 ( .B1(n1921), .B2(B[13]), .C1(n1920), .C2(B[12]), .A(n1946), 
        .ZN(n1945) );
  OAI22_X1 U1651 ( .A1(n1628), .A2(n1917), .B1(n1629), .B2(n1924), .ZN(n1946)
         );
  XNOR2_X1 U1652 ( .A(n1542), .B(n1947), .ZN(n760) );
  AOI221_X1 U1653 ( .B1(n1921), .B2(B[14]), .C1(n1920), .C2(B[13]), .A(n1948), 
        .ZN(n1947) );
  OAI22_X1 U1654 ( .A1(n1632), .A2(n1917), .B1(n1633), .B2(n1924), .ZN(n1948)
         );
  XNOR2_X1 U1655 ( .A(n1542), .B(n1949), .ZN(n759) );
  AOI221_X1 U1656 ( .B1(n1921), .B2(B[15]), .C1(n1920), .C2(B[14]), .A(n1950), 
        .ZN(n1949) );
  OAI22_X1 U1657 ( .A1(n1636), .A2(n1917), .B1(n1637), .B2(n1924), .ZN(n1950)
         );
  XNOR2_X1 U1658 ( .A(n1542), .B(n1951), .ZN(n758) );
  AOI221_X1 U1659 ( .B1(n1921), .B2(B[16]), .C1(n1920), .C2(B[15]), .A(n1952), 
        .ZN(n1951) );
  OAI22_X1 U1660 ( .A1(n1640), .A2(n1917), .B1(n1641), .B2(n1924), .ZN(n1952)
         );
  XNOR2_X1 U1661 ( .A(n1542), .B(n1953), .ZN(n757) );
  AOI221_X1 U1662 ( .B1(n1921), .B2(B[17]), .C1(n1920), .C2(B[16]), .A(n1954), 
        .ZN(n1953) );
  OAI22_X1 U1663 ( .A1(n1644), .A2(n1917), .B1(n1645), .B2(n1924), .ZN(n1954)
         );
  XNOR2_X1 U1664 ( .A(n1542), .B(n1955), .ZN(n756) );
  AOI221_X1 U1665 ( .B1(n1921), .B2(B[18]), .C1(n1920), .C2(B[17]), .A(n1956), 
        .ZN(n1955) );
  OAI22_X1 U1666 ( .A1(n1648), .A2(n1917), .B1(n1649), .B2(n1924), .ZN(n1956)
         );
  XNOR2_X1 U1667 ( .A(n1542), .B(n1957), .ZN(n755) );
  AOI221_X1 U1668 ( .B1(n1921), .B2(B[19]), .C1(n1920), .C2(B[18]), .A(n1958), 
        .ZN(n1957) );
  OAI22_X1 U1669 ( .A1(n1652), .A2(n1917), .B1(n1653), .B2(n1924), .ZN(n1958)
         );
  XNOR2_X1 U1670 ( .A(n1542), .B(n1959), .ZN(n754) );
  AOI221_X1 U1671 ( .B1(n1921), .B2(B[20]), .C1(n1920), .C2(B[19]), .A(n1960), 
        .ZN(n1959) );
  OAI22_X1 U1672 ( .A1(n1656), .A2(n1917), .B1(n1657), .B2(n1924), .ZN(n1960)
         );
  XNOR2_X1 U1673 ( .A(A[20]), .B(n1961), .ZN(n753) );
  AOI221_X1 U1674 ( .B1(n1921), .B2(B[21]), .C1(n1920), .C2(B[20]), .A(n1962), 
        .ZN(n1961) );
  OAI22_X1 U1675 ( .A1(n1660), .A2(n1917), .B1(n1661), .B2(n1924), .ZN(n1962)
         );
  XNOR2_X1 U1676 ( .A(A[20]), .B(n1963), .ZN(n752) );
  AOI221_X1 U1677 ( .B1(n1921), .B2(B[22]), .C1(n1920), .C2(B[21]), .A(n1964), 
        .ZN(n1963) );
  OAI22_X1 U1678 ( .A1(n1562), .A2(n1917), .B1(n1564), .B2(n1924), .ZN(n1964)
         );
  XNOR2_X1 U1679 ( .A(A[20]), .B(n1965), .ZN(n751) );
  AOI221_X1 U1680 ( .B1(n1921), .B2(n1554), .C1(n1920), .C2(B[22]), .A(n1966), 
        .ZN(n1965) );
  OAI22_X1 U1681 ( .A1(n1567), .A2(n1917), .B1(n1568), .B2(n1924), .ZN(n1966)
         );
  XNOR2_X1 U1682 ( .A(A[20]), .B(n1967), .ZN(n750) );
  AOI221_X1 U1683 ( .B1(n1921), .B2(B[23]), .C1(n1920), .C2(n1554), .A(n1968), 
        .ZN(n1967) );
  OAI22_X1 U1684 ( .A1(n1571), .A2(n1917), .B1(n1572), .B2(n1924), .ZN(n1968)
         );
  XNOR2_X1 U1685 ( .A(A[20]), .B(n1969), .ZN(n749) );
  OAI221_X1 U1686 ( .B1(n1556), .B2(n1924), .C1(n1556), .C2(n1917), .A(n1970), 
        .ZN(n1969) );
  OAI21_X1 U1687 ( .B1(n1921), .B2(n1920), .A(n1554), .ZN(n1970) );
  INV_X1 U1688 ( .A(n1974), .ZN(n1971) );
  XNOR2_X1 U1689 ( .A(A[18]), .B(A[19]), .ZN(n1972) );
  XNOR2_X1 U1690 ( .A(A[19]), .B(n1543), .ZN(n1973) );
  XOR2_X1 U1691 ( .A(A[18]), .B(n1545), .Z(n1974) );
  XNOR2_X1 U1692 ( .A(n1975), .B(n1541), .ZN(n748) );
  OAI22_X1 U1693 ( .A1(n1574), .A2(n1535), .B1(n1574), .B2(n1976), .ZN(n1975)
         );
  XNOR2_X1 U1694 ( .A(n1977), .B(n1541), .ZN(n747) );
  OAI222_X1 U1695 ( .A1(n1578), .A2(n1535), .B1(n1574), .B2(n1534), .C1(n1580), 
        .C2(n1976), .ZN(n1977) );
  INV_X1 U1696 ( .A(n1397), .ZN(n1580) );
  XNOR2_X1 U1697 ( .A(n1540), .B(n1978), .ZN(n746) );
  AOI221_X1 U1698 ( .B1(n1537), .B2(B[2]), .C1(n1536), .C2(B[1]), .A(n1979), 
        .ZN(n1978) );
  OAI22_X1 U1699 ( .A1(n1585), .A2(n1976), .B1(n1574), .B2(n1538), .ZN(n1979)
         );
  INV_X1 U1700 ( .A(n1396), .ZN(n1585) );
  XNOR2_X1 U1701 ( .A(n1540), .B(n1981), .ZN(n745) );
  AOI221_X1 U1702 ( .B1(n1537), .B2(B[3]), .C1(n1536), .C2(B[2]), .A(n1982), 
        .ZN(n1981) );
  OAI22_X1 U1703 ( .A1(n1589), .A2(n1976), .B1(n1578), .B2(n1539), .ZN(n1982)
         );
  XNOR2_X1 U1704 ( .A(n1540), .B(n1983), .ZN(n744) );
  AOI221_X1 U1705 ( .B1(n1537), .B2(B[4]), .C1(n1536), .C2(B[3]), .A(n1984), 
        .ZN(n1983) );
  OAI22_X1 U1706 ( .A1(n1592), .A2(n1976), .B1(n1593), .B2(n1539), .ZN(n1984)
         );
  XNOR2_X1 U1707 ( .A(n1540), .B(n1985), .ZN(n743) );
  AOI221_X1 U1708 ( .B1(n1537), .B2(B[5]), .C1(n1536), .C2(B[4]), .A(n1986), 
        .ZN(n1985) );
  OAI22_X1 U1709 ( .A1(n1596), .A2(n1976), .B1(n1597), .B2(n1539), .ZN(n1986)
         );
  XNOR2_X1 U1710 ( .A(n1540), .B(n1987), .ZN(n742) );
  AOI221_X1 U1711 ( .B1(n1537), .B2(B[6]), .C1(n1536), .C2(B[5]), .A(n1988), 
        .ZN(n1987) );
  OAI22_X1 U1712 ( .A1(n1600), .A2(n1976), .B1(n1601), .B2(n1539), .ZN(n1988)
         );
  XNOR2_X1 U1713 ( .A(n1540), .B(n1989), .ZN(n741) );
  AOI221_X1 U1714 ( .B1(n1537), .B2(B[7]), .C1(n1536), .C2(B[6]), .A(n1990), 
        .ZN(n1989) );
  OAI22_X1 U1715 ( .A1(n1604), .A2(n1976), .B1(n1605), .B2(n1539), .ZN(n1990)
         );
  XNOR2_X1 U1716 ( .A(n1540), .B(n1991), .ZN(n740) );
  AOI221_X1 U1717 ( .B1(n1537), .B2(B[9]), .C1(n1536), .C2(B[8]), .A(n1992), 
        .ZN(n1991) );
  OAI22_X1 U1718 ( .A1(n1612), .A2(n1976), .B1(n1613), .B2(n1539), .ZN(n1992)
         );
  XNOR2_X1 U1719 ( .A(n1540), .B(n1993), .ZN(n739) );
  AOI221_X1 U1720 ( .B1(n1537), .B2(B[10]), .C1(n1536), .C2(B[9]), .A(n1994), 
        .ZN(n1993) );
  OAI22_X1 U1721 ( .A1(n1616), .A2(n1976), .B1(n1617), .B2(n1539), .ZN(n1994)
         );
  XNOR2_X1 U1722 ( .A(n1540), .B(n1995), .ZN(n738) );
  AOI221_X1 U1723 ( .B1(n1537), .B2(B[12]), .C1(n1536), .C2(B[11]), .A(n1996), 
        .ZN(n1995) );
  OAI22_X1 U1724 ( .A1(n1624), .A2(n1976), .B1(n1625), .B2(n1539), .ZN(n1996)
         );
  XNOR2_X1 U1725 ( .A(n1540), .B(n1997), .ZN(n737) );
  AOI221_X1 U1726 ( .B1(n1537), .B2(B[13]), .C1(n1536), .C2(B[12]), .A(n1998), 
        .ZN(n1997) );
  OAI22_X1 U1727 ( .A1(n1628), .A2(n1976), .B1(n1629), .B2(n1539), .ZN(n1998)
         );
  XNOR2_X1 U1728 ( .A(n1540), .B(n1999), .ZN(n736) );
  AOI221_X1 U1729 ( .B1(n1537), .B2(B[14]), .C1(n1536), .C2(B[13]), .A(n2000), 
        .ZN(n1999) );
  OAI22_X1 U1730 ( .A1(n1632), .A2(n1976), .B1(n1633), .B2(n1539), .ZN(n2000)
         );
  XNOR2_X1 U1731 ( .A(n1540), .B(n2001), .ZN(n735) );
  AOI221_X1 U1732 ( .B1(n1537), .B2(B[15]), .C1(n1536), .C2(B[14]), .A(n2002), 
        .ZN(n2001) );
  OAI22_X1 U1733 ( .A1(n1636), .A2(n1976), .B1(n1637), .B2(n1539), .ZN(n2002)
         );
  XNOR2_X1 U1734 ( .A(n1540), .B(n2003), .ZN(n734) );
  AOI221_X1 U1735 ( .B1(n1537), .B2(B[16]), .C1(n1536), .C2(B[15]), .A(n2004), 
        .ZN(n2003) );
  OAI22_X1 U1736 ( .A1(n1640), .A2(n1976), .B1(n1641), .B2(n1538), .ZN(n2004)
         );
  XNOR2_X1 U1737 ( .A(n1540), .B(n2005), .ZN(n733) );
  AOI221_X1 U1738 ( .B1(n1537), .B2(B[18]), .C1(n1536), .C2(B[17]), .A(n2006), 
        .ZN(n2005) );
  OAI22_X1 U1739 ( .A1(n1648), .A2(n1976), .B1(n1649), .B2(n1538), .ZN(n2006)
         );
  XNOR2_X1 U1740 ( .A(n1540), .B(n2007), .ZN(n732) );
  AOI221_X1 U1741 ( .B1(n1537), .B2(B[19]), .C1(n1536), .C2(B[18]), .A(n2008), 
        .ZN(n2007) );
  OAI22_X1 U1742 ( .A1(n1652), .A2(n1976), .B1(n1653), .B2(n1538), .ZN(n2008)
         );
  XNOR2_X1 U1743 ( .A(n1540), .B(n2009), .ZN(n731) );
  AOI221_X1 U1744 ( .B1(n1537), .B2(B[20]), .C1(n1536), .C2(B[19]), .A(n2010), 
        .ZN(n2009) );
  OAI22_X1 U1745 ( .A1(n1656), .A2(n1976), .B1(n1657), .B2(n1538), .ZN(n2010)
         );
  XNOR2_X1 U1746 ( .A(A[23]), .B(n2011), .ZN(n730) );
  AOI221_X1 U1747 ( .B1(n1537), .B2(B[21]), .C1(n1536), .C2(B[20]), .A(n2012), 
        .ZN(n2011) );
  OAI22_X1 U1748 ( .A1(n1660), .A2(n1976), .B1(n1661), .B2(n1538), .ZN(n2012)
         );
  XNOR2_X1 U1749 ( .A(A[23]), .B(n2013), .ZN(n729) );
  AOI221_X1 U1750 ( .B1(n1537), .B2(B[22]), .C1(n1536), .C2(B[21]), .A(n2014), 
        .ZN(n2013) );
  OAI22_X1 U1751 ( .A1(n1562), .A2(n1976), .B1(n1564), .B2(n1538), .ZN(n2014)
         );
  INV_X1 U1752 ( .A(B[20]), .ZN(n1564) );
  INV_X1 U1753 ( .A(n1376), .ZN(n1562) );
  XNOR2_X1 U1754 ( .A(n519), .B(n2015), .ZN(n506) );
  INV_X1 U1755 ( .A(n493), .ZN(n479) );
  NOR2_X1 U1756 ( .A1(n2015), .A2(n519), .ZN(n493) );
  XOR2_X1 U1757 ( .A(n2016), .B(n1674), .Z(n2015) );
  OAI221_X1 U1758 ( .B1(n1563), .B2(n1556), .C1(n1561), .C2(n1556), .A(n2017), 
        .ZN(n2016) );
  OAI21_X1 U1759 ( .B1(n1558), .B2(n1559), .A(n1554), .ZN(n2017) );
  INV_X1 U1760 ( .A(n454), .ZN(n442) );
  XOR2_X1 U1761 ( .A(n1540), .B(n2018), .Z(n454) );
  AOI221_X1 U1762 ( .B1(n1537), .B2(B[8]), .C1(n1536), .C2(B[7]), .A(n2019), 
        .ZN(n2018) );
  OAI22_X1 U1763 ( .A1(n1608), .A2(n1976), .B1(n1609), .B2(n1538), .ZN(n2019)
         );
  INV_X1 U1764 ( .A(n421), .ZN(n411) );
  XOR2_X1 U1765 ( .A(n1540), .B(n2020), .Z(n421) );
  AOI221_X1 U1766 ( .B1(n1537), .B2(B[11]), .C1(n1536), .C2(B[10]), .A(n2021), 
        .ZN(n2020) );
  OAI22_X1 U1767 ( .A1(n1620), .A2(n1976), .B1(n1621), .B2(n1538), .ZN(n2021)
         );
  INV_X1 U1768 ( .A(n387), .ZN(n395) );
  INV_X1 U1769 ( .A(n374), .ZN(n368) );
  XOR2_X1 U1770 ( .A(n1540), .B(n2022), .Z(n374) );
  AOI221_X1 U1771 ( .B1(n1537), .B2(B[17]), .C1(n1536), .C2(B[16]), .A(n2023), 
        .ZN(n2022) );
  OAI22_X1 U1772 ( .A1(n1644), .A2(n1976), .B1(n1645), .B2(n1538), .ZN(n2023)
         );
  INV_X1 U1773 ( .A(n356), .ZN(n360) );
  INV_X1 U1774 ( .A(n2024), .ZN(n351) );
  OAI222_X1 U1775 ( .A1(n2025), .A2(n2026), .B1(n2025), .B2(n2027), .C1(n2027), 
        .C2(n2026), .ZN(n326) );
  INV_X1 U1776 ( .A(n550), .ZN(n2027) );
  XNOR2_X1 U1777 ( .A(n1674), .B(n2028), .ZN(n2026) );
  AOI221_X1 U1778 ( .B1(B[21]), .B2(n1558), .C1(B[20]), .C2(n1559), .A(n2029), 
        .ZN(n2028) );
  OAI22_X1 U1779 ( .A1(n1561), .A2(n1660), .B1(n1563), .B2(n1661), .ZN(n2029)
         );
  INV_X1 U1780 ( .A(B[19]), .ZN(n1661) );
  INV_X1 U1781 ( .A(n1377), .ZN(n1660) );
  AOI222_X1 U1782 ( .A1(n2030), .A2(n2031), .B1(n2030), .B2(n564), .C1(n564), 
        .C2(n2031), .ZN(n2025) );
  XNOR2_X1 U1783 ( .A(A[2]), .B(n2032), .ZN(n2031) );
  AOI221_X1 U1784 ( .B1(B[20]), .B2(n1558), .C1(B[19]), .C2(n1559), .A(n2033), 
        .ZN(n2032) );
  OAI22_X1 U1785 ( .A1(n1561), .A2(n1656), .B1(n1563), .B2(n1657), .ZN(n2033)
         );
  INV_X1 U1786 ( .A(B[18]), .ZN(n1657) );
  INV_X1 U1787 ( .A(n1378), .ZN(n1656) );
  INV_X1 U1788 ( .A(n2034), .ZN(n2030) );
  AOI222_X1 U1789 ( .A1(n2035), .A2(n2036), .B1(n2035), .B2(n576), .C1(n576), 
        .C2(n2036), .ZN(n2034) );
  XNOR2_X1 U1790 ( .A(A[2]), .B(n2037), .ZN(n2036) );
  AOI221_X1 U1791 ( .B1(B[19]), .B2(n1558), .C1(B[18]), .C2(n1559), .A(n2038), 
        .ZN(n2037) );
  OAI22_X1 U1792 ( .A1(n1561), .A2(n1652), .B1(n1563), .B2(n1653), .ZN(n2038)
         );
  INV_X1 U1793 ( .A(B[17]), .ZN(n1653) );
  INV_X1 U1794 ( .A(n1379), .ZN(n1652) );
  OAI222_X1 U1795 ( .A1(n2039), .A2(n2040), .B1(n2039), .B2(n2041), .C1(n2041), 
        .C2(n2040), .ZN(n2035) );
  INV_X1 U1796 ( .A(n588), .ZN(n2041) );
  XNOR2_X1 U1797 ( .A(n1674), .B(n2042), .ZN(n2040) );
  AOI221_X1 U1798 ( .B1(B[18]), .B2(n1558), .C1(B[17]), .C2(n1559), .A(n2043), 
        .ZN(n2042) );
  OAI22_X1 U1799 ( .A1(n1561), .A2(n1648), .B1(n1563), .B2(n1649), .ZN(n2043)
         );
  INV_X1 U1800 ( .A(B[16]), .ZN(n1649) );
  INV_X1 U1801 ( .A(n1380), .ZN(n1648) );
  AOI222_X1 U1802 ( .A1(n2044), .A2(n2045), .B1(n2044), .B2(n600), .C1(n600), 
        .C2(n2045), .ZN(n2039) );
  XNOR2_X1 U1803 ( .A(A[2]), .B(n2046), .ZN(n2045) );
  AOI221_X1 U1804 ( .B1(B[17]), .B2(n1558), .C1(B[16]), .C2(n1559), .A(n2047), 
        .ZN(n2046) );
  OAI22_X1 U1805 ( .A1(n1561), .A2(n1644), .B1(n1563), .B2(n1645), .ZN(n2047)
         );
  INV_X1 U1806 ( .A(B[15]), .ZN(n1645) );
  INV_X1 U1807 ( .A(n1381), .ZN(n1644) );
  OAI222_X1 U1808 ( .A1(n2048), .A2(n2049), .B1(n2048), .B2(n2050), .C1(n2050), 
        .C2(n2049), .ZN(n2044) );
  INV_X1 U1809 ( .A(n610), .ZN(n2050) );
  XNOR2_X1 U1810 ( .A(n1674), .B(n2051), .ZN(n2049) );
  AOI221_X1 U1811 ( .B1(B[16]), .B2(n1558), .C1(B[15]), .C2(n1559), .A(n2052), 
        .ZN(n2051) );
  OAI22_X1 U1812 ( .A1(n1561), .A2(n1640), .B1(n1563), .B2(n1641), .ZN(n2052)
         );
  INV_X1 U1813 ( .A(B[14]), .ZN(n1641) );
  INV_X1 U1814 ( .A(n1382), .ZN(n1640) );
  AOI222_X1 U1815 ( .A1(n2053), .A2(n2054), .B1(n2053), .B2(n620), .C1(n620), 
        .C2(n2054), .ZN(n2048) );
  XNOR2_X1 U1816 ( .A(A[2]), .B(n2055), .ZN(n2054) );
  AOI221_X1 U1817 ( .B1(B[15]), .B2(n1558), .C1(B[14]), .C2(n1559), .A(n2056), 
        .ZN(n2055) );
  OAI22_X1 U1818 ( .A1(n1561), .A2(n1636), .B1(n1563), .B2(n1637), .ZN(n2056)
         );
  INV_X1 U1819 ( .A(B[13]), .ZN(n1637) );
  INV_X1 U1820 ( .A(n1383), .ZN(n1636) );
  OAI222_X1 U1821 ( .A1(n2057), .A2(n2058), .B1(n2057), .B2(n2059), .C1(n2059), 
        .C2(n2058), .ZN(n2053) );
  INV_X1 U1822 ( .A(n630), .ZN(n2059) );
  XNOR2_X1 U1823 ( .A(n1674), .B(n2060), .ZN(n2058) );
  AOI221_X1 U1824 ( .B1(B[14]), .B2(n1558), .C1(B[13]), .C2(n1559), .A(n2061), 
        .ZN(n2060) );
  OAI22_X1 U1825 ( .A1(n1561), .A2(n1632), .B1(n1563), .B2(n1633), .ZN(n2061)
         );
  INV_X1 U1826 ( .A(B[12]), .ZN(n1633) );
  INV_X1 U1827 ( .A(n1384), .ZN(n1632) );
  AOI222_X1 U1828 ( .A1(n2062), .A2(n2063), .B1(n2062), .B2(n638), .C1(n638), 
        .C2(n2063), .ZN(n2057) );
  XNOR2_X1 U1829 ( .A(A[2]), .B(n2064), .ZN(n2063) );
  AOI221_X1 U1830 ( .B1(B[13]), .B2(n1558), .C1(B[12]), .C2(n1559), .A(n2065), 
        .ZN(n2064) );
  OAI22_X1 U1831 ( .A1(n1561), .A2(n1628), .B1(n1563), .B2(n1629), .ZN(n2065)
         );
  INV_X1 U1832 ( .A(B[11]), .ZN(n1629) );
  INV_X1 U1833 ( .A(n1385), .ZN(n1628) );
  OAI222_X1 U1834 ( .A1(n2066), .A2(n2067), .B1(n2066), .B2(n2068), .C1(n2068), 
        .C2(n2067), .ZN(n2062) );
  INV_X1 U1835 ( .A(n646), .ZN(n2068) );
  XNOR2_X1 U1836 ( .A(n1674), .B(n2069), .ZN(n2067) );
  AOI221_X1 U1837 ( .B1(B[12]), .B2(n1558), .C1(B[11]), .C2(n1559), .A(n2070), 
        .ZN(n2069) );
  OAI22_X1 U1838 ( .A1(n1561), .A2(n1624), .B1(n1563), .B2(n1625), .ZN(n2070)
         );
  INV_X1 U1839 ( .A(B[10]), .ZN(n1625) );
  INV_X1 U1840 ( .A(n1386), .ZN(n1624) );
  AOI222_X1 U1841 ( .A1(n2071), .A2(n2072), .B1(n2071), .B2(n654), .C1(n654), 
        .C2(n2072), .ZN(n2066) );
  XNOR2_X1 U1842 ( .A(A[2]), .B(n2073), .ZN(n2072) );
  AOI221_X1 U1843 ( .B1(B[11]), .B2(n1558), .C1(B[10]), .C2(n1559), .A(n2074), 
        .ZN(n2073) );
  OAI22_X1 U1844 ( .A1(n1561), .A2(n1620), .B1(n1563), .B2(n1621), .ZN(n2074)
         );
  INV_X1 U1845 ( .A(B[9]), .ZN(n1621) );
  INV_X1 U1846 ( .A(n1387), .ZN(n1620) );
  OAI222_X1 U1847 ( .A1(n2075), .A2(n2076), .B1(n2075), .B2(n2077), .C1(n2077), 
        .C2(n2076), .ZN(n2071) );
  INV_X1 U1848 ( .A(n660), .ZN(n2077) );
  XNOR2_X1 U1849 ( .A(n1674), .B(n2078), .ZN(n2076) );
  AOI221_X1 U1850 ( .B1(B[10]), .B2(n1558), .C1(B[9]), .C2(n1559), .A(n2079), 
        .ZN(n2078) );
  OAI22_X1 U1851 ( .A1(n1561), .A2(n1616), .B1(n1563), .B2(n1617), .ZN(n2079)
         );
  INV_X1 U1852 ( .A(B[8]), .ZN(n1617) );
  INV_X1 U1853 ( .A(n1388), .ZN(n1616) );
  AOI222_X1 U1854 ( .A1(n2080), .A2(n2081), .B1(n2080), .B2(n666), .C1(n666), 
        .C2(n2081), .ZN(n2075) );
  XNOR2_X1 U1855 ( .A(A[2]), .B(n2082), .ZN(n2081) );
  AOI221_X1 U1856 ( .B1(B[9]), .B2(n1558), .C1(B[8]), .C2(n1559), .A(n2083), 
        .ZN(n2082) );
  OAI22_X1 U1857 ( .A1(n1561), .A2(n1612), .B1(n1563), .B2(n1613), .ZN(n2083)
         );
  INV_X1 U1858 ( .A(B[7]), .ZN(n1613) );
  INV_X1 U1859 ( .A(n1389), .ZN(n1612) );
  OAI222_X1 U1860 ( .A1(n2084), .A2(n2085), .B1(n2084), .B2(n2086), .C1(n2086), 
        .C2(n2085), .ZN(n2080) );
  INV_X1 U1861 ( .A(n672), .ZN(n2086) );
  XNOR2_X1 U1862 ( .A(n1674), .B(n2087), .ZN(n2085) );
  AOI221_X1 U1863 ( .B1(B[8]), .B2(n1558), .C1(B[7]), .C2(n1559), .A(n2088), 
        .ZN(n2087) );
  OAI22_X1 U1864 ( .A1(n1561), .A2(n1608), .B1(n1563), .B2(n1609), .ZN(n2088)
         );
  INV_X1 U1865 ( .A(B[6]), .ZN(n1609) );
  INV_X1 U1866 ( .A(n1390), .ZN(n1608) );
  AOI222_X1 U1867 ( .A1(n2089), .A2(n2090), .B1(n2089), .B2(n676), .C1(n676), 
        .C2(n2090), .ZN(n2084) );
  XNOR2_X1 U1868 ( .A(A[2]), .B(n2091), .ZN(n2090) );
  AOI221_X1 U1869 ( .B1(B[7]), .B2(n1558), .C1(B[6]), .C2(n1559), .A(n2092), 
        .ZN(n2091) );
  OAI22_X1 U1870 ( .A1(n1561), .A2(n1604), .B1(n1563), .B2(n1605), .ZN(n2092)
         );
  INV_X1 U1871 ( .A(B[5]), .ZN(n1605) );
  INV_X1 U1872 ( .A(n1391), .ZN(n1604) );
  OAI222_X1 U1873 ( .A1(n2093), .A2(n2094), .B1(n2093), .B2(n2095), .C1(n2095), 
        .C2(n2094), .ZN(n2089) );
  INV_X1 U1874 ( .A(n680), .ZN(n2095) );
  XNOR2_X1 U1875 ( .A(n1674), .B(n2096), .ZN(n2094) );
  AOI221_X1 U1876 ( .B1(B[6]), .B2(n1558), .C1(B[5]), .C2(n1559), .A(n2097), 
        .ZN(n2096) );
  OAI22_X1 U1877 ( .A1(n1561), .A2(n1600), .B1(n1563), .B2(n1601), .ZN(n2097)
         );
  INV_X1 U1878 ( .A(B[4]), .ZN(n1601) );
  INV_X1 U1879 ( .A(n1392), .ZN(n1600) );
  AOI222_X1 U1880 ( .A1(n2098), .A2(n2099), .B1(n2098), .B2(n684), .C1(n684), 
        .C2(n2099), .ZN(n2093) );
  XNOR2_X1 U1881 ( .A(A[2]), .B(n2100), .ZN(n2099) );
  AOI221_X1 U1882 ( .B1(B[5]), .B2(n1558), .C1(B[4]), .C2(n1559), .A(n2101), 
        .ZN(n2100) );
  OAI22_X1 U1883 ( .A1(n1561), .A2(n1596), .B1(n1563), .B2(n1597), .ZN(n2101)
         );
  INV_X1 U1884 ( .A(B[3]), .ZN(n1597) );
  INV_X1 U1885 ( .A(n1393), .ZN(n1596) );
  OAI222_X1 U1886 ( .A1(n2102), .A2(n2103), .B1(n2102), .B2(n2104), .C1(n2104), 
        .C2(n2103), .ZN(n2098) );
  INV_X1 U1887 ( .A(n686), .ZN(n2104) );
  XNOR2_X1 U1888 ( .A(n1674), .B(n2105), .ZN(n2103) );
  AOI221_X1 U1889 ( .B1(B[4]), .B2(n1558), .C1(B[3]), .C2(n1559), .A(n2106), 
        .ZN(n2105) );
  OAI22_X1 U1890 ( .A1(n1561), .A2(n1592), .B1(n1563), .B2(n1593), .ZN(n2106)
         );
  INV_X1 U1891 ( .A(B[2]), .ZN(n1593) );
  INV_X1 U1892 ( .A(n1394), .ZN(n1592) );
  AOI222_X1 U1893 ( .A1(n2107), .A2(n2108), .B1(n2107), .B2(n688), .C1(n688), 
        .C2(n2108), .ZN(n2102) );
  XNOR2_X1 U1894 ( .A(A[2]), .B(n2109), .ZN(n2108) );
  AOI221_X1 U1895 ( .B1(B[3]), .B2(n1558), .C1(B[2]), .C2(n1559), .A(n2110), 
        .ZN(n2109) );
  OAI22_X1 U1896 ( .A1(n1561), .A2(n1589), .B1(n1563), .B2(n1578), .ZN(n2110)
         );
  INV_X1 U1897 ( .A(B[1]), .ZN(n1578) );
  INV_X1 U1898 ( .A(n1395), .ZN(n1589) );
  AND2_X1 U1899 ( .A1(n2114), .A2(n2115), .ZN(n2107) );
  AOI211_X1 U1900 ( .C1(B[1]), .C2(n1558), .A(n2116), .B(B[0]), .ZN(n2115) );
  INV_X1 U1901 ( .A(n2117), .ZN(n2116) );
  AOI22_X1 U1902 ( .A1(n1558), .A2(B[2]), .B1(n2118), .B2(n1397), .ZN(n2117)
         );
  INV_X1 U1903 ( .A(A[0]), .ZN(n2112) );
  AOI221_X1 U1904 ( .B1(B[1]), .B2(n1559), .C1(n1396), .C2(n2118), .A(n1674), 
        .ZN(n2114) );
  INV_X1 U1905 ( .A(n1561), .ZN(n2118) );
  XNOR2_X1 U1906 ( .A(A[1]), .B(n1674), .ZN(n2111) );
  INV_X1 U1907 ( .A(A[2]), .ZN(n1674) );
  INV_X1 U1908 ( .A(A[1]), .ZN(n2113) );
  AOI21_X1 U1909 ( .B1(n2119), .B2(n2120), .A(n2121), .ZN(PRODUCT[47]) );
  OAI22_X1 U1910 ( .A1(n2122), .A2(n2123), .B1(n2122), .B2(n2124), .ZN(n2121)
         );
  INV_X1 U1911 ( .A(n2120), .ZN(n2124) );
  AOI222_X1 U1912 ( .A1(n2024), .A2(n303), .B1(n2123), .B2(n303), .C1(n2024), 
        .C2(n2123), .ZN(n2122) );
  XOR2_X1 U1913 ( .A(n1541), .B(n2125), .Z(n2024) );
  AOI221_X1 U1914 ( .B1(n1537), .B2(B[23]), .C1(n1536), .C2(B[22]), .A(n2126), 
        .ZN(n2125) );
  OAI22_X1 U1915 ( .A1(n1567), .A2(n1976), .B1(n1568), .B2(n1538), .ZN(n2126)
         );
  INV_X1 U1916 ( .A(B[21]), .ZN(n1568) );
  INV_X1 U1917 ( .A(n1375), .ZN(n1567) );
  XOR2_X1 U1918 ( .A(n2127), .B(n1541), .Z(n2120) );
  OAI221_X1 U1919 ( .B1(n1556), .B2(n1539), .C1(n1556), .C2(n1976), .A(n2128), 
        .ZN(n2127) );
  OAI21_X1 U1920 ( .B1(n1537), .B2(n1536), .A(n1554), .ZN(n2128) );
  INV_X1 U1921 ( .A(n2123), .ZN(n2119) );
  XOR2_X1 U1922 ( .A(A[23]), .B(n2129), .Z(n2123) );
  AOI221_X1 U1923 ( .B1(n1537), .B2(n1554), .C1(n1536), .C2(n1554), .A(n2130), 
        .ZN(n2129) );
  OAI22_X1 U1924 ( .A1(n1571), .A2(n1976), .B1(n1572), .B2(n1538), .ZN(n2130)
         );
  NAND3_X1 U1925 ( .A1(n2131), .A2(n2132), .A3(n2133), .ZN(n1980) );
  INV_X1 U1926 ( .A(B[22]), .ZN(n1572) );
  INV_X1 U1927 ( .A(n1374), .ZN(n1571) );
  XNOR2_X1 U1928 ( .A(A[21]), .B(A[22]), .ZN(n2133) );
  INV_X1 U1929 ( .A(n2131), .ZN(n2134) );
  XOR2_X1 U1930 ( .A(A[21]), .B(n1543), .Z(n2131) );
  XNOR2_X1 U1931 ( .A(A[22]), .B(n1541), .ZN(n2132) );
endmodule


module iir_filter_DW02_mult_1 ( A, B, PRODUCT, TC );
  input [23:0] A;
  input [23:0] B;
  output [47:0] PRODUCT;
  input TC;
  wire   n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n351, n352, n353, n354, n355, n356, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n906, n907, n908, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134;

  FA_X1 U182 ( .A(n351), .B(n352), .CI(n304), .CO(n303), .S(PRODUCT[44]) );
  FA_X1 U183 ( .A(n353), .B(n354), .CI(n305), .CO(n304), .S(PRODUCT[43]) );
  FA_X1 U184 ( .A(n355), .B(n358), .CI(n306), .CO(n305), .S(PRODUCT[42]) );
  FA_X1 U185 ( .A(n359), .B(n361), .CI(n307), .CO(n306), .S(PRODUCT[41]) );
  FA_X1 U186 ( .A(n362), .B(n364), .CI(n308), .CO(n307), .S(PRODUCT[40]) );
  FA_X1 U187 ( .A(n365), .B(n370), .CI(n309), .CO(n308), .S(PRODUCT[39]) );
  FA_X1 U188 ( .A(n371), .B(n375), .CI(n310), .CO(n309), .S(PRODUCT[38]) );
  FA_X1 U189 ( .A(n376), .B(n381), .CI(n311), .CO(n310), .S(PRODUCT[37]) );
  FA_X1 U190 ( .A(n382), .B(n389), .CI(n312), .CO(n311), .S(PRODUCT[36]) );
  FA_X1 U191 ( .A(n390), .B(n396), .CI(n313), .CO(n312), .S(PRODUCT[35]) );
  FA_X1 U192 ( .A(n397), .B(n403), .CI(n314), .CO(n313), .S(PRODUCT[34]) );
  FA_X1 U193 ( .A(n404), .B(n413), .CI(n315), .CO(n314), .S(PRODUCT[33]) );
  FA_X1 U194 ( .A(n414), .B(n422), .CI(n316), .CO(n315), .S(PRODUCT[32]) );
  FA_X1 U195 ( .A(n423), .B(n432), .CI(n317), .CO(n316), .S(PRODUCT[31]) );
  FA_X1 U196 ( .A(n433), .B(n444), .CI(n318), .CO(n317), .S(PRODUCT[30]) );
  FA_X1 U197 ( .A(n445), .B(n455), .CI(n319), .CO(n318), .S(PRODUCT[29]) );
  FA_X1 U198 ( .A(n456), .B(n467), .CI(n320), .CO(n319), .S(PRODUCT[28]) );
  FA_X1 U199 ( .A(n468), .B(n481), .CI(n321), .CO(n320), .S(PRODUCT[27]) );
  FA_X1 U200 ( .A(n482), .B(n494), .CI(n322), .CO(n321), .S(PRODUCT[26]) );
  FA_X1 U201 ( .A(n495), .B(n507), .CI(n323), .CO(n322), .S(PRODUCT[25]) );
  FA_X1 U202 ( .A(n508), .B(n906), .CI(n324), .CO(n323), .S(PRODUCT[24]) );
  FA_X1 U203 ( .A(n907), .B(n522), .CI(n325), .CO(n324), .S(PRODUCT[23]) );
  FA_X1 U204 ( .A(n908), .B(n536), .CI(n326), .CO(n325), .S(PRODUCT[22]) );
  FA_X1 U235 ( .A(n356), .B(n749), .CI(n729), .CO(n352), .S(n353) );
  FA_X1 U236 ( .A(n730), .B(n360), .CI(n750), .CO(n354), .S(n355) );
  FA_X1 U238 ( .A(n360), .B(n731), .CI(n751), .CO(n358), .S(n359) );
  FA_X1 U240 ( .A(n752), .B(n363), .CI(n366), .CO(n361), .S(n362) );
  FA_X1 U241 ( .A(n368), .B(n775), .CI(n732), .CO(n356), .S(n363) );
  FA_X1 U242 ( .A(n776), .B(n753), .CI(n367), .CO(n364), .S(n365) );
  FA_X1 U243 ( .A(n733), .B(n374), .CI(n372), .CO(n366), .S(n367) );
  FA_X1 U245 ( .A(n373), .B(n377), .CI(n777), .CO(n370), .S(n371) );
  FA_X1 U246 ( .A(n374), .B(n379), .CI(n754), .CO(n372), .S(n373) );
  FA_X1 U248 ( .A(n778), .B(n378), .CI(n383), .CO(n375), .S(n376) );
  FA_X1 U249 ( .A(n385), .B(n380), .CI(n755), .CO(n377), .S(n378) );
  FA_X1 U250 ( .A(n387), .B(n801), .CI(n734), .CO(n379), .S(n380) );
  FA_X1 U251 ( .A(n802), .B(n779), .CI(n384), .CO(n381), .S(n382) );
  FA_X1 U252 ( .A(n386), .B(n393), .CI(n391), .CO(n383), .S(n384) );
  FA_X1 U253 ( .A(n735), .B(n395), .CI(n756), .CO(n385), .S(n386) );
  FA_X1 U255 ( .A(n392), .B(n398), .CI(n803), .CO(n389), .S(n390) );
  FA_X1 U256 ( .A(n394), .B(n400), .CI(n780), .CO(n391), .S(n392) );
  FA_X1 U257 ( .A(n395), .B(n736), .CI(n757), .CO(n393), .S(n394) );
  FA_X1 U259 ( .A(n804), .B(n399), .CI(n405), .CO(n396), .S(n397) );
  FA_X1 U260 ( .A(n407), .B(n401), .CI(n781), .CO(n398), .S(n399) );
  FA_X1 U261 ( .A(n758), .B(n402), .CI(n409), .CO(n400), .S(n401) );
  FA_X1 U262 ( .A(n411), .B(n827), .CI(n737), .CO(n387), .S(n402) );
  FA_X1 U263 ( .A(n828), .B(n805), .CI(n406), .CO(n403), .S(n404) );
  FA_X1 U264 ( .A(n408), .B(n417), .CI(n415), .CO(n405), .S(n406) );
  FA_X1 U265 ( .A(n410), .B(n759), .CI(n782), .CO(n407), .S(n408) );
  FA_X1 U266 ( .A(n738), .B(n421), .CI(n419), .CO(n409), .S(n410) );
  FA_X1 U268 ( .A(n416), .B(n424), .CI(n829), .CO(n413), .S(n414) );
  FA_X1 U269 ( .A(n418), .B(n426), .CI(n806), .CO(n415), .S(n416) );
  FA_X1 U270 ( .A(n420), .B(n428), .CI(n783), .CO(n417), .S(n418) );
  FA_X1 U271 ( .A(n421), .B(n430), .CI(n760), .CO(n419), .S(n420) );
  FA_X1 U273 ( .A(n830), .B(n425), .CI(n434), .CO(n422), .S(n423) );
  FA_X1 U274 ( .A(n436), .B(n427), .CI(n807), .CO(n424), .S(n425) );
  FA_X1 U275 ( .A(n784), .B(n429), .CI(n438), .CO(n426), .S(n427) );
  FA_X1 U276 ( .A(n440), .B(n431), .CI(n761), .CO(n428), .S(n429) );
  FA_X1 U277 ( .A(n442), .B(n853), .CI(n739), .CO(n430), .S(n431) );
  FA_X1 U278 ( .A(n854), .B(n831), .CI(n435), .CO(n432), .S(n433) );
  FA_X1 U279 ( .A(n437), .B(n448), .CI(n446), .CO(n434), .S(n435) );
  FA_X1 U280 ( .A(n439), .B(n785), .CI(n808), .CO(n436), .S(n437) );
  FA_X1 U281 ( .A(n441), .B(n452), .CI(n450), .CO(n438), .S(n439) );
  FA_X1 U282 ( .A(n740), .B(n454), .CI(n762), .CO(n440), .S(n441) );
  FA_X1 U284 ( .A(n447), .B(n457), .CI(n855), .CO(n444), .S(n445) );
  FA_X1 U285 ( .A(n449), .B(n459), .CI(n832), .CO(n446), .S(n447) );
  FA_X1 U286 ( .A(n451), .B(n461), .CI(n809), .CO(n448), .S(n449) );
  FA_X1 U287 ( .A(n453), .B(n463), .CI(n786), .CO(n450), .S(n451) );
  FA_X1 U288 ( .A(n454), .B(n465), .CI(n763), .CO(n452), .S(n453) );
  FA_X1 U290 ( .A(n856), .B(n458), .CI(n469), .CO(n455), .S(n456) );
  FA_X1 U291 ( .A(n471), .B(n460), .CI(n833), .CO(n457), .S(n458) );
  FA_X1 U292 ( .A(n810), .B(n462), .CI(n473), .CO(n459), .S(n460) );
  FA_X1 U293 ( .A(n475), .B(n464), .CI(n787), .CO(n461), .S(n462) );
  FA_X1 U294 ( .A(n764), .B(n466), .CI(n477), .CO(n463), .S(n464) );
  FA_X1 U295 ( .A(n479), .B(n879), .CI(n741), .CO(n465), .S(n466) );
  FA_X1 U296 ( .A(n880), .B(n857), .CI(n470), .CO(n467), .S(n468) );
  FA_X1 U297 ( .A(n472), .B(n485), .CI(n483), .CO(n469), .S(n470) );
  FA_X1 U298 ( .A(n474), .B(n811), .CI(n834), .CO(n471), .S(n472) );
  FA_X1 U299 ( .A(n476), .B(n489), .CI(n487), .CO(n473), .S(n474) );
  FA_X1 U300 ( .A(n478), .B(n765), .CI(n788), .CO(n475), .S(n476) );
  FA_X1 U301 ( .A(n742), .B(n493), .CI(n491), .CO(n477), .S(n478) );
  FA_X1 U303 ( .A(n484), .B(n858), .CI(n881), .CO(n481), .S(n482) );
  FA_X1 U304 ( .A(n486), .B(n498), .CI(n496), .CO(n483), .S(n484) );
  FA_X1 U305 ( .A(n488), .B(n812), .CI(n835), .CO(n485), .S(n486) );
  FA_X1 U306 ( .A(n490), .B(n502), .CI(n500), .CO(n487), .S(n488) );
  FA_X1 U307 ( .A(n492), .B(n504), .CI(n789), .CO(n489), .S(n490) );
  FA_X1 U308 ( .A(n743), .B(n493), .CI(n766), .CO(n491), .S(n492) );
  FA_X1 U310 ( .A(n497), .B(n509), .CI(n882), .CO(n494), .S(n495) );
  FA_X1 U311 ( .A(n499), .B(n511), .CI(n859), .CO(n496), .S(n497) );
  FA_X1 U312 ( .A(n501), .B(n513), .CI(n836), .CO(n498), .S(n499) );
  FA_X1 U313 ( .A(n503), .B(n515), .CI(n813), .CO(n500), .S(n501) );
  FA_X1 U314 ( .A(n505), .B(n517), .CI(n790), .CO(n502), .S(n503) );
  FA_X1 U315 ( .A(n506), .B(n744), .CI(n767), .CO(n504), .S(n505) );
  FA_X1 U318 ( .A(n883), .B(n510), .CI(n521), .CO(n507), .S(n508) );
  FA_X1 U319 ( .A(n860), .B(n512), .CI(n523), .CO(n509), .S(n510) );
  FA_X1 U320 ( .A(n837), .B(n514), .CI(n525), .CO(n511), .S(n512) );
  FA_X1 U321 ( .A(n814), .B(n516), .CI(n527), .CO(n513), .S(n514) );
  FA_X1 U322 ( .A(n791), .B(n518), .CI(n529), .CO(n515), .S(n516) );
  FA_X1 U323 ( .A(n768), .B(n520), .CI(n531), .CO(n517), .S(n518) );
  HA_X1 U324 ( .A(n533), .B(n745), .CO(n519), .S(n520) );
  FA_X1 U325 ( .A(n884), .B(n524), .CI(n535), .CO(n521), .S(n522) );
  FA_X1 U326 ( .A(n861), .B(n526), .CI(n537), .CO(n523), .S(n524) );
  FA_X1 U327 ( .A(n838), .B(n528), .CI(n539), .CO(n525), .S(n526) );
  FA_X1 U328 ( .A(n815), .B(n530), .CI(n541), .CO(n527), .S(n528) );
  FA_X1 U329 ( .A(n792), .B(n532), .CI(n543), .CO(n529), .S(n530) );
  FA_X1 U330 ( .A(n769), .B(n534), .CI(n545), .CO(n531), .S(n532) );
  HA_X1 U331 ( .A(n547), .B(n746), .CO(n533), .S(n534) );
  FA_X1 U332 ( .A(n885), .B(n538), .CI(n549), .CO(n535), .S(n536) );
  FA_X1 U333 ( .A(n862), .B(n540), .CI(n551), .CO(n537), .S(n538) );
  FA_X1 U334 ( .A(n839), .B(n542), .CI(n553), .CO(n539), .S(n540) );
  FA_X1 U335 ( .A(n816), .B(n544), .CI(n555), .CO(n541), .S(n542) );
  FA_X1 U336 ( .A(n793), .B(n546), .CI(n557), .CO(n543), .S(n544) );
  FA_X1 U337 ( .A(n770), .B(n548), .CI(n559), .CO(n545), .S(n546) );
  HA_X1 U338 ( .A(n561), .B(n747), .CO(n547), .S(n548) );
  FA_X1 U339 ( .A(n886), .B(n552), .CI(n563), .CO(n549), .S(n550) );
  FA_X1 U340 ( .A(n863), .B(n554), .CI(n565), .CO(n551), .S(n552) );
  FA_X1 U341 ( .A(n840), .B(n556), .CI(n567), .CO(n553), .S(n554) );
  FA_X1 U342 ( .A(n817), .B(n558), .CI(n569), .CO(n555), .S(n556) );
  FA_X1 U343 ( .A(n794), .B(n560), .CI(n571), .CO(n557), .S(n558) );
  FA_X1 U344 ( .A(n771), .B(n562), .CI(n573), .CO(n559), .S(n560) );
  HA_X1 U345 ( .A(n748), .B(n1540), .CO(n561), .S(n562) );
  FA_X1 U346 ( .A(n887), .B(n566), .CI(n575), .CO(n563), .S(n564) );
  FA_X1 U347 ( .A(n864), .B(n568), .CI(n577), .CO(n565), .S(n566) );
  FA_X1 U348 ( .A(n841), .B(n570), .CI(n579), .CO(n567), .S(n568) );
  FA_X1 U349 ( .A(n818), .B(n572), .CI(n581), .CO(n569), .S(n570) );
  FA_X1 U350 ( .A(n795), .B(n574), .CI(n583), .CO(n571), .S(n572) );
  HA_X1 U351 ( .A(n585), .B(n772), .CO(n573), .S(n574) );
  FA_X1 U352 ( .A(n888), .B(n578), .CI(n587), .CO(n575), .S(n576) );
  FA_X1 U353 ( .A(n865), .B(n580), .CI(n589), .CO(n577), .S(n578) );
  FA_X1 U354 ( .A(n842), .B(n582), .CI(n591), .CO(n579), .S(n580) );
  FA_X1 U355 ( .A(n819), .B(n584), .CI(n593), .CO(n581), .S(n582) );
  FA_X1 U356 ( .A(n796), .B(n586), .CI(n595), .CO(n583), .S(n584) );
  HA_X1 U357 ( .A(n597), .B(n773), .CO(n585), .S(n586) );
  FA_X1 U358 ( .A(n889), .B(n590), .CI(n599), .CO(n587), .S(n588) );
  FA_X1 U359 ( .A(n866), .B(n592), .CI(n601), .CO(n589), .S(n590) );
  FA_X1 U360 ( .A(n843), .B(n594), .CI(n603), .CO(n591), .S(n592) );
  FA_X1 U361 ( .A(n820), .B(n596), .CI(n605), .CO(n593), .S(n594) );
  FA_X1 U362 ( .A(n797), .B(n598), .CI(n607), .CO(n595), .S(n596) );
  HA_X1 U363 ( .A(n774), .B(n1542), .CO(n597), .S(n598) );
  FA_X1 U364 ( .A(n890), .B(n602), .CI(n609), .CO(n599), .S(n600) );
  FA_X1 U365 ( .A(n867), .B(n604), .CI(n611), .CO(n601), .S(n602) );
  FA_X1 U366 ( .A(n844), .B(n606), .CI(n613), .CO(n603), .S(n604) );
  FA_X1 U367 ( .A(n821), .B(n608), .CI(n615), .CO(n605), .S(n606) );
  HA_X1 U368 ( .A(n617), .B(n798), .CO(n607), .S(n608) );
  FA_X1 U369 ( .A(n891), .B(n612), .CI(n619), .CO(n609), .S(n610) );
  FA_X1 U370 ( .A(n868), .B(n614), .CI(n621), .CO(n611), .S(n612) );
  FA_X1 U371 ( .A(n845), .B(n616), .CI(n623), .CO(n613), .S(n614) );
  FA_X1 U372 ( .A(n822), .B(n618), .CI(n625), .CO(n615), .S(n616) );
  HA_X1 U373 ( .A(n627), .B(n799), .CO(n617), .S(n618) );
  FA_X1 U374 ( .A(n892), .B(n622), .CI(n629), .CO(n619), .S(n620) );
  FA_X1 U375 ( .A(n869), .B(n624), .CI(n631), .CO(n621), .S(n622) );
  FA_X1 U376 ( .A(n846), .B(n626), .CI(n633), .CO(n623), .S(n624) );
  FA_X1 U377 ( .A(n823), .B(n628), .CI(n635), .CO(n625), .S(n626) );
  HA_X1 U378 ( .A(n800), .B(n1544), .CO(n627), .S(n628) );
  FA_X1 U379 ( .A(n893), .B(n632), .CI(n637), .CO(n629), .S(n630) );
  FA_X1 U380 ( .A(n870), .B(n634), .CI(n639), .CO(n631), .S(n632) );
  FA_X1 U381 ( .A(n847), .B(n636), .CI(n641), .CO(n633), .S(n634) );
  HA_X1 U382 ( .A(n643), .B(n824), .CO(n635), .S(n636) );
  FA_X1 U383 ( .A(n894), .B(n640), .CI(n645), .CO(n637), .S(n638) );
  FA_X1 U384 ( .A(n871), .B(n642), .CI(n647), .CO(n639), .S(n640) );
  FA_X1 U385 ( .A(n848), .B(n644), .CI(n649), .CO(n641), .S(n642) );
  HA_X1 U386 ( .A(n651), .B(n825), .CO(n643), .S(n644) );
  FA_X1 U387 ( .A(n895), .B(n648), .CI(n653), .CO(n645), .S(n646) );
  FA_X1 U388 ( .A(n872), .B(n650), .CI(n655), .CO(n647), .S(n648) );
  FA_X1 U389 ( .A(n849), .B(n652), .CI(n657), .CO(n649), .S(n650) );
  HA_X1 U390 ( .A(n826), .B(n1546), .CO(n651), .S(n652) );
  FA_X1 U391 ( .A(n896), .B(n656), .CI(n659), .CO(n653), .S(n654) );
  FA_X1 U392 ( .A(n873), .B(n658), .CI(n661), .CO(n655), .S(n656) );
  HA_X1 U393 ( .A(n663), .B(n850), .CO(n657), .S(n658) );
  FA_X1 U394 ( .A(n897), .B(n662), .CI(n665), .CO(n659), .S(n660) );
  FA_X1 U395 ( .A(n874), .B(n664), .CI(n667), .CO(n661), .S(n662) );
  HA_X1 U396 ( .A(n669), .B(n851), .CO(n663), .S(n664) );
  FA_X1 U397 ( .A(n898), .B(n668), .CI(n671), .CO(n665), .S(n666) );
  FA_X1 U398 ( .A(n875), .B(n670), .CI(n673), .CO(n667), .S(n668) );
  HA_X1 U399 ( .A(n852), .B(n1548), .CO(n669), .S(n670) );
  FA_X1 U400 ( .A(n899), .B(n674), .CI(n675), .CO(n671), .S(n672) );
  HA_X1 U401 ( .A(n677), .B(n876), .CO(n673), .S(n674) );
  FA_X1 U402 ( .A(n900), .B(n678), .CI(n679), .CO(n675), .S(n676) );
  HA_X1 U403 ( .A(n681), .B(n877), .CO(n677), .S(n678) );
  FA_X1 U404 ( .A(n901), .B(n682), .CI(n683), .CO(n679), .S(n680) );
  HA_X1 U405 ( .A(n878), .B(n1550), .CO(n681), .S(n682) );
  HA_X1 U406 ( .A(n685), .B(n902), .CO(n683), .S(n684) );
  HA_X1 U407 ( .A(n687), .B(n903), .CO(n685), .S(n686) );
  HA_X1 U408 ( .A(n904), .B(n1552), .CO(n687), .S(n688) );
  FA_X1 U1112 ( .A(B[22]), .B(n1554), .CI(n706), .CO(n1374), .S(n1375) );
  FA_X1 U1113 ( .A(B[21]), .B(B[22]), .CI(n707), .CO(n706), .S(n1376) );
  FA_X1 U1114 ( .A(B[20]), .B(B[21]), .CI(n708), .CO(n707), .S(n1377) );
  FA_X1 U1115 ( .A(B[19]), .B(B[20]), .CI(n709), .CO(n708), .S(n1378) );
  FA_X1 U1116 ( .A(B[18]), .B(B[19]), .CI(n710), .CO(n709), .S(n1379) );
  FA_X1 U1117 ( .A(B[17]), .B(B[18]), .CI(n711), .CO(n710), .S(n1380) );
  FA_X1 U1118 ( .A(B[16]), .B(B[17]), .CI(n712), .CO(n711), .S(n1381) );
  FA_X1 U1119 ( .A(B[15]), .B(B[16]), .CI(n713), .CO(n712), .S(n1382) );
  FA_X1 U1120 ( .A(B[14]), .B(B[15]), .CI(n714), .CO(n713), .S(n1383) );
  FA_X1 U1121 ( .A(B[13]), .B(B[14]), .CI(n715), .CO(n714), .S(n1384) );
  FA_X1 U1122 ( .A(B[12]), .B(B[13]), .CI(n716), .CO(n715), .S(n1385) );
  FA_X1 U1123 ( .A(B[11]), .B(B[12]), .CI(n717), .CO(n716), .S(n1386) );
  FA_X1 U1124 ( .A(B[10]), .B(B[11]), .CI(n718), .CO(n717), .S(n1387) );
  FA_X1 U1125 ( .A(B[9]), .B(B[10]), .CI(n719), .CO(n718), .S(n1388) );
  FA_X1 U1126 ( .A(B[8]), .B(B[9]), .CI(n720), .CO(n719), .S(n1389) );
  FA_X1 U1127 ( .A(B[7]), .B(B[8]), .CI(n721), .CO(n720), .S(n1390) );
  FA_X1 U1128 ( .A(B[6]), .B(B[7]), .CI(n722), .CO(n721), .S(n1391) );
  FA_X1 U1129 ( .A(B[5]), .B(B[6]), .CI(n723), .CO(n722), .S(n1392) );
  FA_X1 U1130 ( .A(B[4]), .B(B[5]), .CI(n724), .CO(n723), .S(n1393) );
  FA_X1 U1131 ( .A(B[3]), .B(B[4]), .CI(n725), .CO(n724), .S(n1394) );
  FA_X1 U1132 ( .A(B[2]), .B(B[3]), .CI(n726), .CO(n725), .S(n1395) );
  FA_X1 U1133 ( .A(B[1]), .B(B[2]), .CI(n727), .CO(n726), .S(n1396) );
  HA_X1 U1134 ( .A(B[0]), .B(B[1]), .CO(n727), .S(n1397) );
  OR2_X1 U1138 ( .A1(n2134), .A2(n2133), .ZN(n1534) );
  INV_X1 U1139 ( .A(n1534), .ZN(n1536) );
  INV_X1 U1140 ( .A(n1535), .ZN(n1537) );
  BUF_X1 U1141 ( .A(n1980), .Z(n1538) );
  BUF_X1 U1142 ( .A(n1980), .Z(n1539) );
  NAND3_X1 U1143 ( .A1(n1673), .A2(n1672), .A3(n1671), .ZN(n1586) );
  NAND3_X1 U1144 ( .A1(n1854), .A2(n1853), .A3(n1852), .ZN(n1804) );
  NAND3_X1 U1145 ( .A1(n1794), .A2(n1793), .A3(n1792), .ZN(n1744) );
  NAND3_X1 U1146 ( .A1(n1734), .A2(n1733), .A3(n1732), .ZN(n1684) );
  NAND3_X1 U1147 ( .A1(n2111), .A2(n2112), .A3(n2113), .ZN(n1563) );
  NAND2_X1 U1148 ( .A1(n1911), .A2(n1913), .ZN(n1857) );
  NAND2_X1 U1149 ( .A1(n1851), .A2(n1853), .ZN(n1797) );
  NAND2_X1 U1150 ( .A1(n1791), .A2(n1793), .ZN(n1737) );
  NAND2_X1 U1151 ( .A1(n1731), .A2(n1733), .ZN(n1677) );
  INV_X1 U1152 ( .A(n1553), .ZN(n1552) );
  INV_X1 U1153 ( .A(n1549), .ZN(n1548) );
  INV_X1 U1154 ( .A(n1551), .ZN(n1550) );
  NAND3_X1 U1155 ( .A1(n1914), .A2(n1913), .A3(n1912), .ZN(n1864) );
  NAND3_X1 U1156 ( .A1(n1974), .A2(n1973), .A3(n1972), .ZN(n1924) );
  NAND2_X1 U1157 ( .A1(n2134), .A2(n2132), .ZN(n1976) );
  NAND2_X1 U1158 ( .A1(n1971), .A2(n1973), .ZN(n1917) );
  INV_X1 U1159 ( .A(n1541), .ZN(n1540) );
  INV_X1 U1160 ( .A(n1543), .ZN(n1542) );
  INV_X1 U1161 ( .A(n1545), .ZN(n1544) );
  INV_X1 U1162 ( .A(n1547), .ZN(n1546) );
  INV_X1 U1163 ( .A(n1555), .ZN(n1554) );
  OR2_X1 U1164 ( .A1(n2132), .A2(n2131), .ZN(n1535) );
  NAND2_X1 U1165 ( .A1(A[0]), .A2(n2111), .ZN(n1561) );
  INV_X2 U1166 ( .A(B[0]), .ZN(n1574) );
  INV_X1 U1167 ( .A(A[5]), .ZN(n1553) );
  INV_X1 U1168 ( .A(A[11]), .ZN(n1549) );
  INV_X1 U1169 ( .A(A[8]), .ZN(n1551) );
  INV_X1 U1170 ( .A(A[17]), .ZN(n1545) );
  INV_X1 U1171 ( .A(A[14]), .ZN(n1547) );
  INV_X1 U1172 ( .A(A[23]), .ZN(n1541) );
  INV_X1 U1173 ( .A(A[20]), .ZN(n1543) );
  NOR2_X4 U1174 ( .A1(n1670), .A2(n1671), .ZN(n1581) );
  NOR2_X4 U1175 ( .A1(n1672), .A2(n1673), .ZN(n1582) );
  NAND2_X2 U1176 ( .A1(n1670), .A2(n1672), .ZN(n1576) );
  NOR2_X4 U1177 ( .A1(n1731), .A2(n1732), .ZN(n1680) );
  NOR2_X4 U1178 ( .A1(n1733), .A2(n1734), .ZN(n1681) );
  NOR2_X4 U1179 ( .A1(n1791), .A2(n1792), .ZN(n1740) );
  NOR2_X4 U1180 ( .A1(n1793), .A2(n1794), .ZN(n1741) );
  NOR2_X4 U1181 ( .A1(n1851), .A2(n1852), .ZN(n1800) );
  NOR2_X4 U1182 ( .A1(n1853), .A2(n1854), .ZN(n1801) );
  NOR2_X4 U1183 ( .A1(n1911), .A2(n1912), .ZN(n1860) );
  NOR2_X4 U1184 ( .A1(n1913), .A2(n1914), .ZN(n1861) );
  NOR2_X4 U1185 ( .A1(n1971), .A2(n1972), .ZN(n1920) );
  NOR2_X4 U1186 ( .A1(n1973), .A2(n1974), .ZN(n1921) );
  NOR2_X4 U1187 ( .A1(n2112), .A2(n2111), .ZN(n1558) );
  NOR2_X4 U1188 ( .A1(n2113), .A2(A[0]), .ZN(n1559) );
  INV_X1 U1189 ( .A(B[23]), .ZN(n1555) );
  INV_X1 U1190 ( .A(B[23]), .ZN(n1556) );
  XNOR2_X1 U1191 ( .A(A[2]), .B(n1557), .ZN(n908) );
  AOI221_X1 U1192 ( .B1(B[22]), .B2(n1558), .C1(B[21]), .C2(n1559), .A(n1560), 
        .ZN(n1557) );
  OAI22_X1 U1193 ( .A1(n1561), .A2(n1562), .B1(n1563), .B2(n1564), .ZN(n1560)
         );
  XNOR2_X1 U1194 ( .A(A[2]), .B(n1565), .ZN(n907) );
  AOI221_X1 U1195 ( .B1(B[23]), .B2(n1558), .C1(n1559), .C2(B[22]), .A(n1566), 
        .ZN(n1565) );
  OAI22_X1 U1196 ( .A1(n1561), .A2(n1567), .B1(n1568), .B2(n1563), .ZN(n1566)
         );
  XNOR2_X1 U1197 ( .A(A[2]), .B(n1569), .ZN(n906) );
  AOI221_X1 U1198 ( .B1(B[23]), .B2(n1558), .C1(n1554), .C2(n1559), .A(n1570), 
        .ZN(n1569) );
  OAI22_X1 U1199 ( .A1(n1561), .A2(n1571), .B1(n1572), .B2(n1563), .ZN(n1570)
         );
  XNOR2_X1 U1200 ( .A(n1573), .B(n1553), .ZN(n904) );
  OAI22_X1 U1201 ( .A1(n1574), .A2(n1575), .B1(n1576), .B2(n1574), .ZN(n1573)
         );
  XNOR2_X1 U1202 ( .A(n1577), .B(n1553), .ZN(n903) );
  OAI222_X1 U1203 ( .A1(n1575), .A2(n1578), .B1(n1574), .B2(n1579), .C1(n1576), 
        .C2(n1580), .ZN(n1577) );
  INV_X1 U1204 ( .A(n1581), .ZN(n1579) );
  INV_X1 U1205 ( .A(n1582), .ZN(n1575) );
  XNOR2_X1 U1206 ( .A(n1552), .B(n1583), .ZN(n902) );
  AOI221_X1 U1207 ( .B1(B[2]), .B2(n1582), .C1(B[1]), .C2(n1581), .A(n1584), 
        .ZN(n1583) );
  OAI22_X1 U1208 ( .A1(n1576), .A2(n1585), .B1(n1574), .B2(n1586), .ZN(n1584)
         );
  XNOR2_X1 U1209 ( .A(n1552), .B(n1587), .ZN(n901) );
  AOI221_X1 U1210 ( .B1(B[3]), .B2(n1582), .C1(B[2]), .C2(n1581), .A(n1588), 
        .ZN(n1587) );
  OAI22_X1 U1211 ( .A1(n1576), .A2(n1589), .B1(n1578), .B2(n1586), .ZN(n1588)
         );
  XNOR2_X1 U1212 ( .A(n1552), .B(n1590), .ZN(n900) );
  AOI221_X1 U1213 ( .B1(B[4]), .B2(n1582), .C1(B[3]), .C2(n1581), .A(n1591), 
        .ZN(n1590) );
  OAI22_X1 U1214 ( .A1(n1576), .A2(n1592), .B1(n1593), .B2(n1586), .ZN(n1591)
         );
  XNOR2_X1 U1215 ( .A(n1552), .B(n1594), .ZN(n899) );
  AOI221_X1 U1216 ( .B1(B[5]), .B2(n1582), .C1(B[4]), .C2(n1581), .A(n1595), 
        .ZN(n1594) );
  OAI22_X1 U1217 ( .A1(n1576), .A2(n1596), .B1(n1586), .B2(n1597), .ZN(n1595)
         );
  XNOR2_X1 U1218 ( .A(n1552), .B(n1598), .ZN(n898) );
  AOI221_X1 U1219 ( .B1(B[6]), .B2(n1582), .C1(B[5]), .C2(n1581), .A(n1599), 
        .ZN(n1598) );
  OAI22_X1 U1220 ( .A1(n1576), .A2(n1600), .B1(n1586), .B2(n1601), .ZN(n1599)
         );
  XNOR2_X1 U1221 ( .A(n1552), .B(n1602), .ZN(n897) );
  AOI221_X1 U1222 ( .B1(B[7]), .B2(n1582), .C1(B[6]), .C2(n1581), .A(n1603), 
        .ZN(n1602) );
  OAI22_X1 U1223 ( .A1(n1576), .A2(n1604), .B1(n1586), .B2(n1605), .ZN(n1603)
         );
  XNOR2_X1 U1224 ( .A(n1552), .B(n1606), .ZN(n896) );
  AOI221_X1 U1225 ( .B1(B[8]), .B2(n1582), .C1(B[7]), .C2(n1581), .A(n1607), 
        .ZN(n1606) );
  OAI22_X1 U1226 ( .A1(n1576), .A2(n1608), .B1(n1586), .B2(n1609), .ZN(n1607)
         );
  XNOR2_X1 U1227 ( .A(n1552), .B(n1610), .ZN(n895) );
  AOI221_X1 U1228 ( .B1(B[9]), .B2(n1582), .C1(B[8]), .C2(n1581), .A(n1611), 
        .ZN(n1610) );
  OAI22_X1 U1229 ( .A1(n1576), .A2(n1612), .B1(n1586), .B2(n1613), .ZN(n1611)
         );
  XNOR2_X1 U1230 ( .A(n1552), .B(n1614), .ZN(n894) );
  AOI221_X1 U1231 ( .B1(B[10]), .B2(n1582), .C1(B[9]), .C2(n1581), .A(n1615), 
        .ZN(n1614) );
  OAI22_X1 U1232 ( .A1(n1576), .A2(n1616), .B1(n1586), .B2(n1617), .ZN(n1615)
         );
  XNOR2_X1 U1233 ( .A(n1552), .B(n1618), .ZN(n893) );
  AOI221_X1 U1234 ( .B1(B[11]), .B2(n1582), .C1(B[10]), .C2(n1581), .A(n1619), 
        .ZN(n1618) );
  OAI22_X1 U1235 ( .A1(n1576), .A2(n1620), .B1(n1586), .B2(n1621), .ZN(n1619)
         );
  XNOR2_X1 U1236 ( .A(n1552), .B(n1622), .ZN(n892) );
  AOI221_X1 U1237 ( .B1(B[12]), .B2(n1582), .C1(B[11]), .C2(n1581), .A(n1623), 
        .ZN(n1622) );
  OAI22_X1 U1238 ( .A1(n1576), .A2(n1624), .B1(n1586), .B2(n1625), .ZN(n1623)
         );
  XNOR2_X1 U1239 ( .A(n1552), .B(n1626), .ZN(n891) );
  AOI221_X1 U1240 ( .B1(B[13]), .B2(n1582), .C1(B[12]), .C2(n1581), .A(n1627), 
        .ZN(n1626) );
  OAI22_X1 U1241 ( .A1(n1576), .A2(n1628), .B1(n1586), .B2(n1629), .ZN(n1627)
         );
  XNOR2_X1 U1242 ( .A(n1552), .B(n1630), .ZN(n890) );
  AOI221_X1 U1243 ( .B1(B[14]), .B2(n1582), .C1(B[13]), .C2(n1581), .A(n1631), 
        .ZN(n1630) );
  OAI22_X1 U1244 ( .A1(n1576), .A2(n1632), .B1(n1586), .B2(n1633), .ZN(n1631)
         );
  XNOR2_X1 U1245 ( .A(n1552), .B(n1634), .ZN(n889) );
  AOI221_X1 U1246 ( .B1(B[15]), .B2(n1582), .C1(B[14]), .C2(n1581), .A(n1635), 
        .ZN(n1634) );
  OAI22_X1 U1247 ( .A1(n1576), .A2(n1636), .B1(n1586), .B2(n1637), .ZN(n1635)
         );
  XNOR2_X1 U1248 ( .A(n1552), .B(n1638), .ZN(n888) );
  AOI221_X1 U1249 ( .B1(B[16]), .B2(n1582), .C1(B[15]), .C2(n1581), .A(n1639), 
        .ZN(n1638) );
  OAI22_X1 U1250 ( .A1(n1576), .A2(n1640), .B1(n1586), .B2(n1641), .ZN(n1639)
         );
  XNOR2_X1 U1251 ( .A(n1552), .B(n1642), .ZN(n887) );
  AOI221_X1 U1252 ( .B1(B[17]), .B2(n1582), .C1(B[16]), .C2(n1581), .A(n1643), 
        .ZN(n1642) );
  OAI22_X1 U1253 ( .A1(n1576), .A2(n1644), .B1(n1586), .B2(n1645), .ZN(n1643)
         );
  XNOR2_X1 U1254 ( .A(n1552), .B(n1646), .ZN(n886) );
  AOI221_X1 U1255 ( .B1(B[18]), .B2(n1582), .C1(B[17]), .C2(n1581), .A(n1647), 
        .ZN(n1646) );
  OAI22_X1 U1256 ( .A1(n1576), .A2(n1648), .B1(n1586), .B2(n1649), .ZN(n1647)
         );
  XNOR2_X1 U1257 ( .A(n1552), .B(n1650), .ZN(n885) );
  AOI221_X1 U1258 ( .B1(B[19]), .B2(n1582), .C1(B[18]), .C2(n1581), .A(n1651), 
        .ZN(n1650) );
  OAI22_X1 U1259 ( .A1(n1576), .A2(n1652), .B1(n1586), .B2(n1653), .ZN(n1651)
         );
  XNOR2_X1 U1260 ( .A(A[5]), .B(n1654), .ZN(n884) );
  AOI221_X1 U1261 ( .B1(n1582), .B2(B[20]), .C1(B[19]), .C2(n1581), .A(n1655), 
        .ZN(n1654) );
  OAI22_X1 U1262 ( .A1(n1576), .A2(n1656), .B1(n1586), .B2(n1657), .ZN(n1655)
         );
  XNOR2_X1 U1263 ( .A(A[5]), .B(n1658), .ZN(n883) );
  AOI221_X1 U1264 ( .B1(n1582), .B2(B[21]), .C1(n1581), .C2(B[20]), .A(n1659), 
        .ZN(n1658) );
  OAI22_X1 U1265 ( .A1(n1576), .A2(n1660), .B1(n1586), .B2(n1661), .ZN(n1659)
         );
  XNOR2_X1 U1266 ( .A(A[5]), .B(n1662), .ZN(n882) );
  AOI221_X1 U1267 ( .B1(n1582), .B2(B[22]), .C1(n1581), .C2(B[21]), .A(n1663), 
        .ZN(n1662) );
  OAI22_X1 U1268 ( .A1(n1562), .A2(n1576), .B1(n1564), .B2(n1586), .ZN(n1663)
         );
  XNOR2_X1 U1269 ( .A(A[5]), .B(n1664), .ZN(n881) );
  AOI221_X1 U1270 ( .B1(n1582), .B2(B[23]), .C1(n1581), .C2(B[22]), .A(n1665), 
        .ZN(n1664) );
  OAI22_X1 U1271 ( .A1(n1567), .A2(n1576), .B1(n1568), .B2(n1586), .ZN(n1665)
         );
  XNOR2_X1 U1272 ( .A(A[5]), .B(n1666), .ZN(n880) );
  AOI221_X1 U1273 ( .B1(n1582), .B2(B[23]), .C1(n1581), .C2(n1554), .A(n1667), 
        .ZN(n1666) );
  OAI22_X1 U1274 ( .A1(n1571), .A2(n1576), .B1(n1572), .B2(n1586), .ZN(n1667)
         );
  XNOR2_X1 U1275 ( .A(n1552), .B(n1668), .ZN(n879) );
  OAI221_X1 U1276 ( .B1(n1556), .B2(n1586), .C1(n1556), .C2(n1576), .A(n1669), 
        .ZN(n1668) );
  OAI21_X1 U1277 ( .B1(n1582), .B2(n1581), .A(n1554), .ZN(n1669) );
  INV_X1 U1278 ( .A(n1673), .ZN(n1670) );
  XNOR2_X1 U1279 ( .A(A[3]), .B(A[4]), .ZN(n1671) );
  XNOR2_X1 U1280 ( .A(A[4]), .B(n1553), .ZN(n1672) );
  XOR2_X1 U1281 ( .A(A[3]), .B(n1674), .Z(n1673) );
  XNOR2_X1 U1282 ( .A(n1675), .B(n1551), .ZN(n878) );
  OAI22_X1 U1283 ( .A1(n1574), .A2(n1676), .B1(n1574), .B2(n1677), .ZN(n1675)
         );
  XNOR2_X1 U1284 ( .A(n1678), .B(n1551), .ZN(n877) );
  OAI222_X1 U1285 ( .A1(n1578), .A2(n1676), .B1(n1574), .B2(n1679), .C1(n1580), 
        .C2(n1677), .ZN(n1678) );
  INV_X1 U1286 ( .A(n1680), .ZN(n1679) );
  INV_X1 U1287 ( .A(n1681), .ZN(n1676) );
  XNOR2_X1 U1288 ( .A(n1550), .B(n1682), .ZN(n876) );
  AOI221_X1 U1289 ( .B1(n1681), .B2(B[2]), .C1(n1680), .C2(B[1]), .A(n1683), 
        .ZN(n1682) );
  OAI22_X1 U1290 ( .A1(n1585), .A2(n1677), .B1(n1574), .B2(n1684), .ZN(n1683)
         );
  XNOR2_X1 U1291 ( .A(n1550), .B(n1685), .ZN(n875) );
  AOI221_X1 U1292 ( .B1(n1681), .B2(B[3]), .C1(n1680), .C2(B[2]), .A(n1686), 
        .ZN(n1685) );
  OAI22_X1 U1293 ( .A1(n1589), .A2(n1677), .B1(n1578), .B2(n1684), .ZN(n1686)
         );
  XNOR2_X1 U1294 ( .A(n1550), .B(n1687), .ZN(n874) );
  AOI221_X1 U1295 ( .B1(n1681), .B2(B[4]), .C1(n1680), .C2(B[3]), .A(n1688), 
        .ZN(n1687) );
  OAI22_X1 U1296 ( .A1(n1592), .A2(n1677), .B1(n1593), .B2(n1684), .ZN(n1688)
         );
  XNOR2_X1 U1297 ( .A(n1550), .B(n1689), .ZN(n873) );
  AOI221_X1 U1298 ( .B1(n1681), .B2(B[5]), .C1(n1680), .C2(B[4]), .A(n1690), 
        .ZN(n1689) );
  OAI22_X1 U1299 ( .A1(n1596), .A2(n1677), .B1(n1597), .B2(n1684), .ZN(n1690)
         );
  XNOR2_X1 U1300 ( .A(n1550), .B(n1691), .ZN(n872) );
  AOI221_X1 U1301 ( .B1(n1681), .B2(B[6]), .C1(n1680), .C2(B[5]), .A(n1692), 
        .ZN(n1691) );
  OAI22_X1 U1302 ( .A1(n1600), .A2(n1677), .B1(n1601), .B2(n1684), .ZN(n1692)
         );
  XNOR2_X1 U1303 ( .A(n1550), .B(n1693), .ZN(n871) );
  AOI221_X1 U1304 ( .B1(n1681), .B2(B[7]), .C1(n1680), .C2(B[6]), .A(n1694), 
        .ZN(n1693) );
  OAI22_X1 U1305 ( .A1(n1604), .A2(n1677), .B1(n1605), .B2(n1684), .ZN(n1694)
         );
  XNOR2_X1 U1306 ( .A(n1550), .B(n1695), .ZN(n870) );
  AOI221_X1 U1307 ( .B1(n1681), .B2(B[8]), .C1(n1680), .C2(B[7]), .A(n1696), 
        .ZN(n1695) );
  OAI22_X1 U1308 ( .A1(n1608), .A2(n1677), .B1(n1609), .B2(n1684), .ZN(n1696)
         );
  XNOR2_X1 U1309 ( .A(n1550), .B(n1697), .ZN(n869) );
  AOI221_X1 U1310 ( .B1(n1681), .B2(B[9]), .C1(n1680), .C2(B[8]), .A(n1698), 
        .ZN(n1697) );
  OAI22_X1 U1311 ( .A1(n1612), .A2(n1677), .B1(n1613), .B2(n1684), .ZN(n1698)
         );
  XNOR2_X1 U1312 ( .A(n1550), .B(n1699), .ZN(n868) );
  AOI221_X1 U1313 ( .B1(n1681), .B2(B[10]), .C1(n1680), .C2(B[9]), .A(n1700), 
        .ZN(n1699) );
  OAI22_X1 U1314 ( .A1(n1616), .A2(n1677), .B1(n1617), .B2(n1684), .ZN(n1700)
         );
  XNOR2_X1 U1315 ( .A(n1550), .B(n1701), .ZN(n867) );
  AOI221_X1 U1316 ( .B1(n1681), .B2(B[11]), .C1(n1680), .C2(B[10]), .A(n1702), 
        .ZN(n1701) );
  OAI22_X1 U1317 ( .A1(n1620), .A2(n1677), .B1(n1621), .B2(n1684), .ZN(n1702)
         );
  XNOR2_X1 U1318 ( .A(n1550), .B(n1703), .ZN(n866) );
  AOI221_X1 U1319 ( .B1(n1681), .B2(B[12]), .C1(n1680), .C2(B[11]), .A(n1704), 
        .ZN(n1703) );
  OAI22_X1 U1320 ( .A1(n1624), .A2(n1677), .B1(n1625), .B2(n1684), .ZN(n1704)
         );
  XNOR2_X1 U1321 ( .A(n1550), .B(n1705), .ZN(n865) );
  AOI221_X1 U1322 ( .B1(n1681), .B2(B[13]), .C1(n1680), .C2(B[12]), .A(n1706), 
        .ZN(n1705) );
  OAI22_X1 U1323 ( .A1(n1628), .A2(n1677), .B1(n1629), .B2(n1684), .ZN(n1706)
         );
  XNOR2_X1 U1324 ( .A(n1550), .B(n1707), .ZN(n864) );
  AOI221_X1 U1325 ( .B1(n1681), .B2(B[14]), .C1(n1680), .C2(B[13]), .A(n1708), 
        .ZN(n1707) );
  OAI22_X1 U1326 ( .A1(n1632), .A2(n1677), .B1(n1633), .B2(n1684), .ZN(n1708)
         );
  XNOR2_X1 U1327 ( .A(n1550), .B(n1709), .ZN(n863) );
  AOI221_X1 U1328 ( .B1(n1681), .B2(B[15]), .C1(n1680), .C2(B[14]), .A(n1710), 
        .ZN(n1709) );
  OAI22_X1 U1329 ( .A1(n1636), .A2(n1677), .B1(n1637), .B2(n1684), .ZN(n1710)
         );
  XNOR2_X1 U1330 ( .A(n1550), .B(n1711), .ZN(n862) );
  AOI221_X1 U1331 ( .B1(n1681), .B2(B[16]), .C1(n1680), .C2(B[15]), .A(n1712), 
        .ZN(n1711) );
  OAI22_X1 U1332 ( .A1(n1640), .A2(n1677), .B1(n1641), .B2(n1684), .ZN(n1712)
         );
  XNOR2_X1 U1333 ( .A(n1550), .B(n1713), .ZN(n861) );
  AOI221_X1 U1334 ( .B1(n1681), .B2(B[17]), .C1(n1680), .C2(B[16]), .A(n1714), 
        .ZN(n1713) );
  OAI22_X1 U1335 ( .A1(n1644), .A2(n1677), .B1(n1645), .B2(n1684), .ZN(n1714)
         );
  XNOR2_X1 U1336 ( .A(n1550), .B(n1715), .ZN(n860) );
  AOI221_X1 U1337 ( .B1(n1681), .B2(B[18]), .C1(n1680), .C2(B[17]), .A(n1716), 
        .ZN(n1715) );
  OAI22_X1 U1338 ( .A1(n1648), .A2(n1677), .B1(n1649), .B2(n1684), .ZN(n1716)
         );
  XNOR2_X1 U1339 ( .A(n1550), .B(n1717), .ZN(n859) );
  AOI221_X1 U1340 ( .B1(n1681), .B2(B[19]), .C1(n1680), .C2(B[18]), .A(n1718), 
        .ZN(n1717) );
  OAI22_X1 U1341 ( .A1(n1652), .A2(n1677), .B1(n1653), .B2(n1684), .ZN(n1718)
         );
  XNOR2_X1 U1342 ( .A(A[8]), .B(n1719), .ZN(n858) );
  AOI221_X1 U1343 ( .B1(n1681), .B2(B[20]), .C1(n1680), .C2(B[19]), .A(n1720), 
        .ZN(n1719) );
  OAI22_X1 U1344 ( .A1(n1656), .A2(n1677), .B1(n1657), .B2(n1684), .ZN(n1720)
         );
  XNOR2_X1 U1345 ( .A(A[8]), .B(n1721), .ZN(n857) );
  AOI221_X1 U1346 ( .B1(n1681), .B2(B[21]), .C1(n1680), .C2(B[20]), .A(n1722), 
        .ZN(n1721) );
  OAI22_X1 U1347 ( .A1(n1660), .A2(n1677), .B1(n1661), .B2(n1684), .ZN(n1722)
         );
  XNOR2_X1 U1348 ( .A(A[8]), .B(n1723), .ZN(n856) );
  AOI221_X1 U1349 ( .B1(n1681), .B2(B[22]), .C1(n1680), .C2(B[21]), .A(n1724), 
        .ZN(n1723) );
  OAI22_X1 U1350 ( .A1(n1562), .A2(n1677), .B1(n1564), .B2(n1684), .ZN(n1724)
         );
  XNOR2_X1 U1351 ( .A(A[8]), .B(n1725), .ZN(n855) );
  AOI221_X1 U1352 ( .B1(n1681), .B2(B[23]), .C1(n1680), .C2(B[22]), .A(n1726), 
        .ZN(n1725) );
  OAI22_X1 U1353 ( .A1(n1567), .A2(n1677), .B1(n1568), .B2(n1684), .ZN(n1726)
         );
  XNOR2_X1 U1354 ( .A(A[8]), .B(n1727), .ZN(n854) );
  AOI221_X1 U1355 ( .B1(n1681), .B2(B[23]), .C1(n1680), .C2(n1554), .A(n1728), 
        .ZN(n1727) );
  OAI22_X1 U1356 ( .A1(n1571), .A2(n1677), .B1(n1572), .B2(n1684), .ZN(n1728)
         );
  XNOR2_X1 U1357 ( .A(n1550), .B(n1729), .ZN(n853) );
  OAI221_X1 U1358 ( .B1(n1555), .B2(n1684), .C1(n1556), .C2(n1677), .A(n1730), 
        .ZN(n1729) );
  OAI21_X1 U1359 ( .B1(n1681), .B2(n1680), .A(n1554), .ZN(n1730) );
  INV_X1 U1360 ( .A(n1734), .ZN(n1731) );
  XNOR2_X1 U1361 ( .A(A[6]), .B(A[7]), .ZN(n1732) );
  XNOR2_X1 U1362 ( .A(A[7]), .B(n1551), .ZN(n1733) );
  XOR2_X1 U1363 ( .A(A[6]), .B(n1553), .Z(n1734) );
  XNOR2_X1 U1364 ( .A(n1735), .B(n1549), .ZN(n852) );
  OAI22_X1 U1365 ( .A1(n1574), .A2(n1736), .B1(n1574), .B2(n1737), .ZN(n1735)
         );
  XNOR2_X1 U1366 ( .A(n1738), .B(n1549), .ZN(n851) );
  OAI222_X1 U1367 ( .A1(n1578), .A2(n1736), .B1(n1574), .B2(n1739), .C1(n1580), 
        .C2(n1737), .ZN(n1738) );
  INV_X1 U1368 ( .A(n1740), .ZN(n1739) );
  INV_X1 U1369 ( .A(n1741), .ZN(n1736) );
  XNOR2_X1 U1370 ( .A(n1548), .B(n1742), .ZN(n850) );
  AOI221_X1 U1371 ( .B1(n1741), .B2(B[2]), .C1(n1740), .C2(B[1]), .A(n1743), 
        .ZN(n1742) );
  OAI22_X1 U1372 ( .A1(n1585), .A2(n1737), .B1(n1574), .B2(n1744), .ZN(n1743)
         );
  XNOR2_X1 U1373 ( .A(n1548), .B(n1745), .ZN(n849) );
  AOI221_X1 U1374 ( .B1(n1741), .B2(B[3]), .C1(n1740), .C2(B[2]), .A(n1746), 
        .ZN(n1745) );
  OAI22_X1 U1375 ( .A1(n1589), .A2(n1737), .B1(n1578), .B2(n1744), .ZN(n1746)
         );
  XNOR2_X1 U1376 ( .A(n1548), .B(n1747), .ZN(n848) );
  AOI221_X1 U1377 ( .B1(n1741), .B2(B[4]), .C1(n1740), .C2(B[3]), .A(n1748), 
        .ZN(n1747) );
  OAI22_X1 U1378 ( .A1(n1592), .A2(n1737), .B1(n1593), .B2(n1744), .ZN(n1748)
         );
  XNOR2_X1 U1379 ( .A(n1548), .B(n1749), .ZN(n847) );
  AOI221_X1 U1380 ( .B1(n1741), .B2(B[5]), .C1(n1740), .C2(B[4]), .A(n1750), 
        .ZN(n1749) );
  OAI22_X1 U1381 ( .A1(n1596), .A2(n1737), .B1(n1597), .B2(n1744), .ZN(n1750)
         );
  XNOR2_X1 U1382 ( .A(n1548), .B(n1751), .ZN(n846) );
  AOI221_X1 U1383 ( .B1(n1741), .B2(B[6]), .C1(n1740), .C2(B[5]), .A(n1752), 
        .ZN(n1751) );
  OAI22_X1 U1384 ( .A1(n1600), .A2(n1737), .B1(n1601), .B2(n1744), .ZN(n1752)
         );
  XNOR2_X1 U1385 ( .A(n1548), .B(n1753), .ZN(n845) );
  AOI221_X1 U1386 ( .B1(n1741), .B2(B[7]), .C1(n1740), .C2(B[6]), .A(n1754), 
        .ZN(n1753) );
  OAI22_X1 U1387 ( .A1(n1604), .A2(n1737), .B1(n1605), .B2(n1744), .ZN(n1754)
         );
  XNOR2_X1 U1388 ( .A(n1548), .B(n1755), .ZN(n844) );
  AOI221_X1 U1389 ( .B1(n1741), .B2(B[8]), .C1(n1740), .C2(B[7]), .A(n1756), 
        .ZN(n1755) );
  OAI22_X1 U1390 ( .A1(n1608), .A2(n1737), .B1(n1609), .B2(n1744), .ZN(n1756)
         );
  XNOR2_X1 U1391 ( .A(n1548), .B(n1757), .ZN(n843) );
  AOI221_X1 U1392 ( .B1(n1741), .B2(B[9]), .C1(n1740), .C2(B[8]), .A(n1758), 
        .ZN(n1757) );
  OAI22_X1 U1393 ( .A1(n1612), .A2(n1737), .B1(n1613), .B2(n1744), .ZN(n1758)
         );
  XNOR2_X1 U1394 ( .A(n1548), .B(n1759), .ZN(n842) );
  AOI221_X1 U1395 ( .B1(n1741), .B2(B[10]), .C1(n1740), .C2(B[9]), .A(n1760), 
        .ZN(n1759) );
  OAI22_X1 U1396 ( .A1(n1616), .A2(n1737), .B1(n1617), .B2(n1744), .ZN(n1760)
         );
  XNOR2_X1 U1397 ( .A(n1548), .B(n1761), .ZN(n841) );
  AOI221_X1 U1398 ( .B1(n1741), .B2(B[11]), .C1(n1740), .C2(B[10]), .A(n1762), 
        .ZN(n1761) );
  OAI22_X1 U1399 ( .A1(n1620), .A2(n1737), .B1(n1621), .B2(n1744), .ZN(n1762)
         );
  XNOR2_X1 U1400 ( .A(n1548), .B(n1763), .ZN(n840) );
  AOI221_X1 U1401 ( .B1(n1741), .B2(B[12]), .C1(n1740), .C2(B[11]), .A(n1764), 
        .ZN(n1763) );
  OAI22_X1 U1402 ( .A1(n1624), .A2(n1737), .B1(n1625), .B2(n1744), .ZN(n1764)
         );
  XNOR2_X1 U1403 ( .A(n1548), .B(n1765), .ZN(n839) );
  AOI221_X1 U1404 ( .B1(n1741), .B2(B[13]), .C1(n1740), .C2(B[12]), .A(n1766), 
        .ZN(n1765) );
  OAI22_X1 U1405 ( .A1(n1628), .A2(n1737), .B1(n1629), .B2(n1744), .ZN(n1766)
         );
  XNOR2_X1 U1406 ( .A(n1548), .B(n1767), .ZN(n838) );
  AOI221_X1 U1407 ( .B1(n1741), .B2(B[14]), .C1(n1740), .C2(B[13]), .A(n1768), 
        .ZN(n1767) );
  OAI22_X1 U1408 ( .A1(n1632), .A2(n1737), .B1(n1633), .B2(n1744), .ZN(n1768)
         );
  XNOR2_X1 U1409 ( .A(n1548), .B(n1769), .ZN(n837) );
  AOI221_X1 U1410 ( .B1(n1741), .B2(B[15]), .C1(n1740), .C2(B[14]), .A(n1770), 
        .ZN(n1769) );
  OAI22_X1 U1411 ( .A1(n1636), .A2(n1737), .B1(n1637), .B2(n1744), .ZN(n1770)
         );
  XNOR2_X1 U1412 ( .A(n1548), .B(n1771), .ZN(n836) );
  AOI221_X1 U1413 ( .B1(n1741), .B2(B[16]), .C1(n1740), .C2(B[15]), .A(n1772), 
        .ZN(n1771) );
  OAI22_X1 U1414 ( .A1(n1640), .A2(n1737), .B1(n1641), .B2(n1744), .ZN(n1772)
         );
  XNOR2_X1 U1415 ( .A(n1548), .B(n1773), .ZN(n835) );
  AOI221_X1 U1416 ( .B1(n1741), .B2(B[17]), .C1(n1740), .C2(B[16]), .A(n1774), 
        .ZN(n1773) );
  OAI22_X1 U1417 ( .A1(n1644), .A2(n1737), .B1(n1645), .B2(n1744), .ZN(n1774)
         );
  XNOR2_X1 U1418 ( .A(n1548), .B(n1775), .ZN(n834) );
  AOI221_X1 U1419 ( .B1(n1741), .B2(B[18]), .C1(n1740), .C2(B[17]), .A(n1776), 
        .ZN(n1775) );
  OAI22_X1 U1420 ( .A1(n1648), .A2(n1737), .B1(n1649), .B2(n1744), .ZN(n1776)
         );
  XNOR2_X1 U1421 ( .A(n1548), .B(n1777), .ZN(n833) );
  AOI221_X1 U1422 ( .B1(n1741), .B2(B[19]), .C1(n1740), .C2(B[18]), .A(n1778), 
        .ZN(n1777) );
  OAI22_X1 U1423 ( .A1(n1652), .A2(n1737), .B1(n1653), .B2(n1744), .ZN(n1778)
         );
  XNOR2_X1 U1424 ( .A(n1548), .B(n1779), .ZN(n832) );
  AOI221_X1 U1425 ( .B1(n1741), .B2(B[20]), .C1(n1740), .C2(B[19]), .A(n1780), 
        .ZN(n1779) );
  OAI22_X1 U1426 ( .A1(n1656), .A2(n1737), .B1(n1657), .B2(n1744), .ZN(n1780)
         );
  XNOR2_X1 U1427 ( .A(A[11]), .B(n1781), .ZN(n831) );
  AOI221_X1 U1428 ( .B1(n1741), .B2(B[21]), .C1(n1740), .C2(B[20]), .A(n1782), 
        .ZN(n1781) );
  OAI22_X1 U1429 ( .A1(n1660), .A2(n1737), .B1(n1661), .B2(n1744), .ZN(n1782)
         );
  XNOR2_X1 U1430 ( .A(A[11]), .B(n1783), .ZN(n830) );
  AOI221_X1 U1431 ( .B1(n1741), .B2(B[22]), .C1(n1740), .C2(B[21]), .A(n1784), 
        .ZN(n1783) );
  OAI22_X1 U1432 ( .A1(n1562), .A2(n1737), .B1(n1564), .B2(n1744), .ZN(n1784)
         );
  XNOR2_X1 U1433 ( .A(A[11]), .B(n1785), .ZN(n829) );
  AOI221_X1 U1434 ( .B1(n1741), .B2(B[23]), .C1(n1740), .C2(B[22]), .A(n1786), 
        .ZN(n1785) );
  OAI22_X1 U1435 ( .A1(n1567), .A2(n1737), .B1(n1568), .B2(n1744), .ZN(n1786)
         );
  XNOR2_X1 U1436 ( .A(A[11]), .B(n1787), .ZN(n828) );
  AOI221_X1 U1437 ( .B1(n1741), .B2(B[23]), .C1(n1740), .C2(n1554), .A(n1788), 
        .ZN(n1787) );
  OAI22_X1 U1438 ( .A1(n1571), .A2(n1737), .B1(n1572), .B2(n1744), .ZN(n1788)
         );
  XNOR2_X1 U1439 ( .A(A[11]), .B(n1789), .ZN(n827) );
  OAI221_X1 U1440 ( .B1(n1556), .B2(n1744), .C1(n1556), .C2(n1737), .A(n1790), 
        .ZN(n1789) );
  OAI21_X1 U1441 ( .B1(n1741), .B2(n1740), .A(n1554), .ZN(n1790) );
  INV_X1 U1442 ( .A(n1794), .ZN(n1791) );
  XNOR2_X1 U1443 ( .A(A[10]), .B(A[9]), .ZN(n1792) );
  XNOR2_X1 U1444 ( .A(A[10]), .B(n1549), .ZN(n1793) );
  XOR2_X1 U1445 ( .A(A[9]), .B(n1551), .Z(n1794) );
  XNOR2_X1 U1446 ( .A(n1795), .B(n1547), .ZN(n826) );
  OAI22_X1 U1447 ( .A1(n1574), .A2(n1796), .B1(n1574), .B2(n1797), .ZN(n1795)
         );
  XNOR2_X1 U1448 ( .A(n1798), .B(n1547), .ZN(n825) );
  OAI222_X1 U1449 ( .A1(n1578), .A2(n1796), .B1(n1574), .B2(n1799), .C1(n1580), 
        .C2(n1797), .ZN(n1798) );
  INV_X1 U1450 ( .A(n1800), .ZN(n1799) );
  INV_X1 U1451 ( .A(n1801), .ZN(n1796) );
  XNOR2_X1 U1452 ( .A(n1546), .B(n1802), .ZN(n824) );
  AOI221_X1 U1453 ( .B1(n1801), .B2(B[2]), .C1(n1800), .C2(B[1]), .A(n1803), 
        .ZN(n1802) );
  OAI22_X1 U1454 ( .A1(n1585), .A2(n1797), .B1(n1574), .B2(n1804), .ZN(n1803)
         );
  XNOR2_X1 U1455 ( .A(n1546), .B(n1805), .ZN(n823) );
  AOI221_X1 U1456 ( .B1(n1801), .B2(B[3]), .C1(n1800), .C2(B[2]), .A(n1806), 
        .ZN(n1805) );
  OAI22_X1 U1457 ( .A1(n1589), .A2(n1797), .B1(n1578), .B2(n1804), .ZN(n1806)
         );
  XNOR2_X1 U1458 ( .A(n1546), .B(n1807), .ZN(n822) );
  AOI221_X1 U1459 ( .B1(n1801), .B2(B[4]), .C1(n1800), .C2(B[3]), .A(n1808), 
        .ZN(n1807) );
  OAI22_X1 U1460 ( .A1(n1592), .A2(n1797), .B1(n1593), .B2(n1804), .ZN(n1808)
         );
  XNOR2_X1 U1461 ( .A(n1546), .B(n1809), .ZN(n821) );
  AOI221_X1 U1462 ( .B1(n1801), .B2(B[5]), .C1(n1800), .C2(B[4]), .A(n1810), 
        .ZN(n1809) );
  OAI22_X1 U1463 ( .A1(n1596), .A2(n1797), .B1(n1597), .B2(n1804), .ZN(n1810)
         );
  XNOR2_X1 U1464 ( .A(n1546), .B(n1811), .ZN(n820) );
  AOI221_X1 U1465 ( .B1(n1801), .B2(B[6]), .C1(n1800), .C2(B[5]), .A(n1812), 
        .ZN(n1811) );
  OAI22_X1 U1466 ( .A1(n1600), .A2(n1797), .B1(n1601), .B2(n1804), .ZN(n1812)
         );
  XNOR2_X1 U1467 ( .A(n1546), .B(n1813), .ZN(n819) );
  AOI221_X1 U1468 ( .B1(n1801), .B2(B[7]), .C1(n1800), .C2(B[6]), .A(n1814), 
        .ZN(n1813) );
  OAI22_X1 U1469 ( .A1(n1604), .A2(n1797), .B1(n1605), .B2(n1804), .ZN(n1814)
         );
  XNOR2_X1 U1470 ( .A(n1546), .B(n1815), .ZN(n818) );
  AOI221_X1 U1471 ( .B1(n1801), .B2(B[8]), .C1(n1800), .C2(B[7]), .A(n1816), 
        .ZN(n1815) );
  OAI22_X1 U1472 ( .A1(n1608), .A2(n1797), .B1(n1609), .B2(n1804), .ZN(n1816)
         );
  XNOR2_X1 U1473 ( .A(n1546), .B(n1817), .ZN(n817) );
  AOI221_X1 U1474 ( .B1(n1801), .B2(B[9]), .C1(n1800), .C2(B[8]), .A(n1818), 
        .ZN(n1817) );
  OAI22_X1 U1475 ( .A1(n1612), .A2(n1797), .B1(n1613), .B2(n1804), .ZN(n1818)
         );
  XNOR2_X1 U1476 ( .A(n1546), .B(n1819), .ZN(n816) );
  AOI221_X1 U1477 ( .B1(n1801), .B2(B[10]), .C1(n1800), .C2(B[9]), .A(n1820), 
        .ZN(n1819) );
  OAI22_X1 U1478 ( .A1(n1616), .A2(n1797), .B1(n1617), .B2(n1804), .ZN(n1820)
         );
  XNOR2_X1 U1479 ( .A(n1546), .B(n1821), .ZN(n815) );
  AOI221_X1 U1480 ( .B1(n1801), .B2(B[11]), .C1(n1800), .C2(B[10]), .A(n1822), 
        .ZN(n1821) );
  OAI22_X1 U1481 ( .A1(n1620), .A2(n1797), .B1(n1621), .B2(n1804), .ZN(n1822)
         );
  XNOR2_X1 U1482 ( .A(n1546), .B(n1823), .ZN(n814) );
  AOI221_X1 U1483 ( .B1(n1801), .B2(B[12]), .C1(n1800), .C2(B[11]), .A(n1824), 
        .ZN(n1823) );
  OAI22_X1 U1484 ( .A1(n1624), .A2(n1797), .B1(n1625), .B2(n1804), .ZN(n1824)
         );
  XNOR2_X1 U1485 ( .A(n1546), .B(n1825), .ZN(n813) );
  AOI221_X1 U1486 ( .B1(n1801), .B2(B[13]), .C1(n1800), .C2(B[12]), .A(n1826), 
        .ZN(n1825) );
  OAI22_X1 U1487 ( .A1(n1628), .A2(n1797), .B1(n1629), .B2(n1804), .ZN(n1826)
         );
  XNOR2_X1 U1488 ( .A(n1546), .B(n1827), .ZN(n812) );
  AOI221_X1 U1489 ( .B1(n1801), .B2(B[14]), .C1(n1800), .C2(B[13]), .A(n1828), 
        .ZN(n1827) );
  OAI22_X1 U1490 ( .A1(n1632), .A2(n1797), .B1(n1633), .B2(n1804), .ZN(n1828)
         );
  XNOR2_X1 U1491 ( .A(n1546), .B(n1829), .ZN(n811) );
  AOI221_X1 U1492 ( .B1(n1801), .B2(B[15]), .C1(n1800), .C2(B[14]), .A(n1830), 
        .ZN(n1829) );
  OAI22_X1 U1493 ( .A1(n1636), .A2(n1797), .B1(n1637), .B2(n1804), .ZN(n1830)
         );
  XNOR2_X1 U1494 ( .A(n1546), .B(n1831), .ZN(n810) );
  AOI221_X1 U1495 ( .B1(n1801), .B2(B[16]), .C1(n1800), .C2(B[15]), .A(n1832), 
        .ZN(n1831) );
  OAI22_X1 U1496 ( .A1(n1640), .A2(n1797), .B1(n1641), .B2(n1804), .ZN(n1832)
         );
  XNOR2_X1 U1497 ( .A(n1546), .B(n1833), .ZN(n809) );
  AOI221_X1 U1498 ( .B1(n1801), .B2(B[17]), .C1(n1800), .C2(B[16]), .A(n1834), 
        .ZN(n1833) );
  OAI22_X1 U1499 ( .A1(n1644), .A2(n1797), .B1(n1645), .B2(n1804), .ZN(n1834)
         );
  XNOR2_X1 U1500 ( .A(n1546), .B(n1835), .ZN(n808) );
  AOI221_X1 U1501 ( .B1(n1801), .B2(B[18]), .C1(n1800), .C2(B[17]), .A(n1836), 
        .ZN(n1835) );
  OAI22_X1 U1502 ( .A1(n1648), .A2(n1797), .B1(n1649), .B2(n1804), .ZN(n1836)
         );
  XNOR2_X1 U1503 ( .A(n1546), .B(n1837), .ZN(n807) );
  AOI221_X1 U1504 ( .B1(n1801), .B2(B[19]), .C1(n1800), .C2(B[18]), .A(n1838), 
        .ZN(n1837) );
  OAI22_X1 U1505 ( .A1(n1652), .A2(n1797), .B1(n1653), .B2(n1804), .ZN(n1838)
         );
  XNOR2_X1 U1506 ( .A(n1546), .B(n1839), .ZN(n806) );
  AOI221_X1 U1507 ( .B1(n1801), .B2(B[20]), .C1(n1800), .C2(B[19]), .A(n1840), 
        .ZN(n1839) );
  OAI22_X1 U1508 ( .A1(n1656), .A2(n1797), .B1(n1657), .B2(n1804), .ZN(n1840)
         );
  XNOR2_X1 U1509 ( .A(A[14]), .B(n1841), .ZN(n805) );
  AOI221_X1 U1510 ( .B1(n1801), .B2(B[21]), .C1(n1800), .C2(B[20]), .A(n1842), 
        .ZN(n1841) );
  OAI22_X1 U1511 ( .A1(n1660), .A2(n1797), .B1(n1661), .B2(n1804), .ZN(n1842)
         );
  XNOR2_X1 U1512 ( .A(A[14]), .B(n1843), .ZN(n804) );
  AOI221_X1 U1513 ( .B1(n1801), .B2(B[22]), .C1(n1800), .C2(B[21]), .A(n1844), 
        .ZN(n1843) );
  OAI22_X1 U1514 ( .A1(n1562), .A2(n1797), .B1(n1564), .B2(n1804), .ZN(n1844)
         );
  XNOR2_X1 U1515 ( .A(A[14]), .B(n1845), .ZN(n803) );
  AOI221_X1 U1516 ( .B1(n1801), .B2(B[23]), .C1(n1800), .C2(B[22]), .A(n1846), 
        .ZN(n1845) );
  OAI22_X1 U1517 ( .A1(n1567), .A2(n1797), .B1(n1568), .B2(n1804), .ZN(n1846)
         );
  XNOR2_X1 U1518 ( .A(A[14]), .B(n1847), .ZN(n802) );
  AOI221_X1 U1519 ( .B1(n1801), .B2(B[23]), .C1(n1800), .C2(n1554), .A(n1848), 
        .ZN(n1847) );
  OAI22_X1 U1520 ( .A1(n1571), .A2(n1797), .B1(n1572), .B2(n1804), .ZN(n1848)
         );
  XNOR2_X1 U1521 ( .A(A[14]), .B(n1849), .ZN(n801) );
  OAI221_X1 U1522 ( .B1(n1556), .B2(n1804), .C1(n1556), .C2(n1797), .A(n1850), 
        .ZN(n1849) );
  OAI21_X1 U1523 ( .B1(n1801), .B2(n1800), .A(n1554), .ZN(n1850) );
  INV_X1 U1524 ( .A(n1854), .ZN(n1851) );
  XNOR2_X1 U1525 ( .A(A[12]), .B(A[13]), .ZN(n1852) );
  XNOR2_X1 U1526 ( .A(A[13]), .B(n1547), .ZN(n1853) );
  XOR2_X1 U1527 ( .A(A[12]), .B(n1549), .Z(n1854) );
  XNOR2_X1 U1528 ( .A(n1855), .B(n1545), .ZN(n800) );
  OAI22_X1 U1529 ( .A1(n1574), .A2(n1856), .B1(n1574), .B2(n1857), .ZN(n1855)
         );
  XNOR2_X1 U1530 ( .A(n1858), .B(n1545), .ZN(n799) );
  OAI222_X1 U1531 ( .A1(n1578), .A2(n1856), .B1(n1574), .B2(n1859), .C1(n1580), 
        .C2(n1857), .ZN(n1858) );
  INV_X1 U1532 ( .A(n1860), .ZN(n1859) );
  INV_X1 U1533 ( .A(n1861), .ZN(n1856) );
  XNOR2_X1 U1534 ( .A(n1544), .B(n1862), .ZN(n798) );
  AOI221_X1 U1535 ( .B1(n1861), .B2(B[2]), .C1(n1860), .C2(B[1]), .A(n1863), 
        .ZN(n1862) );
  OAI22_X1 U1536 ( .A1(n1585), .A2(n1857), .B1(n1574), .B2(n1864), .ZN(n1863)
         );
  XNOR2_X1 U1537 ( .A(n1544), .B(n1865), .ZN(n797) );
  AOI221_X1 U1538 ( .B1(n1861), .B2(B[3]), .C1(n1860), .C2(B[2]), .A(n1866), 
        .ZN(n1865) );
  OAI22_X1 U1539 ( .A1(n1589), .A2(n1857), .B1(n1578), .B2(n1864), .ZN(n1866)
         );
  XNOR2_X1 U1540 ( .A(n1544), .B(n1867), .ZN(n796) );
  AOI221_X1 U1541 ( .B1(n1861), .B2(B[4]), .C1(n1860), .C2(B[3]), .A(n1868), 
        .ZN(n1867) );
  OAI22_X1 U1542 ( .A1(n1592), .A2(n1857), .B1(n1593), .B2(n1864), .ZN(n1868)
         );
  XNOR2_X1 U1543 ( .A(n1544), .B(n1869), .ZN(n795) );
  AOI221_X1 U1544 ( .B1(n1861), .B2(B[5]), .C1(n1860), .C2(B[4]), .A(n1870), 
        .ZN(n1869) );
  OAI22_X1 U1545 ( .A1(n1596), .A2(n1857), .B1(n1597), .B2(n1864), .ZN(n1870)
         );
  XNOR2_X1 U1546 ( .A(n1544), .B(n1871), .ZN(n794) );
  AOI221_X1 U1547 ( .B1(n1861), .B2(B[6]), .C1(n1860), .C2(B[5]), .A(n1872), 
        .ZN(n1871) );
  OAI22_X1 U1548 ( .A1(n1600), .A2(n1857), .B1(n1601), .B2(n1864), .ZN(n1872)
         );
  XNOR2_X1 U1549 ( .A(n1544), .B(n1873), .ZN(n793) );
  AOI221_X1 U1550 ( .B1(n1861), .B2(B[7]), .C1(n1860), .C2(B[6]), .A(n1874), 
        .ZN(n1873) );
  OAI22_X1 U1551 ( .A1(n1604), .A2(n1857), .B1(n1605), .B2(n1864), .ZN(n1874)
         );
  XNOR2_X1 U1552 ( .A(n1544), .B(n1875), .ZN(n792) );
  AOI221_X1 U1553 ( .B1(n1861), .B2(B[8]), .C1(n1860), .C2(B[7]), .A(n1876), 
        .ZN(n1875) );
  OAI22_X1 U1554 ( .A1(n1608), .A2(n1857), .B1(n1609), .B2(n1864), .ZN(n1876)
         );
  XNOR2_X1 U1555 ( .A(n1544), .B(n1877), .ZN(n791) );
  AOI221_X1 U1556 ( .B1(n1861), .B2(B[9]), .C1(n1860), .C2(B[8]), .A(n1878), 
        .ZN(n1877) );
  OAI22_X1 U1557 ( .A1(n1612), .A2(n1857), .B1(n1613), .B2(n1864), .ZN(n1878)
         );
  XNOR2_X1 U1558 ( .A(n1544), .B(n1879), .ZN(n790) );
  AOI221_X1 U1559 ( .B1(n1861), .B2(B[10]), .C1(n1860), .C2(B[9]), .A(n1880), 
        .ZN(n1879) );
  OAI22_X1 U1560 ( .A1(n1616), .A2(n1857), .B1(n1617), .B2(n1864), .ZN(n1880)
         );
  XNOR2_X1 U1561 ( .A(n1544), .B(n1881), .ZN(n789) );
  AOI221_X1 U1562 ( .B1(n1861), .B2(B[11]), .C1(n1860), .C2(B[10]), .A(n1882), 
        .ZN(n1881) );
  OAI22_X1 U1563 ( .A1(n1620), .A2(n1857), .B1(n1621), .B2(n1864), .ZN(n1882)
         );
  XNOR2_X1 U1564 ( .A(n1544), .B(n1883), .ZN(n788) );
  AOI221_X1 U1565 ( .B1(n1861), .B2(B[12]), .C1(n1860), .C2(B[11]), .A(n1884), 
        .ZN(n1883) );
  OAI22_X1 U1566 ( .A1(n1624), .A2(n1857), .B1(n1625), .B2(n1864), .ZN(n1884)
         );
  XNOR2_X1 U1567 ( .A(n1544), .B(n1885), .ZN(n787) );
  AOI221_X1 U1568 ( .B1(n1861), .B2(B[13]), .C1(n1860), .C2(B[12]), .A(n1886), 
        .ZN(n1885) );
  OAI22_X1 U1569 ( .A1(n1628), .A2(n1857), .B1(n1629), .B2(n1864), .ZN(n1886)
         );
  XNOR2_X1 U1570 ( .A(n1544), .B(n1887), .ZN(n786) );
  AOI221_X1 U1571 ( .B1(n1861), .B2(B[14]), .C1(n1860), .C2(B[13]), .A(n1888), 
        .ZN(n1887) );
  OAI22_X1 U1572 ( .A1(n1632), .A2(n1857), .B1(n1633), .B2(n1864), .ZN(n1888)
         );
  XNOR2_X1 U1573 ( .A(n1544), .B(n1889), .ZN(n785) );
  AOI221_X1 U1574 ( .B1(n1861), .B2(B[15]), .C1(n1860), .C2(B[14]), .A(n1890), 
        .ZN(n1889) );
  OAI22_X1 U1575 ( .A1(n1636), .A2(n1857), .B1(n1637), .B2(n1864), .ZN(n1890)
         );
  XNOR2_X1 U1576 ( .A(n1544), .B(n1891), .ZN(n784) );
  AOI221_X1 U1577 ( .B1(n1861), .B2(B[16]), .C1(n1860), .C2(B[15]), .A(n1892), 
        .ZN(n1891) );
  OAI22_X1 U1578 ( .A1(n1640), .A2(n1857), .B1(n1641), .B2(n1864), .ZN(n1892)
         );
  XNOR2_X1 U1579 ( .A(n1544), .B(n1893), .ZN(n783) );
  AOI221_X1 U1580 ( .B1(n1861), .B2(B[17]), .C1(n1860), .C2(B[16]), .A(n1894), 
        .ZN(n1893) );
  OAI22_X1 U1581 ( .A1(n1644), .A2(n1857), .B1(n1645), .B2(n1864), .ZN(n1894)
         );
  XNOR2_X1 U1582 ( .A(n1544), .B(n1895), .ZN(n782) );
  AOI221_X1 U1583 ( .B1(n1861), .B2(B[18]), .C1(n1860), .C2(B[17]), .A(n1896), 
        .ZN(n1895) );
  OAI22_X1 U1584 ( .A1(n1648), .A2(n1857), .B1(n1649), .B2(n1864), .ZN(n1896)
         );
  XNOR2_X1 U1585 ( .A(n1544), .B(n1897), .ZN(n781) );
  AOI221_X1 U1586 ( .B1(n1861), .B2(B[19]), .C1(n1860), .C2(B[18]), .A(n1898), 
        .ZN(n1897) );
  OAI22_X1 U1587 ( .A1(n1652), .A2(n1857), .B1(n1653), .B2(n1864), .ZN(n1898)
         );
  XNOR2_X1 U1588 ( .A(n1544), .B(n1899), .ZN(n780) );
  AOI221_X1 U1589 ( .B1(n1861), .B2(B[20]), .C1(n1860), .C2(B[19]), .A(n1900), 
        .ZN(n1899) );
  OAI22_X1 U1590 ( .A1(n1656), .A2(n1857), .B1(n1657), .B2(n1864), .ZN(n1900)
         );
  XNOR2_X1 U1591 ( .A(A[17]), .B(n1901), .ZN(n779) );
  AOI221_X1 U1592 ( .B1(n1861), .B2(B[21]), .C1(n1860), .C2(B[20]), .A(n1902), 
        .ZN(n1901) );
  OAI22_X1 U1593 ( .A1(n1660), .A2(n1857), .B1(n1661), .B2(n1864), .ZN(n1902)
         );
  XNOR2_X1 U1594 ( .A(A[17]), .B(n1903), .ZN(n778) );
  AOI221_X1 U1595 ( .B1(n1861), .B2(B[22]), .C1(n1860), .C2(B[21]), .A(n1904), 
        .ZN(n1903) );
  OAI22_X1 U1596 ( .A1(n1562), .A2(n1857), .B1(n1564), .B2(n1864), .ZN(n1904)
         );
  XNOR2_X1 U1597 ( .A(A[17]), .B(n1905), .ZN(n777) );
  AOI221_X1 U1598 ( .B1(n1861), .B2(B[23]), .C1(n1860), .C2(B[22]), .A(n1906), 
        .ZN(n1905) );
  OAI22_X1 U1599 ( .A1(n1567), .A2(n1857), .B1(n1568), .B2(n1864), .ZN(n1906)
         );
  XNOR2_X1 U1600 ( .A(A[17]), .B(n1907), .ZN(n776) );
  AOI221_X1 U1601 ( .B1(n1861), .B2(B[23]), .C1(n1860), .C2(n1554), .A(n1908), 
        .ZN(n1907) );
  OAI22_X1 U1602 ( .A1(n1571), .A2(n1857), .B1(n1572), .B2(n1864), .ZN(n1908)
         );
  XNOR2_X1 U1603 ( .A(A[17]), .B(n1909), .ZN(n775) );
  OAI221_X1 U1604 ( .B1(n1556), .B2(n1864), .C1(n1556), .C2(n1857), .A(n1910), 
        .ZN(n1909) );
  OAI21_X1 U1605 ( .B1(n1861), .B2(n1860), .A(n1554), .ZN(n1910) );
  INV_X1 U1606 ( .A(n1914), .ZN(n1911) );
  XNOR2_X1 U1607 ( .A(A[15]), .B(A[16]), .ZN(n1912) );
  XNOR2_X1 U1608 ( .A(A[16]), .B(n1545), .ZN(n1913) );
  XOR2_X1 U1609 ( .A(A[15]), .B(n1547), .Z(n1914) );
  XNOR2_X1 U1610 ( .A(n1915), .B(n1543), .ZN(n774) );
  OAI22_X1 U1611 ( .A1(n1574), .A2(n1916), .B1(n1574), .B2(n1917), .ZN(n1915)
         );
  XNOR2_X1 U1612 ( .A(n1918), .B(n1543), .ZN(n773) );
  OAI222_X1 U1613 ( .A1(n1578), .A2(n1916), .B1(n1574), .B2(n1919), .C1(n1580), 
        .C2(n1917), .ZN(n1918) );
  INV_X1 U1614 ( .A(n1920), .ZN(n1919) );
  INV_X1 U1615 ( .A(n1921), .ZN(n1916) );
  XNOR2_X1 U1616 ( .A(n1542), .B(n1922), .ZN(n772) );
  AOI221_X1 U1617 ( .B1(n1921), .B2(B[2]), .C1(n1920), .C2(B[1]), .A(n1923), 
        .ZN(n1922) );
  OAI22_X1 U1618 ( .A1(n1585), .A2(n1917), .B1(n1574), .B2(n1924), .ZN(n1923)
         );
  XNOR2_X1 U1619 ( .A(n1542), .B(n1925), .ZN(n771) );
  AOI221_X1 U1620 ( .B1(n1921), .B2(B[3]), .C1(n1920), .C2(B[2]), .A(n1926), 
        .ZN(n1925) );
  OAI22_X1 U1621 ( .A1(n1589), .A2(n1917), .B1(n1578), .B2(n1924), .ZN(n1926)
         );
  XNOR2_X1 U1622 ( .A(n1542), .B(n1927), .ZN(n770) );
  AOI221_X1 U1623 ( .B1(n1921), .B2(B[4]), .C1(n1920), .C2(B[3]), .A(n1928), 
        .ZN(n1927) );
  OAI22_X1 U1624 ( .A1(n1592), .A2(n1917), .B1(n1593), .B2(n1924), .ZN(n1928)
         );
  XNOR2_X1 U1625 ( .A(n1542), .B(n1929), .ZN(n769) );
  AOI221_X1 U1626 ( .B1(n1921), .B2(B[5]), .C1(n1920), .C2(B[4]), .A(n1930), 
        .ZN(n1929) );
  OAI22_X1 U1627 ( .A1(n1596), .A2(n1917), .B1(n1597), .B2(n1924), .ZN(n1930)
         );
  XNOR2_X1 U1628 ( .A(n1542), .B(n1931), .ZN(n768) );
  AOI221_X1 U1629 ( .B1(n1921), .B2(B[6]), .C1(n1920), .C2(B[5]), .A(n1932), 
        .ZN(n1931) );
  OAI22_X1 U1630 ( .A1(n1600), .A2(n1917), .B1(n1601), .B2(n1924), .ZN(n1932)
         );
  XNOR2_X1 U1631 ( .A(n1542), .B(n1933), .ZN(n767) );
  AOI221_X1 U1632 ( .B1(n1921), .B2(B[7]), .C1(n1920), .C2(B[6]), .A(n1934), 
        .ZN(n1933) );
  OAI22_X1 U1633 ( .A1(n1604), .A2(n1917), .B1(n1605), .B2(n1924), .ZN(n1934)
         );
  XNOR2_X1 U1634 ( .A(n1542), .B(n1935), .ZN(n766) );
  AOI221_X1 U1635 ( .B1(n1921), .B2(B[8]), .C1(n1920), .C2(B[7]), .A(n1936), 
        .ZN(n1935) );
  OAI22_X1 U1636 ( .A1(n1608), .A2(n1917), .B1(n1609), .B2(n1924), .ZN(n1936)
         );
  XNOR2_X1 U1637 ( .A(n1542), .B(n1937), .ZN(n765) );
  AOI221_X1 U1638 ( .B1(n1921), .B2(B[9]), .C1(n1920), .C2(B[8]), .A(n1938), 
        .ZN(n1937) );
  OAI22_X1 U1639 ( .A1(n1612), .A2(n1917), .B1(n1613), .B2(n1924), .ZN(n1938)
         );
  XNOR2_X1 U1640 ( .A(n1542), .B(n1939), .ZN(n764) );
  AOI221_X1 U1641 ( .B1(n1921), .B2(B[10]), .C1(n1920), .C2(B[9]), .A(n1940), 
        .ZN(n1939) );
  OAI22_X1 U1642 ( .A1(n1616), .A2(n1917), .B1(n1617), .B2(n1924), .ZN(n1940)
         );
  XNOR2_X1 U1643 ( .A(n1542), .B(n1941), .ZN(n763) );
  AOI221_X1 U1644 ( .B1(n1921), .B2(B[11]), .C1(n1920), .C2(B[10]), .A(n1942), 
        .ZN(n1941) );
  OAI22_X1 U1645 ( .A1(n1620), .A2(n1917), .B1(n1621), .B2(n1924), .ZN(n1942)
         );
  XNOR2_X1 U1646 ( .A(n1542), .B(n1943), .ZN(n762) );
  AOI221_X1 U1647 ( .B1(n1921), .B2(B[12]), .C1(n1920), .C2(B[11]), .A(n1944), 
        .ZN(n1943) );
  OAI22_X1 U1648 ( .A1(n1624), .A2(n1917), .B1(n1625), .B2(n1924), .ZN(n1944)
         );
  XNOR2_X1 U1649 ( .A(n1542), .B(n1945), .ZN(n761) );
  AOI221_X1 U1650 ( .B1(n1921), .B2(B[13]), .C1(n1920), .C2(B[12]), .A(n1946), 
        .ZN(n1945) );
  OAI22_X1 U1651 ( .A1(n1628), .A2(n1917), .B1(n1629), .B2(n1924), .ZN(n1946)
         );
  XNOR2_X1 U1652 ( .A(n1542), .B(n1947), .ZN(n760) );
  AOI221_X1 U1653 ( .B1(n1921), .B2(B[14]), .C1(n1920), .C2(B[13]), .A(n1948), 
        .ZN(n1947) );
  OAI22_X1 U1654 ( .A1(n1632), .A2(n1917), .B1(n1633), .B2(n1924), .ZN(n1948)
         );
  XNOR2_X1 U1655 ( .A(n1542), .B(n1949), .ZN(n759) );
  AOI221_X1 U1656 ( .B1(n1921), .B2(B[15]), .C1(n1920), .C2(B[14]), .A(n1950), 
        .ZN(n1949) );
  OAI22_X1 U1657 ( .A1(n1636), .A2(n1917), .B1(n1637), .B2(n1924), .ZN(n1950)
         );
  XNOR2_X1 U1658 ( .A(n1542), .B(n1951), .ZN(n758) );
  AOI221_X1 U1659 ( .B1(n1921), .B2(B[16]), .C1(n1920), .C2(B[15]), .A(n1952), 
        .ZN(n1951) );
  OAI22_X1 U1660 ( .A1(n1640), .A2(n1917), .B1(n1641), .B2(n1924), .ZN(n1952)
         );
  XNOR2_X1 U1661 ( .A(n1542), .B(n1953), .ZN(n757) );
  AOI221_X1 U1662 ( .B1(n1921), .B2(B[17]), .C1(n1920), .C2(B[16]), .A(n1954), 
        .ZN(n1953) );
  OAI22_X1 U1663 ( .A1(n1644), .A2(n1917), .B1(n1645), .B2(n1924), .ZN(n1954)
         );
  XNOR2_X1 U1664 ( .A(n1542), .B(n1955), .ZN(n756) );
  AOI221_X1 U1665 ( .B1(n1921), .B2(B[18]), .C1(n1920), .C2(B[17]), .A(n1956), 
        .ZN(n1955) );
  OAI22_X1 U1666 ( .A1(n1648), .A2(n1917), .B1(n1649), .B2(n1924), .ZN(n1956)
         );
  XNOR2_X1 U1667 ( .A(n1542), .B(n1957), .ZN(n755) );
  AOI221_X1 U1668 ( .B1(n1921), .B2(B[19]), .C1(n1920), .C2(B[18]), .A(n1958), 
        .ZN(n1957) );
  OAI22_X1 U1669 ( .A1(n1652), .A2(n1917), .B1(n1653), .B2(n1924), .ZN(n1958)
         );
  XNOR2_X1 U1670 ( .A(n1542), .B(n1959), .ZN(n754) );
  AOI221_X1 U1671 ( .B1(n1921), .B2(B[20]), .C1(n1920), .C2(B[19]), .A(n1960), 
        .ZN(n1959) );
  OAI22_X1 U1672 ( .A1(n1656), .A2(n1917), .B1(n1657), .B2(n1924), .ZN(n1960)
         );
  XNOR2_X1 U1673 ( .A(A[20]), .B(n1961), .ZN(n753) );
  AOI221_X1 U1674 ( .B1(n1921), .B2(B[21]), .C1(n1920), .C2(B[20]), .A(n1962), 
        .ZN(n1961) );
  OAI22_X1 U1675 ( .A1(n1660), .A2(n1917), .B1(n1661), .B2(n1924), .ZN(n1962)
         );
  XNOR2_X1 U1676 ( .A(A[20]), .B(n1963), .ZN(n752) );
  AOI221_X1 U1677 ( .B1(n1921), .B2(B[22]), .C1(n1920), .C2(B[21]), .A(n1964), 
        .ZN(n1963) );
  OAI22_X1 U1678 ( .A1(n1562), .A2(n1917), .B1(n1564), .B2(n1924), .ZN(n1964)
         );
  XNOR2_X1 U1679 ( .A(A[20]), .B(n1965), .ZN(n751) );
  AOI221_X1 U1680 ( .B1(n1921), .B2(n1554), .C1(n1920), .C2(B[22]), .A(n1966), 
        .ZN(n1965) );
  OAI22_X1 U1681 ( .A1(n1567), .A2(n1917), .B1(n1568), .B2(n1924), .ZN(n1966)
         );
  XNOR2_X1 U1682 ( .A(A[20]), .B(n1967), .ZN(n750) );
  AOI221_X1 U1683 ( .B1(n1921), .B2(B[23]), .C1(n1920), .C2(n1554), .A(n1968), 
        .ZN(n1967) );
  OAI22_X1 U1684 ( .A1(n1571), .A2(n1917), .B1(n1572), .B2(n1924), .ZN(n1968)
         );
  XNOR2_X1 U1685 ( .A(A[20]), .B(n1969), .ZN(n749) );
  OAI221_X1 U1686 ( .B1(n1556), .B2(n1924), .C1(n1556), .C2(n1917), .A(n1970), 
        .ZN(n1969) );
  OAI21_X1 U1687 ( .B1(n1921), .B2(n1920), .A(n1554), .ZN(n1970) );
  INV_X1 U1688 ( .A(n1974), .ZN(n1971) );
  XNOR2_X1 U1689 ( .A(A[18]), .B(A[19]), .ZN(n1972) );
  XNOR2_X1 U1690 ( .A(A[19]), .B(n1543), .ZN(n1973) );
  XOR2_X1 U1691 ( .A(A[18]), .B(n1545), .Z(n1974) );
  XNOR2_X1 U1692 ( .A(n1975), .B(n1541), .ZN(n748) );
  OAI22_X1 U1693 ( .A1(n1574), .A2(n1535), .B1(n1574), .B2(n1976), .ZN(n1975)
         );
  XNOR2_X1 U1694 ( .A(n1977), .B(n1541), .ZN(n747) );
  OAI222_X1 U1695 ( .A1(n1578), .A2(n1535), .B1(n1574), .B2(n1534), .C1(n1580), 
        .C2(n1976), .ZN(n1977) );
  INV_X1 U1696 ( .A(n1397), .ZN(n1580) );
  XNOR2_X1 U1697 ( .A(n1540), .B(n1978), .ZN(n746) );
  AOI221_X1 U1698 ( .B1(n1537), .B2(B[2]), .C1(n1536), .C2(B[1]), .A(n1979), 
        .ZN(n1978) );
  OAI22_X1 U1699 ( .A1(n1585), .A2(n1976), .B1(n1574), .B2(n1538), .ZN(n1979)
         );
  INV_X1 U1700 ( .A(n1396), .ZN(n1585) );
  XNOR2_X1 U1701 ( .A(n1540), .B(n1981), .ZN(n745) );
  AOI221_X1 U1702 ( .B1(n1537), .B2(B[3]), .C1(n1536), .C2(B[2]), .A(n1982), 
        .ZN(n1981) );
  OAI22_X1 U1703 ( .A1(n1589), .A2(n1976), .B1(n1578), .B2(n1539), .ZN(n1982)
         );
  XNOR2_X1 U1704 ( .A(n1540), .B(n1983), .ZN(n744) );
  AOI221_X1 U1705 ( .B1(n1537), .B2(B[4]), .C1(n1536), .C2(B[3]), .A(n1984), 
        .ZN(n1983) );
  OAI22_X1 U1706 ( .A1(n1592), .A2(n1976), .B1(n1593), .B2(n1539), .ZN(n1984)
         );
  XNOR2_X1 U1707 ( .A(n1540), .B(n1985), .ZN(n743) );
  AOI221_X1 U1708 ( .B1(n1537), .B2(B[5]), .C1(n1536), .C2(B[4]), .A(n1986), 
        .ZN(n1985) );
  OAI22_X1 U1709 ( .A1(n1596), .A2(n1976), .B1(n1597), .B2(n1539), .ZN(n1986)
         );
  XNOR2_X1 U1710 ( .A(n1540), .B(n1987), .ZN(n742) );
  AOI221_X1 U1711 ( .B1(n1537), .B2(B[6]), .C1(n1536), .C2(B[5]), .A(n1988), 
        .ZN(n1987) );
  OAI22_X1 U1712 ( .A1(n1600), .A2(n1976), .B1(n1601), .B2(n1539), .ZN(n1988)
         );
  XNOR2_X1 U1713 ( .A(n1540), .B(n1989), .ZN(n741) );
  AOI221_X1 U1714 ( .B1(n1537), .B2(B[7]), .C1(n1536), .C2(B[6]), .A(n1990), 
        .ZN(n1989) );
  OAI22_X1 U1715 ( .A1(n1604), .A2(n1976), .B1(n1605), .B2(n1539), .ZN(n1990)
         );
  XNOR2_X1 U1716 ( .A(n1540), .B(n1991), .ZN(n740) );
  AOI221_X1 U1717 ( .B1(n1537), .B2(B[9]), .C1(n1536), .C2(B[8]), .A(n1992), 
        .ZN(n1991) );
  OAI22_X1 U1718 ( .A1(n1612), .A2(n1976), .B1(n1613), .B2(n1539), .ZN(n1992)
         );
  XNOR2_X1 U1719 ( .A(n1540), .B(n1993), .ZN(n739) );
  AOI221_X1 U1720 ( .B1(n1537), .B2(B[10]), .C1(n1536), .C2(B[9]), .A(n1994), 
        .ZN(n1993) );
  OAI22_X1 U1721 ( .A1(n1616), .A2(n1976), .B1(n1617), .B2(n1539), .ZN(n1994)
         );
  XNOR2_X1 U1722 ( .A(n1540), .B(n1995), .ZN(n738) );
  AOI221_X1 U1723 ( .B1(n1537), .B2(B[12]), .C1(n1536), .C2(B[11]), .A(n1996), 
        .ZN(n1995) );
  OAI22_X1 U1724 ( .A1(n1624), .A2(n1976), .B1(n1625), .B2(n1539), .ZN(n1996)
         );
  XNOR2_X1 U1725 ( .A(n1540), .B(n1997), .ZN(n737) );
  AOI221_X1 U1726 ( .B1(n1537), .B2(B[13]), .C1(n1536), .C2(B[12]), .A(n1998), 
        .ZN(n1997) );
  OAI22_X1 U1727 ( .A1(n1628), .A2(n1976), .B1(n1629), .B2(n1539), .ZN(n1998)
         );
  XNOR2_X1 U1728 ( .A(n1540), .B(n1999), .ZN(n736) );
  AOI221_X1 U1729 ( .B1(n1537), .B2(B[14]), .C1(n1536), .C2(B[13]), .A(n2000), 
        .ZN(n1999) );
  OAI22_X1 U1730 ( .A1(n1632), .A2(n1976), .B1(n1633), .B2(n1539), .ZN(n2000)
         );
  XNOR2_X1 U1731 ( .A(n1540), .B(n2001), .ZN(n735) );
  AOI221_X1 U1732 ( .B1(n1537), .B2(B[15]), .C1(n1536), .C2(B[14]), .A(n2002), 
        .ZN(n2001) );
  OAI22_X1 U1733 ( .A1(n1636), .A2(n1976), .B1(n1637), .B2(n1539), .ZN(n2002)
         );
  XNOR2_X1 U1734 ( .A(n1540), .B(n2003), .ZN(n734) );
  AOI221_X1 U1735 ( .B1(n1537), .B2(B[16]), .C1(n1536), .C2(B[15]), .A(n2004), 
        .ZN(n2003) );
  OAI22_X1 U1736 ( .A1(n1640), .A2(n1976), .B1(n1641), .B2(n1538), .ZN(n2004)
         );
  XNOR2_X1 U1737 ( .A(n1540), .B(n2005), .ZN(n733) );
  AOI221_X1 U1738 ( .B1(n1537), .B2(B[18]), .C1(n1536), .C2(B[17]), .A(n2006), 
        .ZN(n2005) );
  OAI22_X1 U1739 ( .A1(n1648), .A2(n1976), .B1(n1649), .B2(n1538), .ZN(n2006)
         );
  XNOR2_X1 U1740 ( .A(n1540), .B(n2007), .ZN(n732) );
  AOI221_X1 U1741 ( .B1(n1537), .B2(B[19]), .C1(n1536), .C2(B[18]), .A(n2008), 
        .ZN(n2007) );
  OAI22_X1 U1742 ( .A1(n1652), .A2(n1976), .B1(n1653), .B2(n1538), .ZN(n2008)
         );
  XNOR2_X1 U1743 ( .A(n1540), .B(n2009), .ZN(n731) );
  AOI221_X1 U1744 ( .B1(n1537), .B2(B[20]), .C1(n1536), .C2(B[19]), .A(n2010), 
        .ZN(n2009) );
  OAI22_X1 U1745 ( .A1(n1656), .A2(n1976), .B1(n1657), .B2(n1538), .ZN(n2010)
         );
  XNOR2_X1 U1746 ( .A(A[23]), .B(n2011), .ZN(n730) );
  AOI221_X1 U1747 ( .B1(n1537), .B2(B[21]), .C1(n1536), .C2(B[20]), .A(n2012), 
        .ZN(n2011) );
  OAI22_X1 U1748 ( .A1(n1660), .A2(n1976), .B1(n1661), .B2(n1538), .ZN(n2012)
         );
  XNOR2_X1 U1749 ( .A(A[23]), .B(n2013), .ZN(n729) );
  AOI221_X1 U1750 ( .B1(n1537), .B2(B[22]), .C1(n1536), .C2(B[21]), .A(n2014), 
        .ZN(n2013) );
  OAI22_X1 U1751 ( .A1(n1562), .A2(n1976), .B1(n1564), .B2(n1538), .ZN(n2014)
         );
  INV_X1 U1752 ( .A(B[20]), .ZN(n1564) );
  INV_X1 U1753 ( .A(n1376), .ZN(n1562) );
  XNOR2_X1 U1754 ( .A(n519), .B(n2015), .ZN(n506) );
  INV_X1 U1755 ( .A(n493), .ZN(n479) );
  NOR2_X1 U1756 ( .A1(n2015), .A2(n519), .ZN(n493) );
  XOR2_X1 U1757 ( .A(n2016), .B(n1674), .Z(n2015) );
  OAI221_X1 U1758 ( .B1(n1563), .B2(n1556), .C1(n1561), .C2(n1556), .A(n2017), 
        .ZN(n2016) );
  OAI21_X1 U1759 ( .B1(n1558), .B2(n1559), .A(n1554), .ZN(n2017) );
  INV_X1 U1760 ( .A(n454), .ZN(n442) );
  XOR2_X1 U1761 ( .A(n1540), .B(n2018), .Z(n454) );
  AOI221_X1 U1762 ( .B1(n1537), .B2(B[8]), .C1(n1536), .C2(B[7]), .A(n2019), 
        .ZN(n2018) );
  OAI22_X1 U1763 ( .A1(n1608), .A2(n1976), .B1(n1609), .B2(n1538), .ZN(n2019)
         );
  INV_X1 U1764 ( .A(n421), .ZN(n411) );
  XOR2_X1 U1765 ( .A(n1540), .B(n2020), .Z(n421) );
  AOI221_X1 U1766 ( .B1(n1537), .B2(B[11]), .C1(n1536), .C2(B[10]), .A(n2021), 
        .ZN(n2020) );
  OAI22_X1 U1767 ( .A1(n1620), .A2(n1976), .B1(n1621), .B2(n1538), .ZN(n2021)
         );
  INV_X1 U1768 ( .A(n387), .ZN(n395) );
  INV_X1 U1769 ( .A(n374), .ZN(n368) );
  XOR2_X1 U1770 ( .A(n1540), .B(n2022), .Z(n374) );
  AOI221_X1 U1771 ( .B1(n1537), .B2(B[17]), .C1(n1536), .C2(B[16]), .A(n2023), 
        .ZN(n2022) );
  OAI22_X1 U1772 ( .A1(n1644), .A2(n1976), .B1(n1645), .B2(n1538), .ZN(n2023)
         );
  INV_X1 U1773 ( .A(n356), .ZN(n360) );
  INV_X1 U1774 ( .A(n2024), .ZN(n351) );
  OAI222_X1 U1775 ( .A1(n2025), .A2(n2026), .B1(n2025), .B2(n2027), .C1(n2027), 
        .C2(n2026), .ZN(n326) );
  INV_X1 U1776 ( .A(n550), .ZN(n2027) );
  XNOR2_X1 U1777 ( .A(n1674), .B(n2028), .ZN(n2026) );
  AOI221_X1 U1778 ( .B1(B[21]), .B2(n1558), .C1(B[20]), .C2(n1559), .A(n2029), 
        .ZN(n2028) );
  OAI22_X1 U1779 ( .A1(n1561), .A2(n1660), .B1(n1563), .B2(n1661), .ZN(n2029)
         );
  INV_X1 U1780 ( .A(B[19]), .ZN(n1661) );
  INV_X1 U1781 ( .A(n1377), .ZN(n1660) );
  AOI222_X1 U1782 ( .A1(n2030), .A2(n2031), .B1(n2030), .B2(n564), .C1(n564), 
        .C2(n2031), .ZN(n2025) );
  XNOR2_X1 U1783 ( .A(A[2]), .B(n2032), .ZN(n2031) );
  AOI221_X1 U1784 ( .B1(B[20]), .B2(n1558), .C1(B[19]), .C2(n1559), .A(n2033), 
        .ZN(n2032) );
  OAI22_X1 U1785 ( .A1(n1561), .A2(n1656), .B1(n1563), .B2(n1657), .ZN(n2033)
         );
  INV_X1 U1786 ( .A(B[18]), .ZN(n1657) );
  INV_X1 U1787 ( .A(n1378), .ZN(n1656) );
  INV_X1 U1788 ( .A(n2034), .ZN(n2030) );
  AOI222_X1 U1789 ( .A1(n2035), .A2(n2036), .B1(n2035), .B2(n576), .C1(n576), 
        .C2(n2036), .ZN(n2034) );
  XNOR2_X1 U1790 ( .A(A[2]), .B(n2037), .ZN(n2036) );
  AOI221_X1 U1791 ( .B1(B[19]), .B2(n1558), .C1(B[18]), .C2(n1559), .A(n2038), 
        .ZN(n2037) );
  OAI22_X1 U1792 ( .A1(n1561), .A2(n1652), .B1(n1563), .B2(n1653), .ZN(n2038)
         );
  INV_X1 U1793 ( .A(B[17]), .ZN(n1653) );
  INV_X1 U1794 ( .A(n1379), .ZN(n1652) );
  OAI222_X1 U1795 ( .A1(n2039), .A2(n2040), .B1(n2039), .B2(n2041), .C1(n2041), 
        .C2(n2040), .ZN(n2035) );
  INV_X1 U1796 ( .A(n588), .ZN(n2041) );
  XNOR2_X1 U1797 ( .A(n1674), .B(n2042), .ZN(n2040) );
  AOI221_X1 U1798 ( .B1(B[18]), .B2(n1558), .C1(B[17]), .C2(n1559), .A(n2043), 
        .ZN(n2042) );
  OAI22_X1 U1799 ( .A1(n1561), .A2(n1648), .B1(n1563), .B2(n1649), .ZN(n2043)
         );
  INV_X1 U1800 ( .A(B[16]), .ZN(n1649) );
  INV_X1 U1801 ( .A(n1380), .ZN(n1648) );
  AOI222_X1 U1802 ( .A1(n2044), .A2(n2045), .B1(n2044), .B2(n600), .C1(n600), 
        .C2(n2045), .ZN(n2039) );
  XNOR2_X1 U1803 ( .A(A[2]), .B(n2046), .ZN(n2045) );
  AOI221_X1 U1804 ( .B1(B[17]), .B2(n1558), .C1(B[16]), .C2(n1559), .A(n2047), 
        .ZN(n2046) );
  OAI22_X1 U1805 ( .A1(n1561), .A2(n1644), .B1(n1563), .B2(n1645), .ZN(n2047)
         );
  INV_X1 U1806 ( .A(B[15]), .ZN(n1645) );
  INV_X1 U1807 ( .A(n1381), .ZN(n1644) );
  OAI222_X1 U1808 ( .A1(n2048), .A2(n2049), .B1(n2048), .B2(n2050), .C1(n2050), 
        .C2(n2049), .ZN(n2044) );
  INV_X1 U1809 ( .A(n610), .ZN(n2050) );
  XNOR2_X1 U1810 ( .A(n1674), .B(n2051), .ZN(n2049) );
  AOI221_X1 U1811 ( .B1(B[16]), .B2(n1558), .C1(B[15]), .C2(n1559), .A(n2052), 
        .ZN(n2051) );
  OAI22_X1 U1812 ( .A1(n1561), .A2(n1640), .B1(n1563), .B2(n1641), .ZN(n2052)
         );
  INV_X1 U1813 ( .A(B[14]), .ZN(n1641) );
  INV_X1 U1814 ( .A(n1382), .ZN(n1640) );
  AOI222_X1 U1815 ( .A1(n2053), .A2(n2054), .B1(n2053), .B2(n620), .C1(n620), 
        .C2(n2054), .ZN(n2048) );
  XNOR2_X1 U1816 ( .A(A[2]), .B(n2055), .ZN(n2054) );
  AOI221_X1 U1817 ( .B1(B[15]), .B2(n1558), .C1(B[14]), .C2(n1559), .A(n2056), 
        .ZN(n2055) );
  OAI22_X1 U1818 ( .A1(n1561), .A2(n1636), .B1(n1563), .B2(n1637), .ZN(n2056)
         );
  INV_X1 U1819 ( .A(B[13]), .ZN(n1637) );
  INV_X1 U1820 ( .A(n1383), .ZN(n1636) );
  OAI222_X1 U1821 ( .A1(n2057), .A2(n2058), .B1(n2057), .B2(n2059), .C1(n2059), 
        .C2(n2058), .ZN(n2053) );
  INV_X1 U1822 ( .A(n630), .ZN(n2059) );
  XNOR2_X1 U1823 ( .A(n1674), .B(n2060), .ZN(n2058) );
  AOI221_X1 U1824 ( .B1(B[14]), .B2(n1558), .C1(B[13]), .C2(n1559), .A(n2061), 
        .ZN(n2060) );
  OAI22_X1 U1825 ( .A1(n1561), .A2(n1632), .B1(n1563), .B2(n1633), .ZN(n2061)
         );
  INV_X1 U1826 ( .A(B[12]), .ZN(n1633) );
  INV_X1 U1827 ( .A(n1384), .ZN(n1632) );
  AOI222_X1 U1828 ( .A1(n2062), .A2(n2063), .B1(n2062), .B2(n638), .C1(n638), 
        .C2(n2063), .ZN(n2057) );
  XNOR2_X1 U1829 ( .A(A[2]), .B(n2064), .ZN(n2063) );
  AOI221_X1 U1830 ( .B1(B[13]), .B2(n1558), .C1(B[12]), .C2(n1559), .A(n2065), 
        .ZN(n2064) );
  OAI22_X1 U1831 ( .A1(n1561), .A2(n1628), .B1(n1563), .B2(n1629), .ZN(n2065)
         );
  INV_X1 U1832 ( .A(B[11]), .ZN(n1629) );
  INV_X1 U1833 ( .A(n1385), .ZN(n1628) );
  OAI222_X1 U1834 ( .A1(n2066), .A2(n2067), .B1(n2066), .B2(n2068), .C1(n2068), 
        .C2(n2067), .ZN(n2062) );
  INV_X1 U1835 ( .A(n646), .ZN(n2068) );
  XNOR2_X1 U1836 ( .A(n1674), .B(n2069), .ZN(n2067) );
  AOI221_X1 U1837 ( .B1(B[12]), .B2(n1558), .C1(B[11]), .C2(n1559), .A(n2070), 
        .ZN(n2069) );
  OAI22_X1 U1838 ( .A1(n1561), .A2(n1624), .B1(n1563), .B2(n1625), .ZN(n2070)
         );
  INV_X1 U1839 ( .A(B[10]), .ZN(n1625) );
  INV_X1 U1840 ( .A(n1386), .ZN(n1624) );
  AOI222_X1 U1841 ( .A1(n2071), .A2(n2072), .B1(n2071), .B2(n654), .C1(n654), 
        .C2(n2072), .ZN(n2066) );
  XNOR2_X1 U1842 ( .A(A[2]), .B(n2073), .ZN(n2072) );
  AOI221_X1 U1843 ( .B1(B[11]), .B2(n1558), .C1(B[10]), .C2(n1559), .A(n2074), 
        .ZN(n2073) );
  OAI22_X1 U1844 ( .A1(n1561), .A2(n1620), .B1(n1563), .B2(n1621), .ZN(n2074)
         );
  INV_X1 U1845 ( .A(B[9]), .ZN(n1621) );
  INV_X1 U1846 ( .A(n1387), .ZN(n1620) );
  OAI222_X1 U1847 ( .A1(n2075), .A2(n2076), .B1(n2075), .B2(n2077), .C1(n2077), 
        .C2(n2076), .ZN(n2071) );
  INV_X1 U1848 ( .A(n660), .ZN(n2077) );
  XNOR2_X1 U1849 ( .A(n1674), .B(n2078), .ZN(n2076) );
  AOI221_X1 U1850 ( .B1(B[10]), .B2(n1558), .C1(B[9]), .C2(n1559), .A(n2079), 
        .ZN(n2078) );
  OAI22_X1 U1851 ( .A1(n1561), .A2(n1616), .B1(n1563), .B2(n1617), .ZN(n2079)
         );
  INV_X1 U1852 ( .A(B[8]), .ZN(n1617) );
  INV_X1 U1853 ( .A(n1388), .ZN(n1616) );
  AOI222_X1 U1854 ( .A1(n2080), .A2(n2081), .B1(n2080), .B2(n666), .C1(n666), 
        .C2(n2081), .ZN(n2075) );
  XNOR2_X1 U1855 ( .A(A[2]), .B(n2082), .ZN(n2081) );
  AOI221_X1 U1856 ( .B1(B[9]), .B2(n1558), .C1(B[8]), .C2(n1559), .A(n2083), 
        .ZN(n2082) );
  OAI22_X1 U1857 ( .A1(n1561), .A2(n1612), .B1(n1563), .B2(n1613), .ZN(n2083)
         );
  INV_X1 U1858 ( .A(B[7]), .ZN(n1613) );
  INV_X1 U1859 ( .A(n1389), .ZN(n1612) );
  OAI222_X1 U1860 ( .A1(n2084), .A2(n2085), .B1(n2084), .B2(n2086), .C1(n2086), 
        .C2(n2085), .ZN(n2080) );
  INV_X1 U1861 ( .A(n672), .ZN(n2086) );
  XNOR2_X1 U1862 ( .A(n1674), .B(n2087), .ZN(n2085) );
  AOI221_X1 U1863 ( .B1(B[8]), .B2(n1558), .C1(B[7]), .C2(n1559), .A(n2088), 
        .ZN(n2087) );
  OAI22_X1 U1864 ( .A1(n1561), .A2(n1608), .B1(n1563), .B2(n1609), .ZN(n2088)
         );
  INV_X1 U1865 ( .A(B[6]), .ZN(n1609) );
  INV_X1 U1866 ( .A(n1390), .ZN(n1608) );
  AOI222_X1 U1867 ( .A1(n2089), .A2(n2090), .B1(n2089), .B2(n676), .C1(n676), 
        .C2(n2090), .ZN(n2084) );
  XNOR2_X1 U1868 ( .A(A[2]), .B(n2091), .ZN(n2090) );
  AOI221_X1 U1869 ( .B1(B[7]), .B2(n1558), .C1(B[6]), .C2(n1559), .A(n2092), 
        .ZN(n2091) );
  OAI22_X1 U1870 ( .A1(n1561), .A2(n1604), .B1(n1563), .B2(n1605), .ZN(n2092)
         );
  INV_X1 U1871 ( .A(B[5]), .ZN(n1605) );
  INV_X1 U1872 ( .A(n1391), .ZN(n1604) );
  OAI222_X1 U1873 ( .A1(n2093), .A2(n2094), .B1(n2093), .B2(n2095), .C1(n2095), 
        .C2(n2094), .ZN(n2089) );
  INV_X1 U1874 ( .A(n680), .ZN(n2095) );
  XNOR2_X1 U1875 ( .A(n1674), .B(n2096), .ZN(n2094) );
  AOI221_X1 U1876 ( .B1(B[6]), .B2(n1558), .C1(B[5]), .C2(n1559), .A(n2097), 
        .ZN(n2096) );
  OAI22_X1 U1877 ( .A1(n1561), .A2(n1600), .B1(n1563), .B2(n1601), .ZN(n2097)
         );
  INV_X1 U1878 ( .A(B[4]), .ZN(n1601) );
  INV_X1 U1879 ( .A(n1392), .ZN(n1600) );
  AOI222_X1 U1880 ( .A1(n2098), .A2(n2099), .B1(n2098), .B2(n684), .C1(n684), 
        .C2(n2099), .ZN(n2093) );
  XNOR2_X1 U1881 ( .A(A[2]), .B(n2100), .ZN(n2099) );
  AOI221_X1 U1882 ( .B1(B[5]), .B2(n1558), .C1(B[4]), .C2(n1559), .A(n2101), 
        .ZN(n2100) );
  OAI22_X1 U1883 ( .A1(n1561), .A2(n1596), .B1(n1563), .B2(n1597), .ZN(n2101)
         );
  INV_X1 U1884 ( .A(B[3]), .ZN(n1597) );
  INV_X1 U1885 ( .A(n1393), .ZN(n1596) );
  OAI222_X1 U1886 ( .A1(n2102), .A2(n2103), .B1(n2102), .B2(n2104), .C1(n2104), 
        .C2(n2103), .ZN(n2098) );
  INV_X1 U1887 ( .A(n686), .ZN(n2104) );
  XNOR2_X1 U1888 ( .A(n1674), .B(n2105), .ZN(n2103) );
  AOI221_X1 U1889 ( .B1(B[4]), .B2(n1558), .C1(B[3]), .C2(n1559), .A(n2106), 
        .ZN(n2105) );
  OAI22_X1 U1890 ( .A1(n1561), .A2(n1592), .B1(n1563), .B2(n1593), .ZN(n2106)
         );
  INV_X1 U1891 ( .A(B[2]), .ZN(n1593) );
  INV_X1 U1892 ( .A(n1394), .ZN(n1592) );
  AOI222_X1 U1893 ( .A1(n2107), .A2(n2108), .B1(n2107), .B2(n688), .C1(n688), 
        .C2(n2108), .ZN(n2102) );
  XNOR2_X1 U1894 ( .A(A[2]), .B(n2109), .ZN(n2108) );
  AOI221_X1 U1895 ( .B1(B[3]), .B2(n1558), .C1(B[2]), .C2(n1559), .A(n2110), 
        .ZN(n2109) );
  OAI22_X1 U1896 ( .A1(n1561), .A2(n1589), .B1(n1563), .B2(n1578), .ZN(n2110)
         );
  INV_X1 U1897 ( .A(B[1]), .ZN(n1578) );
  INV_X1 U1898 ( .A(n1395), .ZN(n1589) );
  AND2_X1 U1899 ( .A1(n2114), .A2(n2115), .ZN(n2107) );
  AOI211_X1 U1900 ( .C1(B[1]), .C2(n1558), .A(n2116), .B(B[0]), .ZN(n2115) );
  INV_X1 U1901 ( .A(n2117), .ZN(n2116) );
  AOI22_X1 U1902 ( .A1(n1558), .A2(B[2]), .B1(n2118), .B2(n1397), .ZN(n2117)
         );
  INV_X1 U1903 ( .A(A[0]), .ZN(n2112) );
  AOI221_X1 U1904 ( .B1(B[1]), .B2(n1559), .C1(n1396), .C2(n2118), .A(n1674), 
        .ZN(n2114) );
  INV_X1 U1905 ( .A(n1561), .ZN(n2118) );
  XNOR2_X1 U1906 ( .A(A[1]), .B(n1674), .ZN(n2111) );
  INV_X1 U1907 ( .A(A[2]), .ZN(n1674) );
  INV_X1 U1908 ( .A(A[1]), .ZN(n2113) );
  AOI21_X1 U1909 ( .B1(n2119), .B2(n2120), .A(n2121), .ZN(PRODUCT[47]) );
  OAI22_X1 U1910 ( .A1(n2122), .A2(n2123), .B1(n2122), .B2(n2124), .ZN(n2121)
         );
  INV_X1 U1911 ( .A(n2120), .ZN(n2124) );
  AOI222_X1 U1912 ( .A1(n2024), .A2(n303), .B1(n2123), .B2(n303), .C1(n2024), 
        .C2(n2123), .ZN(n2122) );
  XOR2_X1 U1913 ( .A(n1541), .B(n2125), .Z(n2024) );
  AOI221_X1 U1914 ( .B1(n1537), .B2(B[23]), .C1(n1536), .C2(B[22]), .A(n2126), 
        .ZN(n2125) );
  OAI22_X1 U1915 ( .A1(n1567), .A2(n1976), .B1(n1568), .B2(n1538), .ZN(n2126)
         );
  INV_X1 U1916 ( .A(B[21]), .ZN(n1568) );
  INV_X1 U1917 ( .A(n1375), .ZN(n1567) );
  XOR2_X1 U1918 ( .A(n2127), .B(n1541), .Z(n2120) );
  OAI221_X1 U1919 ( .B1(n1556), .B2(n1539), .C1(n1556), .C2(n1976), .A(n2128), 
        .ZN(n2127) );
  OAI21_X1 U1920 ( .B1(n1537), .B2(n1536), .A(n1554), .ZN(n2128) );
  INV_X1 U1921 ( .A(n2123), .ZN(n2119) );
  XOR2_X1 U1922 ( .A(A[23]), .B(n2129), .Z(n2123) );
  AOI221_X1 U1923 ( .B1(n1537), .B2(n1554), .C1(n1536), .C2(n1554), .A(n2130), 
        .ZN(n2129) );
  OAI22_X1 U1924 ( .A1(n1571), .A2(n1976), .B1(n1572), .B2(n1538), .ZN(n2130)
         );
  NAND3_X1 U1925 ( .A1(n2131), .A2(n2132), .A3(n2133), .ZN(n1980) );
  INV_X1 U1926 ( .A(B[22]), .ZN(n1572) );
  INV_X1 U1927 ( .A(n1374), .ZN(n1571) );
  XNOR2_X1 U1928 ( .A(A[21]), .B(A[22]), .ZN(n2133) );
  INV_X1 U1929 ( .A(n2131), .ZN(n2134) );
  XOR2_X1 U1930 ( .A(A[21]), .B(n1543), .Z(n2131) );
  XNOR2_X1 U1931 ( .A(A[22]), .B(n1541), .ZN(n2132) );
endmodule


module iir_filter_DW02_mult_0 ( A, B, PRODUCT, TC );
  input [23:0] A;
  input [23:0] B;
  output [47:0] PRODUCT;
  input TC;
  wire   n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n351, n352, n353, n354, n355, n356, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n906, n907, n908, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134;

  FA_X1 U182 ( .A(n351), .B(n352), .CI(n304), .CO(n303), .S(PRODUCT[44]) );
  FA_X1 U183 ( .A(n353), .B(n354), .CI(n305), .CO(n304), .S(PRODUCT[43]) );
  FA_X1 U184 ( .A(n355), .B(n358), .CI(n306), .CO(n305), .S(PRODUCT[42]) );
  FA_X1 U185 ( .A(n359), .B(n361), .CI(n307), .CO(n306), .S(PRODUCT[41]) );
  FA_X1 U186 ( .A(n362), .B(n364), .CI(n308), .CO(n307), .S(PRODUCT[40]) );
  FA_X1 U187 ( .A(n365), .B(n370), .CI(n309), .CO(n308), .S(PRODUCT[39]) );
  FA_X1 U188 ( .A(n371), .B(n375), .CI(n310), .CO(n309), .S(PRODUCT[38]) );
  FA_X1 U189 ( .A(n376), .B(n381), .CI(n311), .CO(n310), .S(PRODUCT[37]) );
  FA_X1 U190 ( .A(n382), .B(n389), .CI(n312), .CO(n311), .S(PRODUCT[36]) );
  FA_X1 U191 ( .A(n390), .B(n396), .CI(n313), .CO(n312), .S(PRODUCT[35]) );
  FA_X1 U192 ( .A(n397), .B(n403), .CI(n314), .CO(n313), .S(PRODUCT[34]) );
  FA_X1 U193 ( .A(n404), .B(n413), .CI(n315), .CO(n314), .S(PRODUCT[33]) );
  FA_X1 U194 ( .A(n414), .B(n422), .CI(n316), .CO(n315), .S(PRODUCT[32]) );
  FA_X1 U195 ( .A(n423), .B(n432), .CI(n317), .CO(n316), .S(PRODUCT[31]) );
  FA_X1 U196 ( .A(n433), .B(n444), .CI(n318), .CO(n317), .S(PRODUCT[30]) );
  FA_X1 U197 ( .A(n445), .B(n455), .CI(n319), .CO(n318), .S(PRODUCT[29]) );
  FA_X1 U198 ( .A(n456), .B(n467), .CI(n320), .CO(n319), .S(PRODUCT[28]) );
  FA_X1 U199 ( .A(n468), .B(n481), .CI(n321), .CO(n320), .S(PRODUCT[27]) );
  FA_X1 U200 ( .A(n482), .B(n494), .CI(n322), .CO(n321), .S(PRODUCT[26]) );
  FA_X1 U201 ( .A(n495), .B(n507), .CI(n323), .CO(n322), .S(PRODUCT[25]) );
  FA_X1 U202 ( .A(n508), .B(n906), .CI(n324), .CO(n323), .S(PRODUCT[24]) );
  FA_X1 U203 ( .A(n907), .B(n522), .CI(n325), .CO(n324), .S(PRODUCT[23]) );
  FA_X1 U204 ( .A(n908), .B(n536), .CI(n326), .CO(n325), .S(PRODUCT[22]) );
  FA_X1 U235 ( .A(n356), .B(n749), .CI(n729), .CO(n352), .S(n353) );
  FA_X1 U236 ( .A(n730), .B(n360), .CI(n750), .CO(n354), .S(n355) );
  FA_X1 U238 ( .A(n360), .B(n731), .CI(n751), .CO(n358), .S(n359) );
  FA_X1 U240 ( .A(n752), .B(n363), .CI(n366), .CO(n361), .S(n362) );
  FA_X1 U241 ( .A(n368), .B(n775), .CI(n732), .CO(n356), .S(n363) );
  FA_X1 U242 ( .A(n776), .B(n753), .CI(n367), .CO(n364), .S(n365) );
  FA_X1 U243 ( .A(n733), .B(n374), .CI(n372), .CO(n366), .S(n367) );
  FA_X1 U245 ( .A(n373), .B(n377), .CI(n777), .CO(n370), .S(n371) );
  FA_X1 U246 ( .A(n374), .B(n379), .CI(n754), .CO(n372), .S(n373) );
  FA_X1 U248 ( .A(n778), .B(n378), .CI(n383), .CO(n375), .S(n376) );
  FA_X1 U249 ( .A(n385), .B(n380), .CI(n755), .CO(n377), .S(n378) );
  FA_X1 U250 ( .A(n387), .B(n801), .CI(n734), .CO(n379), .S(n380) );
  FA_X1 U251 ( .A(n802), .B(n779), .CI(n384), .CO(n381), .S(n382) );
  FA_X1 U252 ( .A(n386), .B(n393), .CI(n391), .CO(n383), .S(n384) );
  FA_X1 U253 ( .A(n735), .B(n395), .CI(n756), .CO(n385), .S(n386) );
  FA_X1 U255 ( .A(n392), .B(n398), .CI(n803), .CO(n389), .S(n390) );
  FA_X1 U256 ( .A(n394), .B(n400), .CI(n780), .CO(n391), .S(n392) );
  FA_X1 U257 ( .A(n395), .B(n736), .CI(n757), .CO(n393), .S(n394) );
  FA_X1 U259 ( .A(n804), .B(n399), .CI(n405), .CO(n396), .S(n397) );
  FA_X1 U260 ( .A(n407), .B(n401), .CI(n781), .CO(n398), .S(n399) );
  FA_X1 U261 ( .A(n758), .B(n402), .CI(n409), .CO(n400), .S(n401) );
  FA_X1 U262 ( .A(n411), .B(n827), .CI(n737), .CO(n387), .S(n402) );
  FA_X1 U263 ( .A(n828), .B(n805), .CI(n406), .CO(n403), .S(n404) );
  FA_X1 U264 ( .A(n408), .B(n417), .CI(n415), .CO(n405), .S(n406) );
  FA_X1 U265 ( .A(n410), .B(n759), .CI(n782), .CO(n407), .S(n408) );
  FA_X1 U266 ( .A(n738), .B(n421), .CI(n419), .CO(n409), .S(n410) );
  FA_X1 U268 ( .A(n416), .B(n424), .CI(n829), .CO(n413), .S(n414) );
  FA_X1 U269 ( .A(n418), .B(n426), .CI(n806), .CO(n415), .S(n416) );
  FA_X1 U270 ( .A(n420), .B(n428), .CI(n783), .CO(n417), .S(n418) );
  FA_X1 U271 ( .A(n421), .B(n430), .CI(n760), .CO(n419), .S(n420) );
  FA_X1 U273 ( .A(n830), .B(n425), .CI(n434), .CO(n422), .S(n423) );
  FA_X1 U274 ( .A(n436), .B(n427), .CI(n807), .CO(n424), .S(n425) );
  FA_X1 U275 ( .A(n784), .B(n429), .CI(n438), .CO(n426), .S(n427) );
  FA_X1 U276 ( .A(n440), .B(n431), .CI(n761), .CO(n428), .S(n429) );
  FA_X1 U277 ( .A(n442), .B(n853), .CI(n739), .CO(n430), .S(n431) );
  FA_X1 U278 ( .A(n854), .B(n831), .CI(n435), .CO(n432), .S(n433) );
  FA_X1 U279 ( .A(n437), .B(n448), .CI(n446), .CO(n434), .S(n435) );
  FA_X1 U280 ( .A(n439), .B(n785), .CI(n808), .CO(n436), .S(n437) );
  FA_X1 U281 ( .A(n441), .B(n452), .CI(n450), .CO(n438), .S(n439) );
  FA_X1 U282 ( .A(n740), .B(n454), .CI(n762), .CO(n440), .S(n441) );
  FA_X1 U284 ( .A(n447), .B(n457), .CI(n855), .CO(n444), .S(n445) );
  FA_X1 U285 ( .A(n449), .B(n459), .CI(n832), .CO(n446), .S(n447) );
  FA_X1 U286 ( .A(n451), .B(n461), .CI(n809), .CO(n448), .S(n449) );
  FA_X1 U287 ( .A(n453), .B(n463), .CI(n786), .CO(n450), .S(n451) );
  FA_X1 U288 ( .A(n454), .B(n465), .CI(n763), .CO(n452), .S(n453) );
  FA_X1 U290 ( .A(n856), .B(n458), .CI(n469), .CO(n455), .S(n456) );
  FA_X1 U291 ( .A(n471), .B(n460), .CI(n833), .CO(n457), .S(n458) );
  FA_X1 U292 ( .A(n810), .B(n462), .CI(n473), .CO(n459), .S(n460) );
  FA_X1 U293 ( .A(n475), .B(n464), .CI(n787), .CO(n461), .S(n462) );
  FA_X1 U294 ( .A(n764), .B(n466), .CI(n477), .CO(n463), .S(n464) );
  FA_X1 U295 ( .A(n479), .B(n879), .CI(n741), .CO(n465), .S(n466) );
  FA_X1 U296 ( .A(n880), .B(n857), .CI(n470), .CO(n467), .S(n468) );
  FA_X1 U297 ( .A(n472), .B(n485), .CI(n483), .CO(n469), .S(n470) );
  FA_X1 U298 ( .A(n474), .B(n811), .CI(n834), .CO(n471), .S(n472) );
  FA_X1 U299 ( .A(n476), .B(n489), .CI(n487), .CO(n473), .S(n474) );
  FA_X1 U300 ( .A(n478), .B(n765), .CI(n788), .CO(n475), .S(n476) );
  FA_X1 U301 ( .A(n742), .B(n493), .CI(n491), .CO(n477), .S(n478) );
  FA_X1 U303 ( .A(n484), .B(n858), .CI(n881), .CO(n481), .S(n482) );
  FA_X1 U304 ( .A(n486), .B(n498), .CI(n496), .CO(n483), .S(n484) );
  FA_X1 U305 ( .A(n488), .B(n812), .CI(n835), .CO(n485), .S(n486) );
  FA_X1 U306 ( .A(n490), .B(n502), .CI(n500), .CO(n487), .S(n488) );
  FA_X1 U307 ( .A(n492), .B(n504), .CI(n789), .CO(n489), .S(n490) );
  FA_X1 U308 ( .A(n743), .B(n493), .CI(n766), .CO(n491), .S(n492) );
  FA_X1 U310 ( .A(n497), .B(n509), .CI(n882), .CO(n494), .S(n495) );
  FA_X1 U311 ( .A(n499), .B(n511), .CI(n859), .CO(n496), .S(n497) );
  FA_X1 U312 ( .A(n501), .B(n513), .CI(n836), .CO(n498), .S(n499) );
  FA_X1 U313 ( .A(n503), .B(n515), .CI(n813), .CO(n500), .S(n501) );
  FA_X1 U314 ( .A(n505), .B(n517), .CI(n790), .CO(n502), .S(n503) );
  FA_X1 U315 ( .A(n506), .B(n744), .CI(n767), .CO(n504), .S(n505) );
  FA_X1 U318 ( .A(n883), .B(n510), .CI(n521), .CO(n507), .S(n508) );
  FA_X1 U319 ( .A(n860), .B(n512), .CI(n523), .CO(n509), .S(n510) );
  FA_X1 U320 ( .A(n837), .B(n514), .CI(n525), .CO(n511), .S(n512) );
  FA_X1 U321 ( .A(n814), .B(n516), .CI(n527), .CO(n513), .S(n514) );
  FA_X1 U322 ( .A(n791), .B(n518), .CI(n529), .CO(n515), .S(n516) );
  FA_X1 U323 ( .A(n768), .B(n520), .CI(n531), .CO(n517), .S(n518) );
  HA_X1 U324 ( .A(n533), .B(n745), .CO(n519), .S(n520) );
  FA_X1 U325 ( .A(n884), .B(n524), .CI(n535), .CO(n521), .S(n522) );
  FA_X1 U326 ( .A(n861), .B(n526), .CI(n537), .CO(n523), .S(n524) );
  FA_X1 U327 ( .A(n838), .B(n528), .CI(n539), .CO(n525), .S(n526) );
  FA_X1 U328 ( .A(n815), .B(n530), .CI(n541), .CO(n527), .S(n528) );
  FA_X1 U329 ( .A(n792), .B(n532), .CI(n543), .CO(n529), .S(n530) );
  FA_X1 U330 ( .A(n769), .B(n534), .CI(n545), .CO(n531), .S(n532) );
  HA_X1 U331 ( .A(n547), .B(n746), .CO(n533), .S(n534) );
  FA_X1 U332 ( .A(n885), .B(n538), .CI(n549), .CO(n535), .S(n536) );
  FA_X1 U333 ( .A(n862), .B(n540), .CI(n551), .CO(n537), .S(n538) );
  FA_X1 U334 ( .A(n839), .B(n542), .CI(n553), .CO(n539), .S(n540) );
  FA_X1 U335 ( .A(n816), .B(n544), .CI(n555), .CO(n541), .S(n542) );
  FA_X1 U336 ( .A(n793), .B(n546), .CI(n557), .CO(n543), .S(n544) );
  FA_X1 U337 ( .A(n770), .B(n548), .CI(n559), .CO(n545), .S(n546) );
  HA_X1 U338 ( .A(n561), .B(n747), .CO(n547), .S(n548) );
  FA_X1 U339 ( .A(n886), .B(n552), .CI(n563), .CO(n549), .S(n550) );
  FA_X1 U340 ( .A(n863), .B(n554), .CI(n565), .CO(n551), .S(n552) );
  FA_X1 U341 ( .A(n840), .B(n556), .CI(n567), .CO(n553), .S(n554) );
  FA_X1 U342 ( .A(n817), .B(n558), .CI(n569), .CO(n555), .S(n556) );
  FA_X1 U343 ( .A(n794), .B(n560), .CI(n571), .CO(n557), .S(n558) );
  FA_X1 U344 ( .A(n771), .B(n562), .CI(n573), .CO(n559), .S(n560) );
  HA_X1 U345 ( .A(n748), .B(n1540), .CO(n561), .S(n562) );
  FA_X1 U346 ( .A(n887), .B(n566), .CI(n575), .CO(n563), .S(n564) );
  FA_X1 U347 ( .A(n864), .B(n568), .CI(n577), .CO(n565), .S(n566) );
  FA_X1 U348 ( .A(n841), .B(n570), .CI(n579), .CO(n567), .S(n568) );
  FA_X1 U349 ( .A(n818), .B(n572), .CI(n581), .CO(n569), .S(n570) );
  FA_X1 U350 ( .A(n795), .B(n574), .CI(n583), .CO(n571), .S(n572) );
  HA_X1 U351 ( .A(n585), .B(n772), .CO(n573), .S(n574) );
  FA_X1 U352 ( .A(n888), .B(n578), .CI(n587), .CO(n575), .S(n576) );
  FA_X1 U353 ( .A(n865), .B(n580), .CI(n589), .CO(n577), .S(n578) );
  FA_X1 U354 ( .A(n842), .B(n582), .CI(n591), .CO(n579), .S(n580) );
  FA_X1 U355 ( .A(n819), .B(n584), .CI(n593), .CO(n581), .S(n582) );
  FA_X1 U356 ( .A(n796), .B(n586), .CI(n595), .CO(n583), .S(n584) );
  HA_X1 U357 ( .A(n597), .B(n773), .CO(n585), .S(n586) );
  FA_X1 U358 ( .A(n889), .B(n590), .CI(n599), .CO(n587), .S(n588) );
  FA_X1 U359 ( .A(n866), .B(n592), .CI(n601), .CO(n589), .S(n590) );
  FA_X1 U360 ( .A(n843), .B(n594), .CI(n603), .CO(n591), .S(n592) );
  FA_X1 U361 ( .A(n820), .B(n596), .CI(n605), .CO(n593), .S(n594) );
  FA_X1 U362 ( .A(n797), .B(n598), .CI(n607), .CO(n595), .S(n596) );
  HA_X1 U363 ( .A(n774), .B(n1542), .CO(n597), .S(n598) );
  FA_X1 U364 ( .A(n890), .B(n602), .CI(n609), .CO(n599), .S(n600) );
  FA_X1 U365 ( .A(n867), .B(n604), .CI(n611), .CO(n601), .S(n602) );
  FA_X1 U366 ( .A(n844), .B(n606), .CI(n613), .CO(n603), .S(n604) );
  FA_X1 U367 ( .A(n821), .B(n608), .CI(n615), .CO(n605), .S(n606) );
  HA_X1 U368 ( .A(n617), .B(n798), .CO(n607), .S(n608) );
  FA_X1 U369 ( .A(n891), .B(n612), .CI(n619), .CO(n609), .S(n610) );
  FA_X1 U370 ( .A(n868), .B(n614), .CI(n621), .CO(n611), .S(n612) );
  FA_X1 U371 ( .A(n845), .B(n616), .CI(n623), .CO(n613), .S(n614) );
  FA_X1 U372 ( .A(n822), .B(n618), .CI(n625), .CO(n615), .S(n616) );
  HA_X1 U373 ( .A(n627), .B(n799), .CO(n617), .S(n618) );
  FA_X1 U374 ( .A(n892), .B(n622), .CI(n629), .CO(n619), .S(n620) );
  FA_X1 U375 ( .A(n869), .B(n624), .CI(n631), .CO(n621), .S(n622) );
  FA_X1 U376 ( .A(n846), .B(n626), .CI(n633), .CO(n623), .S(n624) );
  FA_X1 U377 ( .A(n823), .B(n628), .CI(n635), .CO(n625), .S(n626) );
  HA_X1 U378 ( .A(n800), .B(n1544), .CO(n627), .S(n628) );
  FA_X1 U379 ( .A(n893), .B(n632), .CI(n637), .CO(n629), .S(n630) );
  FA_X1 U380 ( .A(n870), .B(n634), .CI(n639), .CO(n631), .S(n632) );
  FA_X1 U381 ( .A(n847), .B(n636), .CI(n641), .CO(n633), .S(n634) );
  HA_X1 U382 ( .A(n643), .B(n824), .CO(n635), .S(n636) );
  FA_X1 U383 ( .A(n894), .B(n640), .CI(n645), .CO(n637), .S(n638) );
  FA_X1 U384 ( .A(n871), .B(n642), .CI(n647), .CO(n639), .S(n640) );
  FA_X1 U385 ( .A(n848), .B(n644), .CI(n649), .CO(n641), .S(n642) );
  HA_X1 U386 ( .A(n651), .B(n825), .CO(n643), .S(n644) );
  FA_X1 U387 ( .A(n895), .B(n648), .CI(n653), .CO(n645), .S(n646) );
  FA_X1 U388 ( .A(n872), .B(n650), .CI(n655), .CO(n647), .S(n648) );
  FA_X1 U389 ( .A(n849), .B(n652), .CI(n657), .CO(n649), .S(n650) );
  HA_X1 U390 ( .A(n826), .B(n1546), .CO(n651), .S(n652) );
  FA_X1 U391 ( .A(n896), .B(n656), .CI(n659), .CO(n653), .S(n654) );
  FA_X1 U392 ( .A(n873), .B(n658), .CI(n661), .CO(n655), .S(n656) );
  HA_X1 U393 ( .A(n663), .B(n850), .CO(n657), .S(n658) );
  FA_X1 U394 ( .A(n897), .B(n662), .CI(n665), .CO(n659), .S(n660) );
  FA_X1 U395 ( .A(n874), .B(n664), .CI(n667), .CO(n661), .S(n662) );
  HA_X1 U396 ( .A(n669), .B(n851), .CO(n663), .S(n664) );
  FA_X1 U397 ( .A(n898), .B(n668), .CI(n671), .CO(n665), .S(n666) );
  FA_X1 U398 ( .A(n875), .B(n670), .CI(n673), .CO(n667), .S(n668) );
  HA_X1 U399 ( .A(n852), .B(n1548), .CO(n669), .S(n670) );
  FA_X1 U400 ( .A(n899), .B(n674), .CI(n675), .CO(n671), .S(n672) );
  HA_X1 U401 ( .A(n677), .B(n876), .CO(n673), .S(n674) );
  FA_X1 U402 ( .A(n900), .B(n678), .CI(n679), .CO(n675), .S(n676) );
  HA_X1 U403 ( .A(n681), .B(n877), .CO(n677), .S(n678) );
  FA_X1 U404 ( .A(n901), .B(n682), .CI(n683), .CO(n679), .S(n680) );
  HA_X1 U405 ( .A(n878), .B(n1550), .CO(n681), .S(n682) );
  HA_X1 U406 ( .A(n685), .B(n902), .CO(n683), .S(n684) );
  HA_X1 U407 ( .A(n687), .B(n903), .CO(n685), .S(n686) );
  HA_X1 U408 ( .A(n904), .B(n1552), .CO(n687), .S(n688) );
  FA_X1 U1112 ( .A(B[22]), .B(n1554), .CI(n706), .CO(n1374), .S(n1375) );
  FA_X1 U1113 ( .A(B[21]), .B(B[22]), .CI(n707), .CO(n706), .S(n1376) );
  FA_X1 U1114 ( .A(B[20]), .B(B[21]), .CI(n708), .CO(n707), .S(n1377) );
  FA_X1 U1115 ( .A(B[19]), .B(B[20]), .CI(n709), .CO(n708), .S(n1378) );
  FA_X1 U1116 ( .A(B[18]), .B(B[19]), .CI(n710), .CO(n709), .S(n1379) );
  FA_X1 U1117 ( .A(B[17]), .B(B[18]), .CI(n711), .CO(n710), .S(n1380) );
  FA_X1 U1118 ( .A(B[16]), .B(B[17]), .CI(n712), .CO(n711), .S(n1381) );
  FA_X1 U1119 ( .A(B[15]), .B(B[16]), .CI(n713), .CO(n712), .S(n1382) );
  FA_X1 U1120 ( .A(B[14]), .B(B[15]), .CI(n714), .CO(n713), .S(n1383) );
  FA_X1 U1121 ( .A(B[13]), .B(B[14]), .CI(n715), .CO(n714), .S(n1384) );
  FA_X1 U1122 ( .A(B[12]), .B(B[13]), .CI(n716), .CO(n715), .S(n1385) );
  FA_X1 U1123 ( .A(B[11]), .B(B[12]), .CI(n717), .CO(n716), .S(n1386) );
  FA_X1 U1124 ( .A(B[10]), .B(B[11]), .CI(n718), .CO(n717), .S(n1387) );
  FA_X1 U1125 ( .A(B[9]), .B(B[10]), .CI(n719), .CO(n718), .S(n1388) );
  FA_X1 U1126 ( .A(B[8]), .B(B[9]), .CI(n720), .CO(n719), .S(n1389) );
  FA_X1 U1127 ( .A(B[7]), .B(B[8]), .CI(n721), .CO(n720), .S(n1390) );
  FA_X1 U1128 ( .A(B[6]), .B(B[7]), .CI(n722), .CO(n721), .S(n1391) );
  FA_X1 U1129 ( .A(B[5]), .B(B[6]), .CI(n723), .CO(n722), .S(n1392) );
  FA_X1 U1130 ( .A(B[4]), .B(B[5]), .CI(n724), .CO(n723), .S(n1393) );
  FA_X1 U1131 ( .A(B[3]), .B(B[4]), .CI(n725), .CO(n724), .S(n1394) );
  FA_X1 U1132 ( .A(B[2]), .B(B[3]), .CI(n726), .CO(n725), .S(n1395) );
  FA_X1 U1133 ( .A(B[1]), .B(B[2]), .CI(n727), .CO(n726), .S(n1396) );
  HA_X1 U1134 ( .A(B[0]), .B(B[1]), .CO(n727), .S(n1397) );
  OR2_X1 U1138 ( .A1(n2134), .A2(n2133), .ZN(n1534) );
  INV_X1 U1139 ( .A(n1534), .ZN(n1536) );
  INV_X1 U1140 ( .A(n1535), .ZN(n1537) );
  BUF_X1 U1141 ( .A(n1980), .Z(n1538) );
  BUF_X1 U1142 ( .A(n1980), .Z(n1539) );
  NAND3_X1 U1143 ( .A1(n1673), .A2(n1672), .A3(n1671), .ZN(n1586) );
  NAND3_X1 U1144 ( .A1(n1854), .A2(n1853), .A3(n1852), .ZN(n1804) );
  NAND3_X1 U1145 ( .A1(n1794), .A2(n1793), .A3(n1792), .ZN(n1744) );
  NAND3_X1 U1146 ( .A1(n1734), .A2(n1733), .A3(n1732), .ZN(n1684) );
  NAND3_X1 U1147 ( .A1(n2111), .A2(n2112), .A3(n2113), .ZN(n1563) );
  NAND2_X1 U1148 ( .A1(n1911), .A2(n1913), .ZN(n1857) );
  NAND2_X1 U1149 ( .A1(n1851), .A2(n1853), .ZN(n1797) );
  NAND2_X1 U1150 ( .A1(n1791), .A2(n1793), .ZN(n1737) );
  NAND2_X1 U1151 ( .A1(n1731), .A2(n1733), .ZN(n1677) );
  INV_X1 U1152 ( .A(n1553), .ZN(n1552) );
  INV_X1 U1153 ( .A(n1549), .ZN(n1548) );
  INV_X1 U1154 ( .A(n1551), .ZN(n1550) );
  NAND3_X1 U1155 ( .A1(n1914), .A2(n1913), .A3(n1912), .ZN(n1864) );
  NAND3_X1 U1156 ( .A1(n1974), .A2(n1973), .A3(n1972), .ZN(n1924) );
  NAND2_X1 U1157 ( .A1(n2134), .A2(n2132), .ZN(n1976) );
  NAND2_X1 U1158 ( .A1(n1971), .A2(n1973), .ZN(n1917) );
  INV_X1 U1159 ( .A(n1541), .ZN(n1540) );
  INV_X1 U1160 ( .A(n1543), .ZN(n1542) );
  INV_X1 U1161 ( .A(n1545), .ZN(n1544) );
  INV_X1 U1162 ( .A(n1547), .ZN(n1546) );
  INV_X1 U1163 ( .A(n1555), .ZN(n1554) );
  OR2_X1 U1164 ( .A1(n2132), .A2(n2131), .ZN(n1535) );
  NAND2_X1 U1165 ( .A1(A[0]), .A2(n2111), .ZN(n1561) );
  INV_X2 U1166 ( .A(B[0]), .ZN(n1574) );
  INV_X1 U1167 ( .A(A[5]), .ZN(n1553) );
  INV_X1 U1168 ( .A(A[11]), .ZN(n1549) );
  INV_X1 U1169 ( .A(A[8]), .ZN(n1551) );
  INV_X1 U1170 ( .A(A[17]), .ZN(n1545) );
  INV_X1 U1171 ( .A(A[14]), .ZN(n1547) );
  INV_X1 U1172 ( .A(A[23]), .ZN(n1541) );
  INV_X1 U1173 ( .A(A[20]), .ZN(n1543) );
  NOR2_X4 U1174 ( .A1(n1670), .A2(n1671), .ZN(n1581) );
  NOR2_X4 U1175 ( .A1(n1672), .A2(n1673), .ZN(n1582) );
  NAND2_X2 U1176 ( .A1(n1670), .A2(n1672), .ZN(n1576) );
  NOR2_X4 U1177 ( .A1(n1731), .A2(n1732), .ZN(n1680) );
  NOR2_X4 U1178 ( .A1(n1733), .A2(n1734), .ZN(n1681) );
  NOR2_X4 U1179 ( .A1(n1791), .A2(n1792), .ZN(n1740) );
  NOR2_X4 U1180 ( .A1(n1793), .A2(n1794), .ZN(n1741) );
  NOR2_X4 U1181 ( .A1(n1851), .A2(n1852), .ZN(n1800) );
  NOR2_X4 U1182 ( .A1(n1853), .A2(n1854), .ZN(n1801) );
  NOR2_X4 U1183 ( .A1(n1911), .A2(n1912), .ZN(n1860) );
  NOR2_X4 U1184 ( .A1(n1913), .A2(n1914), .ZN(n1861) );
  NOR2_X4 U1185 ( .A1(n1971), .A2(n1972), .ZN(n1920) );
  NOR2_X4 U1186 ( .A1(n1973), .A2(n1974), .ZN(n1921) );
  NOR2_X4 U1187 ( .A1(n2112), .A2(n2111), .ZN(n1558) );
  NOR2_X4 U1188 ( .A1(n2113), .A2(A[0]), .ZN(n1559) );
  INV_X1 U1189 ( .A(B[23]), .ZN(n1555) );
  INV_X1 U1190 ( .A(B[23]), .ZN(n1556) );
  XNOR2_X1 U1191 ( .A(A[2]), .B(n1557), .ZN(n908) );
  AOI221_X1 U1192 ( .B1(B[22]), .B2(n1558), .C1(B[21]), .C2(n1559), .A(n1560), 
        .ZN(n1557) );
  OAI22_X1 U1193 ( .A1(n1561), .A2(n1562), .B1(n1563), .B2(n1564), .ZN(n1560)
         );
  XNOR2_X1 U1194 ( .A(A[2]), .B(n1565), .ZN(n907) );
  AOI221_X1 U1195 ( .B1(B[23]), .B2(n1558), .C1(n1559), .C2(B[22]), .A(n1566), 
        .ZN(n1565) );
  OAI22_X1 U1196 ( .A1(n1561), .A2(n1567), .B1(n1568), .B2(n1563), .ZN(n1566)
         );
  XNOR2_X1 U1197 ( .A(A[2]), .B(n1569), .ZN(n906) );
  AOI221_X1 U1198 ( .B1(B[23]), .B2(n1558), .C1(n1554), .C2(n1559), .A(n1570), 
        .ZN(n1569) );
  OAI22_X1 U1199 ( .A1(n1561), .A2(n1571), .B1(n1572), .B2(n1563), .ZN(n1570)
         );
  XNOR2_X1 U1200 ( .A(n1573), .B(n1553), .ZN(n904) );
  OAI22_X1 U1201 ( .A1(n1574), .A2(n1575), .B1(n1576), .B2(n1574), .ZN(n1573)
         );
  XNOR2_X1 U1202 ( .A(n1577), .B(n1553), .ZN(n903) );
  OAI222_X1 U1203 ( .A1(n1575), .A2(n1578), .B1(n1574), .B2(n1579), .C1(n1576), 
        .C2(n1580), .ZN(n1577) );
  INV_X1 U1204 ( .A(n1581), .ZN(n1579) );
  INV_X1 U1205 ( .A(n1582), .ZN(n1575) );
  XNOR2_X1 U1206 ( .A(n1552), .B(n1583), .ZN(n902) );
  AOI221_X1 U1207 ( .B1(B[2]), .B2(n1582), .C1(B[1]), .C2(n1581), .A(n1584), 
        .ZN(n1583) );
  OAI22_X1 U1208 ( .A1(n1576), .A2(n1585), .B1(n1574), .B2(n1586), .ZN(n1584)
         );
  XNOR2_X1 U1209 ( .A(n1552), .B(n1587), .ZN(n901) );
  AOI221_X1 U1210 ( .B1(B[3]), .B2(n1582), .C1(B[2]), .C2(n1581), .A(n1588), 
        .ZN(n1587) );
  OAI22_X1 U1211 ( .A1(n1576), .A2(n1589), .B1(n1578), .B2(n1586), .ZN(n1588)
         );
  XNOR2_X1 U1212 ( .A(n1552), .B(n1590), .ZN(n900) );
  AOI221_X1 U1213 ( .B1(B[4]), .B2(n1582), .C1(B[3]), .C2(n1581), .A(n1591), 
        .ZN(n1590) );
  OAI22_X1 U1214 ( .A1(n1576), .A2(n1592), .B1(n1593), .B2(n1586), .ZN(n1591)
         );
  XNOR2_X1 U1215 ( .A(n1552), .B(n1594), .ZN(n899) );
  AOI221_X1 U1216 ( .B1(B[5]), .B2(n1582), .C1(B[4]), .C2(n1581), .A(n1595), 
        .ZN(n1594) );
  OAI22_X1 U1217 ( .A1(n1576), .A2(n1596), .B1(n1586), .B2(n1597), .ZN(n1595)
         );
  XNOR2_X1 U1218 ( .A(n1552), .B(n1598), .ZN(n898) );
  AOI221_X1 U1219 ( .B1(B[6]), .B2(n1582), .C1(B[5]), .C2(n1581), .A(n1599), 
        .ZN(n1598) );
  OAI22_X1 U1220 ( .A1(n1576), .A2(n1600), .B1(n1586), .B2(n1601), .ZN(n1599)
         );
  XNOR2_X1 U1221 ( .A(n1552), .B(n1602), .ZN(n897) );
  AOI221_X1 U1222 ( .B1(B[7]), .B2(n1582), .C1(B[6]), .C2(n1581), .A(n1603), 
        .ZN(n1602) );
  OAI22_X1 U1223 ( .A1(n1576), .A2(n1604), .B1(n1586), .B2(n1605), .ZN(n1603)
         );
  XNOR2_X1 U1224 ( .A(n1552), .B(n1606), .ZN(n896) );
  AOI221_X1 U1225 ( .B1(B[8]), .B2(n1582), .C1(B[7]), .C2(n1581), .A(n1607), 
        .ZN(n1606) );
  OAI22_X1 U1226 ( .A1(n1576), .A2(n1608), .B1(n1586), .B2(n1609), .ZN(n1607)
         );
  XNOR2_X1 U1227 ( .A(n1552), .B(n1610), .ZN(n895) );
  AOI221_X1 U1228 ( .B1(B[9]), .B2(n1582), .C1(B[8]), .C2(n1581), .A(n1611), 
        .ZN(n1610) );
  OAI22_X1 U1229 ( .A1(n1576), .A2(n1612), .B1(n1586), .B2(n1613), .ZN(n1611)
         );
  XNOR2_X1 U1230 ( .A(n1552), .B(n1614), .ZN(n894) );
  AOI221_X1 U1231 ( .B1(B[10]), .B2(n1582), .C1(B[9]), .C2(n1581), .A(n1615), 
        .ZN(n1614) );
  OAI22_X1 U1232 ( .A1(n1576), .A2(n1616), .B1(n1586), .B2(n1617), .ZN(n1615)
         );
  XNOR2_X1 U1233 ( .A(n1552), .B(n1618), .ZN(n893) );
  AOI221_X1 U1234 ( .B1(B[11]), .B2(n1582), .C1(B[10]), .C2(n1581), .A(n1619), 
        .ZN(n1618) );
  OAI22_X1 U1235 ( .A1(n1576), .A2(n1620), .B1(n1586), .B2(n1621), .ZN(n1619)
         );
  XNOR2_X1 U1236 ( .A(n1552), .B(n1622), .ZN(n892) );
  AOI221_X1 U1237 ( .B1(B[12]), .B2(n1582), .C1(B[11]), .C2(n1581), .A(n1623), 
        .ZN(n1622) );
  OAI22_X1 U1238 ( .A1(n1576), .A2(n1624), .B1(n1586), .B2(n1625), .ZN(n1623)
         );
  XNOR2_X1 U1239 ( .A(n1552), .B(n1626), .ZN(n891) );
  AOI221_X1 U1240 ( .B1(B[13]), .B2(n1582), .C1(B[12]), .C2(n1581), .A(n1627), 
        .ZN(n1626) );
  OAI22_X1 U1241 ( .A1(n1576), .A2(n1628), .B1(n1586), .B2(n1629), .ZN(n1627)
         );
  XNOR2_X1 U1242 ( .A(n1552), .B(n1630), .ZN(n890) );
  AOI221_X1 U1243 ( .B1(B[14]), .B2(n1582), .C1(B[13]), .C2(n1581), .A(n1631), 
        .ZN(n1630) );
  OAI22_X1 U1244 ( .A1(n1576), .A2(n1632), .B1(n1586), .B2(n1633), .ZN(n1631)
         );
  XNOR2_X1 U1245 ( .A(n1552), .B(n1634), .ZN(n889) );
  AOI221_X1 U1246 ( .B1(B[15]), .B2(n1582), .C1(B[14]), .C2(n1581), .A(n1635), 
        .ZN(n1634) );
  OAI22_X1 U1247 ( .A1(n1576), .A2(n1636), .B1(n1586), .B2(n1637), .ZN(n1635)
         );
  XNOR2_X1 U1248 ( .A(n1552), .B(n1638), .ZN(n888) );
  AOI221_X1 U1249 ( .B1(B[16]), .B2(n1582), .C1(B[15]), .C2(n1581), .A(n1639), 
        .ZN(n1638) );
  OAI22_X1 U1250 ( .A1(n1576), .A2(n1640), .B1(n1586), .B2(n1641), .ZN(n1639)
         );
  XNOR2_X1 U1251 ( .A(n1552), .B(n1642), .ZN(n887) );
  AOI221_X1 U1252 ( .B1(B[17]), .B2(n1582), .C1(B[16]), .C2(n1581), .A(n1643), 
        .ZN(n1642) );
  OAI22_X1 U1253 ( .A1(n1576), .A2(n1644), .B1(n1586), .B2(n1645), .ZN(n1643)
         );
  XNOR2_X1 U1254 ( .A(n1552), .B(n1646), .ZN(n886) );
  AOI221_X1 U1255 ( .B1(B[18]), .B2(n1582), .C1(B[17]), .C2(n1581), .A(n1647), 
        .ZN(n1646) );
  OAI22_X1 U1256 ( .A1(n1576), .A2(n1648), .B1(n1586), .B2(n1649), .ZN(n1647)
         );
  XNOR2_X1 U1257 ( .A(n1552), .B(n1650), .ZN(n885) );
  AOI221_X1 U1258 ( .B1(B[19]), .B2(n1582), .C1(B[18]), .C2(n1581), .A(n1651), 
        .ZN(n1650) );
  OAI22_X1 U1259 ( .A1(n1576), .A2(n1652), .B1(n1586), .B2(n1653), .ZN(n1651)
         );
  XNOR2_X1 U1260 ( .A(A[5]), .B(n1654), .ZN(n884) );
  AOI221_X1 U1261 ( .B1(n1582), .B2(B[20]), .C1(B[19]), .C2(n1581), .A(n1655), 
        .ZN(n1654) );
  OAI22_X1 U1262 ( .A1(n1576), .A2(n1656), .B1(n1586), .B2(n1657), .ZN(n1655)
         );
  XNOR2_X1 U1263 ( .A(A[5]), .B(n1658), .ZN(n883) );
  AOI221_X1 U1264 ( .B1(n1582), .B2(B[21]), .C1(n1581), .C2(B[20]), .A(n1659), 
        .ZN(n1658) );
  OAI22_X1 U1265 ( .A1(n1576), .A2(n1660), .B1(n1586), .B2(n1661), .ZN(n1659)
         );
  XNOR2_X1 U1266 ( .A(A[5]), .B(n1662), .ZN(n882) );
  AOI221_X1 U1267 ( .B1(n1582), .B2(B[22]), .C1(n1581), .C2(B[21]), .A(n1663), 
        .ZN(n1662) );
  OAI22_X1 U1268 ( .A1(n1562), .A2(n1576), .B1(n1564), .B2(n1586), .ZN(n1663)
         );
  XNOR2_X1 U1269 ( .A(A[5]), .B(n1664), .ZN(n881) );
  AOI221_X1 U1270 ( .B1(n1582), .B2(B[23]), .C1(n1581), .C2(B[22]), .A(n1665), 
        .ZN(n1664) );
  OAI22_X1 U1271 ( .A1(n1567), .A2(n1576), .B1(n1568), .B2(n1586), .ZN(n1665)
         );
  XNOR2_X1 U1272 ( .A(A[5]), .B(n1666), .ZN(n880) );
  AOI221_X1 U1273 ( .B1(n1582), .B2(B[23]), .C1(n1581), .C2(n1554), .A(n1667), 
        .ZN(n1666) );
  OAI22_X1 U1274 ( .A1(n1571), .A2(n1576), .B1(n1572), .B2(n1586), .ZN(n1667)
         );
  XNOR2_X1 U1275 ( .A(n1552), .B(n1668), .ZN(n879) );
  OAI221_X1 U1276 ( .B1(n1556), .B2(n1586), .C1(n1556), .C2(n1576), .A(n1669), 
        .ZN(n1668) );
  OAI21_X1 U1277 ( .B1(n1582), .B2(n1581), .A(n1554), .ZN(n1669) );
  INV_X1 U1278 ( .A(n1673), .ZN(n1670) );
  XNOR2_X1 U1279 ( .A(A[3]), .B(A[4]), .ZN(n1671) );
  XNOR2_X1 U1280 ( .A(A[4]), .B(n1553), .ZN(n1672) );
  XOR2_X1 U1281 ( .A(A[3]), .B(n1674), .Z(n1673) );
  XNOR2_X1 U1282 ( .A(n1675), .B(n1551), .ZN(n878) );
  OAI22_X1 U1283 ( .A1(n1574), .A2(n1676), .B1(n1574), .B2(n1677), .ZN(n1675)
         );
  XNOR2_X1 U1284 ( .A(n1678), .B(n1551), .ZN(n877) );
  OAI222_X1 U1285 ( .A1(n1578), .A2(n1676), .B1(n1574), .B2(n1679), .C1(n1580), 
        .C2(n1677), .ZN(n1678) );
  INV_X1 U1286 ( .A(n1680), .ZN(n1679) );
  INV_X1 U1287 ( .A(n1681), .ZN(n1676) );
  XNOR2_X1 U1288 ( .A(n1550), .B(n1682), .ZN(n876) );
  AOI221_X1 U1289 ( .B1(n1681), .B2(B[2]), .C1(n1680), .C2(B[1]), .A(n1683), 
        .ZN(n1682) );
  OAI22_X1 U1290 ( .A1(n1585), .A2(n1677), .B1(n1574), .B2(n1684), .ZN(n1683)
         );
  XNOR2_X1 U1291 ( .A(n1550), .B(n1685), .ZN(n875) );
  AOI221_X1 U1292 ( .B1(n1681), .B2(B[3]), .C1(n1680), .C2(B[2]), .A(n1686), 
        .ZN(n1685) );
  OAI22_X1 U1293 ( .A1(n1589), .A2(n1677), .B1(n1578), .B2(n1684), .ZN(n1686)
         );
  XNOR2_X1 U1294 ( .A(n1550), .B(n1687), .ZN(n874) );
  AOI221_X1 U1295 ( .B1(n1681), .B2(B[4]), .C1(n1680), .C2(B[3]), .A(n1688), 
        .ZN(n1687) );
  OAI22_X1 U1296 ( .A1(n1592), .A2(n1677), .B1(n1593), .B2(n1684), .ZN(n1688)
         );
  XNOR2_X1 U1297 ( .A(n1550), .B(n1689), .ZN(n873) );
  AOI221_X1 U1298 ( .B1(n1681), .B2(B[5]), .C1(n1680), .C2(B[4]), .A(n1690), 
        .ZN(n1689) );
  OAI22_X1 U1299 ( .A1(n1596), .A2(n1677), .B1(n1597), .B2(n1684), .ZN(n1690)
         );
  XNOR2_X1 U1300 ( .A(n1550), .B(n1691), .ZN(n872) );
  AOI221_X1 U1301 ( .B1(n1681), .B2(B[6]), .C1(n1680), .C2(B[5]), .A(n1692), 
        .ZN(n1691) );
  OAI22_X1 U1302 ( .A1(n1600), .A2(n1677), .B1(n1601), .B2(n1684), .ZN(n1692)
         );
  XNOR2_X1 U1303 ( .A(n1550), .B(n1693), .ZN(n871) );
  AOI221_X1 U1304 ( .B1(n1681), .B2(B[7]), .C1(n1680), .C2(B[6]), .A(n1694), 
        .ZN(n1693) );
  OAI22_X1 U1305 ( .A1(n1604), .A2(n1677), .B1(n1605), .B2(n1684), .ZN(n1694)
         );
  XNOR2_X1 U1306 ( .A(n1550), .B(n1695), .ZN(n870) );
  AOI221_X1 U1307 ( .B1(n1681), .B2(B[8]), .C1(n1680), .C2(B[7]), .A(n1696), 
        .ZN(n1695) );
  OAI22_X1 U1308 ( .A1(n1608), .A2(n1677), .B1(n1609), .B2(n1684), .ZN(n1696)
         );
  XNOR2_X1 U1309 ( .A(n1550), .B(n1697), .ZN(n869) );
  AOI221_X1 U1310 ( .B1(n1681), .B2(B[9]), .C1(n1680), .C2(B[8]), .A(n1698), 
        .ZN(n1697) );
  OAI22_X1 U1311 ( .A1(n1612), .A2(n1677), .B1(n1613), .B2(n1684), .ZN(n1698)
         );
  XNOR2_X1 U1312 ( .A(n1550), .B(n1699), .ZN(n868) );
  AOI221_X1 U1313 ( .B1(n1681), .B2(B[10]), .C1(n1680), .C2(B[9]), .A(n1700), 
        .ZN(n1699) );
  OAI22_X1 U1314 ( .A1(n1616), .A2(n1677), .B1(n1617), .B2(n1684), .ZN(n1700)
         );
  XNOR2_X1 U1315 ( .A(n1550), .B(n1701), .ZN(n867) );
  AOI221_X1 U1316 ( .B1(n1681), .B2(B[11]), .C1(n1680), .C2(B[10]), .A(n1702), 
        .ZN(n1701) );
  OAI22_X1 U1317 ( .A1(n1620), .A2(n1677), .B1(n1621), .B2(n1684), .ZN(n1702)
         );
  XNOR2_X1 U1318 ( .A(n1550), .B(n1703), .ZN(n866) );
  AOI221_X1 U1319 ( .B1(n1681), .B2(B[12]), .C1(n1680), .C2(B[11]), .A(n1704), 
        .ZN(n1703) );
  OAI22_X1 U1320 ( .A1(n1624), .A2(n1677), .B1(n1625), .B2(n1684), .ZN(n1704)
         );
  XNOR2_X1 U1321 ( .A(n1550), .B(n1705), .ZN(n865) );
  AOI221_X1 U1322 ( .B1(n1681), .B2(B[13]), .C1(n1680), .C2(B[12]), .A(n1706), 
        .ZN(n1705) );
  OAI22_X1 U1323 ( .A1(n1628), .A2(n1677), .B1(n1629), .B2(n1684), .ZN(n1706)
         );
  XNOR2_X1 U1324 ( .A(n1550), .B(n1707), .ZN(n864) );
  AOI221_X1 U1325 ( .B1(n1681), .B2(B[14]), .C1(n1680), .C2(B[13]), .A(n1708), 
        .ZN(n1707) );
  OAI22_X1 U1326 ( .A1(n1632), .A2(n1677), .B1(n1633), .B2(n1684), .ZN(n1708)
         );
  XNOR2_X1 U1327 ( .A(n1550), .B(n1709), .ZN(n863) );
  AOI221_X1 U1328 ( .B1(n1681), .B2(B[15]), .C1(n1680), .C2(B[14]), .A(n1710), 
        .ZN(n1709) );
  OAI22_X1 U1329 ( .A1(n1636), .A2(n1677), .B1(n1637), .B2(n1684), .ZN(n1710)
         );
  XNOR2_X1 U1330 ( .A(n1550), .B(n1711), .ZN(n862) );
  AOI221_X1 U1331 ( .B1(n1681), .B2(B[16]), .C1(n1680), .C2(B[15]), .A(n1712), 
        .ZN(n1711) );
  OAI22_X1 U1332 ( .A1(n1640), .A2(n1677), .B1(n1641), .B2(n1684), .ZN(n1712)
         );
  XNOR2_X1 U1333 ( .A(n1550), .B(n1713), .ZN(n861) );
  AOI221_X1 U1334 ( .B1(n1681), .B2(B[17]), .C1(n1680), .C2(B[16]), .A(n1714), 
        .ZN(n1713) );
  OAI22_X1 U1335 ( .A1(n1644), .A2(n1677), .B1(n1645), .B2(n1684), .ZN(n1714)
         );
  XNOR2_X1 U1336 ( .A(n1550), .B(n1715), .ZN(n860) );
  AOI221_X1 U1337 ( .B1(n1681), .B2(B[18]), .C1(n1680), .C2(B[17]), .A(n1716), 
        .ZN(n1715) );
  OAI22_X1 U1338 ( .A1(n1648), .A2(n1677), .B1(n1649), .B2(n1684), .ZN(n1716)
         );
  XNOR2_X1 U1339 ( .A(n1550), .B(n1717), .ZN(n859) );
  AOI221_X1 U1340 ( .B1(n1681), .B2(B[19]), .C1(n1680), .C2(B[18]), .A(n1718), 
        .ZN(n1717) );
  OAI22_X1 U1341 ( .A1(n1652), .A2(n1677), .B1(n1653), .B2(n1684), .ZN(n1718)
         );
  XNOR2_X1 U1342 ( .A(A[8]), .B(n1719), .ZN(n858) );
  AOI221_X1 U1343 ( .B1(n1681), .B2(B[20]), .C1(n1680), .C2(B[19]), .A(n1720), 
        .ZN(n1719) );
  OAI22_X1 U1344 ( .A1(n1656), .A2(n1677), .B1(n1657), .B2(n1684), .ZN(n1720)
         );
  XNOR2_X1 U1345 ( .A(A[8]), .B(n1721), .ZN(n857) );
  AOI221_X1 U1346 ( .B1(n1681), .B2(B[21]), .C1(n1680), .C2(B[20]), .A(n1722), 
        .ZN(n1721) );
  OAI22_X1 U1347 ( .A1(n1660), .A2(n1677), .B1(n1661), .B2(n1684), .ZN(n1722)
         );
  XNOR2_X1 U1348 ( .A(A[8]), .B(n1723), .ZN(n856) );
  AOI221_X1 U1349 ( .B1(n1681), .B2(B[22]), .C1(n1680), .C2(B[21]), .A(n1724), 
        .ZN(n1723) );
  OAI22_X1 U1350 ( .A1(n1562), .A2(n1677), .B1(n1564), .B2(n1684), .ZN(n1724)
         );
  XNOR2_X1 U1351 ( .A(A[8]), .B(n1725), .ZN(n855) );
  AOI221_X1 U1352 ( .B1(n1681), .B2(B[23]), .C1(n1680), .C2(B[22]), .A(n1726), 
        .ZN(n1725) );
  OAI22_X1 U1353 ( .A1(n1567), .A2(n1677), .B1(n1568), .B2(n1684), .ZN(n1726)
         );
  XNOR2_X1 U1354 ( .A(A[8]), .B(n1727), .ZN(n854) );
  AOI221_X1 U1355 ( .B1(n1681), .B2(B[23]), .C1(n1680), .C2(n1554), .A(n1728), 
        .ZN(n1727) );
  OAI22_X1 U1356 ( .A1(n1571), .A2(n1677), .B1(n1572), .B2(n1684), .ZN(n1728)
         );
  XNOR2_X1 U1357 ( .A(n1550), .B(n1729), .ZN(n853) );
  OAI221_X1 U1358 ( .B1(n1555), .B2(n1684), .C1(n1556), .C2(n1677), .A(n1730), 
        .ZN(n1729) );
  OAI21_X1 U1359 ( .B1(n1681), .B2(n1680), .A(n1554), .ZN(n1730) );
  INV_X1 U1360 ( .A(n1734), .ZN(n1731) );
  XNOR2_X1 U1361 ( .A(A[6]), .B(A[7]), .ZN(n1732) );
  XNOR2_X1 U1362 ( .A(A[7]), .B(n1551), .ZN(n1733) );
  XOR2_X1 U1363 ( .A(A[6]), .B(n1553), .Z(n1734) );
  XNOR2_X1 U1364 ( .A(n1735), .B(n1549), .ZN(n852) );
  OAI22_X1 U1365 ( .A1(n1574), .A2(n1736), .B1(n1574), .B2(n1737), .ZN(n1735)
         );
  XNOR2_X1 U1366 ( .A(n1738), .B(n1549), .ZN(n851) );
  OAI222_X1 U1367 ( .A1(n1578), .A2(n1736), .B1(n1574), .B2(n1739), .C1(n1580), 
        .C2(n1737), .ZN(n1738) );
  INV_X1 U1368 ( .A(n1740), .ZN(n1739) );
  INV_X1 U1369 ( .A(n1741), .ZN(n1736) );
  XNOR2_X1 U1370 ( .A(n1548), .B(n1742), .ZN(n850) );
  AOI221_X1 U1371 ( .B1(n1741), .B2(B[2]), .C1(n1740), .C2(B[1]), .A(n1743), 
        .ZN(n1742) );
  OAI22_X1 U1372 ( .A1(n1585), .A2(n1737), .B1(n1574), .B2(n1744), .ZN(n1743)
         );
  XNOR2_X1 U1373 ( .A(n1548), .B(n1745), .ZN(n849) );
  AOI221_X1 U1374 ( .B1(n1741), .B2(B[3]), .C1(n1740), .C2(B[2]), .A(n1746), 
        .ZN(n1745) );
  OAI22_X1 U1375 ( .A1(n1589), .A2(n1737), .B1(n1578), .B2(n1744), .ZN(n1746)
         );
  XNOR2_X1 U1376 ( .A(n1548), .B(n1747), .ZN(n848) );
  AOI221_X1 U1377 ( .B1(n1741), .B2(B[4]), .C1(n1740), .C2(B[3]), .A(n1748), 
        .ZN(n1747) );
  OAI22_X1 U1378 ( .A1(n1592), .A2(n1737), .B1(n1593), .B2(n1744), .ZN(n1748)
         );
  XNOR2_X1 U1379 ( .A(n1548), .B(n1749), .ZN(n847) );
  AOI221_X1 U1380 ( .B1(n1741), .B2(B[5]), .C1(n1740), .C2(B[4]), .A(n1750), 
        .ZN(n1749) );
  OAI22_X1 U1381 ( .A1(n1596), .A2(n1737), .B1(n1597), .B2(n1744), .ZN(n1750)
         );
  XNOR2_X1 U1382 ( .A(n1548), .B(n1751), .ZN(n846) );
  AOI221_X1 U1383 ( .B1(n1741), .B2(B[6]), .C1(n1740), .C2(B[5]), .A(n1752), 
        .ZN(n1751) );
  OAI22_X1 U1384 ( .A1(n1600), .A2(n1737), .B1(n1601), .B2(n1744), .ZN(n1752)
         );
  XNOR2_X1 U1385 ( .A(n1548), .B(n1753), .ZN(n845) );
  AOI221_X1 U1386 ( .B1(n1741), .B2(B[7]), .C1(n1740), .C2(B[6]), .A(n1754), 
        .ZN(n1753) );
  OAI22_X1 U1387 ( .A1(n1604), .A2(n1737), .B1(n1605), .B2(n1744), .ZN(n1754)
         );
  XNOR2_X1 U1388 ( .A(n1548), .B(n1755), .ZN(n844) );
  AOI221_X1 U1389 ( .B1(n1741), .B2(B[8]), .C1(n1740), .C2(B[7]), .A(n1756), 
        .ZN(n1755) );
  OAI22_X1 U1390 ( .A1(n1608), .A2(n1737), .B1(n1609), .B2(n1744), .ZN(n1756)
         );
  XNOR2_X1 U1391 ( .A(n1548), .B(n1757), .ZN(n843) );
  AOI221_X1 U1392 ( .B1(n1741), .B2(B[9]), .C1(n1740), .C2(B[8]), .A(n1758), 
        .ZN(n1757) );
  OAI22_X1 U1393 ( .A1(n1612), .A2(n1737), .B1(n1613), .B2(n1744), .ZN(n1758)
         );
  XNOR2_X1 U1394 ( .A(n1548), .B(n1759), .ZN(n842) );
  AOI221_X1 U1395 ( .B1(n1741), .B2(B[10]), .C1(n1740), .C2(B[9]), .A(n1760), 
        .ZN(n1759) );
  OAI22_X1 U1396 ( .A1(n1616), .A2(n1737), .B1(n1617), .B2(n1744), .ZN(n1760)
         );
  XNOR2_X1 U1397 ( .A(n1548), .B(n1761), .ZN(n841) );
  AOI221_X1 U1398 ( .B1(n1741), .B2(B[11]), .C1(n1740), .C2(B[10]), .A(n1762), 
        .ZN(n1761) );
  OAI22_X1 U1399 ( .A1(n1620), .A2(n1737), .B1(n1621), .B2(n1744), .ZN(n1762)
         );
  XNOR2_X1 U1400 ( .A(n1548), .B(n1763), .ZN(n840) );
  AOI221_X1 U1401 ( .B1(n1741), .B2(B[12]), .C1(n1740), .C2(B[11]), .A(n1764), 
        .ZN(n1763) );
  OAI22_X1 U1402 ( .A1(n1624), .A2(n1737), .B1(n1625), .B2(n1744), .ZN(n1764)
         );
  XNOR2_X1 U1403 ( .A(n1548), .B(n1765), .ZN(n839) );
  AOI221_X1 U1404 ( .B1(n1741), .B2(B[13]), .C1(n1740), .C2(B[12]), .A(n1766), 
        .ZN(n1765) );
  OAI22_X1 U1405 ( .A1(n1628), .A2(n1737), .B1(n1629), .B2(n1744), .ZN(n1766)
         );
  XNOR2_X1 U1406 ( .A(n1548), .B(n1767), .ZN(n838) );
  AOI221_X1 U1407 ( .B1(n1741), .B2(B[14]), .C1(n1740), .C2(B[13]), .A(n1768), 
        .ZN(n1767) );
  OAI22_X1 U1408 ( .A1(n1632), .A2(n1737), .B1(n1633), .B2(n1744), .ZN(n1768)
         );
  XNOR2_X1 U1409 ( .A(n1548), .B(n1769), .ZN(n837) );
  AOI221_X1 U1410 ( .B1(n1741), .B2(B[15]), .C1(n1740), .C2(B[14]), .A(n1770), 
        .ZN(n1769) );
  OAI22_X1 U1411 ( .A1(n1636), .A2(n1737), .B1(n1637), .B2(n1744), .ZN(n1770)
         );
  XNOR2_X1 U1412 ( .A(n1548), .B(n1771), .ZN(n836) );
  AOI221_X1 U1413 ( .B1(n1741), .B2(B[16]), .C1(n1740), .C2(B[15]), .A(n1772), 
        .ZN(n1771) );
  OAI22_X1 U1414 ( .A1(n1640), .A2(n1737), .B1(n1641), .B2(n1744), .ZN(n1772)
         );
  XNOR2_X1 U1415 ( .A(n1548), .B(n1773), .ZN(n835) );
  AOI221_X1 U1416 ( .B1(n1741), .B2(B[17]), .C1(n1740), .C2(B[16]), .A(n1774), 
        .ZN(n1773) );
  OAI22_X1 U1417 ( .A1(n1644), .A2(n1737), .B1(n1645), .B2(n1744), .ZN(n1774)
         );
  XNOR2_X1 U1418 ( .A(n1548), .B(n1775), .ZN(n834) );
  AOI221_X1 U1419 ( .B1(n1741), .B2(B[18]), .C1(n1740), .C2(B[17]), .A(n1776), 
        .ZN(n1775) );
  OAI22_X1 U1420 ( .A1(n1648), .A2(n1737), .B1(n1649), .B2(n1744), .ZN(n1776)
         );
  XNOR2_X1 U1421 ( .A(n1548), .B(n1777), .ZN(n833) );
  AOI221_X1 U1422 ( .B1(n1741), .B2(B[19]), .C1(n1740), .C2(B[18]), .A(n1778), 
        .ZN(n1777) );
  OAI22_X1 U1423 ( .A1(n1652), .A2(n1737), .B1(n1653), .B2(n1744), .ZN(n1778)
         );
  XNOR2_X1 U1424 ( .A(n1548), .B(n1779), .ZN(n832) );
  AOI221_X1 U1425 ( .B1(n1741), .B2(B[20]), .C1(n1740), .C2(B[19]), .A(n1780), 
        .ZN(n1779) );
  OAI22_X1 U1426 ( .A1(n1656), .A2(n1737), .B1(n1657), .B2(n1744), .ZN(n1780)
         );
  XNOR2_X1 U1427 ( .A(A[11]), .B(n1781), .ZN(n831) );
  AOI221_X1 U1428 ( .B1(n1741), .B2(B[21]), .C1(n1740), .C2(B[20]), .A(n1782), 
        .ZN(n1781) );
  OAI22_X1 U1429 ( .A1(n1660), .A2(n1737), .B1(n1661), .B2(n1744), .ZN(n1782)
         );
  XNOR2_X1 U1430 ( .A(A[11]), .B(n1783), .ZN(n830) );
  AOI221_X1 U1431 ( .B1(n1741), .B2(B[22]), .C1(n1740), .C2(B[21]), .A(n1784), 
        .ZN(n1783) );
  OAI22_X1 U1432 ( .A1(n1562), .A2(n1737), .B1(n1564), .B2(n1744), .ZN(n1784)
         );
  XNOR2_X1 U1433 ( .A(A[11]), .B(n1785), .ZN(n829) );
  AOI221_X1 U1434 ( .B1(n1741), .B2(B[23]), .C1(n1740), .C2(B[22]), .A(n1786), 
        .ZN(n1785) );
  OAI22_X1 U1435 ( .A1(n1567), .A2(n1737), .B1(n1568), .B2(n1744), .ZN(n1786)
         );
  XNOR2_X1 U1436 ( .A(A[11]), .B(n1787), .ZN(n828) );
  AOI221_X1 U1437 ( .B1(n1741), .B2(B[23]), .C1(n1740), .C2(n1554), .A(n1788), 
        .ZN(n1787) );
  OAI22_X1 U1438 ( .A1(n1571), .A2(n1737), .B1(n1572), .B2(n1744), .ZN(n1788)
         );
  XNOR2_X1 U1439 ( .A(A[11]), .B(n1789), .ZN(n827) );
  OAI221_X1 U1440 ( .B1(n1556), .B2(n1744), .C1(n1556), .C2(n1737), .A(n1790), 
        .ZN(n1789) );
  OAI21_X1 U1441 ( .B1(n1741), .B2(n1740), .A(n1554), .ZN(n1790) );
  INV_X1 U1442 ( .A(n1794), .ZN(n1791) );
  XNOR2_X1 U1443 ( .A(A[10]), .B(A[9]), .ZN(n1792) );
  XNOR2_X1 U1444 ( .A(A[10]), .B(n1549), .ZN(n1793) );
  XOR2_X1 U1445 ( .A(A[9]), .B(n1551), .Z(n1794) );
  XNOR2_X1 U1446 ( .A(n1795), .B(n1547), .ZN(n826) );
  OAI22_X1 U1447 ( .A1(n1574), .A2(n1796), .B1(n1574), .B2(n1797), .ZN(n1795)
         );
  XNOR2_X1 U1448 ( .A(n1798), .B(n1547), .ZN(n825) );
  OAI222_X1 U1449 ( .A1(n1578), .A2(n1796), .B1(n1574), .B2(n1799), .C1(n1580), 
        .C2(n1797), .ZN(n1798) );
  INV_X1 U1450 ( .A(n1800), .ZN(n1799) );
  INV_X1 U1451 ( .A(n1801), .ZN(n1796) );
  XNOR2_X1 U1452 ( .A(n1546), .B(n1802), .ZN(n824) );
  AOI221_X1 U1453 ( .B1(n1801), .B2(B[2]), .C1(n1800), .C2(B[1]), .A(n1803), 
        .ZN(n1802) );
  OAI22_X1 U1454 ( .A1(n1585), .A2(n1797), .B1(n1574), .B2(n1804), .ZN(n1803)
         );
  XNOR2_X1 U1455 ( .A(n1546), .B(n1805), .ZN(n823) );
  AOI221_X1 U1456 ( .B1(n1801), .B2(B[3]), .C1(n1800), .C2(B[2]), .A(n1806), 
        .ZN(n1805) );
  OAI22_X1 U1457 ( .A1(n1589), .A2(n1797), .B1(n1578), .B2(n1804), .ZN(n1806)
         );
  XNOR2_X1 U1458 ( .A(n1546), .B(n1807), .ZN(n822) );
  AOI221_X1 U1459 ( .B1(n1801), .B2(B[4]), .C1(n1800), .C2(B[3]), .A(n1808), 
        .ZN(n1807) );
  OAI22_X1 U1460 ( .A1(n1592), .A2(n1797), .B1(n1593), .B2(n1804), .ZN(n1808)
         );
  XNOR2_X1 U1461 ( .A(n1546), .B(n1809), .ZN(n821) );
  AOI221_X1 U1462 ( .B1(n1801), .B2(B[5]), .C1(n1800), .C2(B[4]), .A(n1810), 
        .ZN(n1809) );
  OAI22_X1 U1463 ( .A1(n1596), .A2(n1797), .B1(n1597), .B2(n1804), .ZN(n1810)
         );
  XNOR2_X1 U1464 ( .A(n1546), .B(n1811), .ZN(n820) );
  AOI221_X1 U1465 ( .B1(n1801), .B2(B[6]), .C1(n1800), .C2(B[5]), .A(n1812), 
        .ZN(n1811) );
  OAI22_X1 U1466 ( .A1(n1600), .A2(n1797), .B1(n1601), .B2(n1804), .ZN(n1812)
         );
  XNOR2_X1 U1467 ( .A(n1546), .B(n1813), .ZN(n819) );
  AOI221_X1 U1468 ( .B1(n1801), .B2(B[7]), .C1(n1800), .C2(B[6]), .A(n1814), 
        .ZN(n1813) );
  OAI22_X1 U1469 ( .A1(n1604), .A2(n1797), .B1(n1605), .B2(n1804), .ZN(n1814)
         );
  XNOR2_X1 U1470 ( .A(n1546), .B(n1815), .ZN(n818) );
  AOI221_X1 U1471 ( .B1(n1801), .B2(B[8]), .C1(n1800), .C2(B[7]), .A(n1816), 
        .ZN(n1815) );
  OAI22_X1 U1472 ( .A1(n1608), .A2(n1797), .B1(n1609), .B2(n1804), .ZN(n1816)
         );
  XNOR2_X1 U1473 ( .A(n1546), .B(n1817), .ZN(n817) );
  AOI221_X1 U1474 ( .B1(n1801), .B2(B[9]), .C1(n1800), .C2(B[8]), .A(n1818), 
        .ZN(n1817) );
  OAI22_X1 U1475 ( .A1(n1612), .A2(n1797), .B1(n1613), .B2(n1804), .ZN(n1818)
         );
  XNOR2_X1 U1476 ( .A(n1546), .B(n1819), .ZN(n816) );
  AOI221_X1 U1477 ( .B1(n1801), .B2(B[10]), .C1(n1800), .C2(B[9]), .A(n1820), 
        .ZN(n1819) );
  OAI22_X1 U1478 ( .A1(n1616), .A2(n1797), .B1(n1617), .B2(n1804), .ZN(n1820)
         );
  XNOR2_X1 U1479 ( .A(n1546), .B(n1821), .ZN(n815) );
  AOI221_X1 U1480 ( .B1(n1801), .B2(B[11]), .C1(n1800), .C2(B[10]), .A(n1822), 
        .ZN(n1821) );
  OAI22_X1 U1481 ( .A1(n1620), .A2(n1797), .B1(n1621), .B2(n1804), .ZN(n1822)
         );
  XNOR2_X1 U1482 ( .A(n1546), .B(n1823), .ZN(n814) );
  AOI221_X1 U1483 ( .B1(n1801), .B2(B[12]), .C1(n1800), .C2(B[11]), .A(n1824), 
        .ZN(n1823) );
  OAI22_X1 U1484 ( .A1(n1624), .A2(n1797), .B1(n1625), .B2(n1804), .ZN(n1824)
         );
  XNOR2_X1 U1485 ( .A(n1546), .B(n1825), .ZN(n813) );
  AOI221_X1 U1486 ( .B1(n1801), .B2(B[13]), .C1(n1800), .C2(B[12]), .A(n1826), 
        .ZN(n1825) );
  OAI22_X1 U1487 ( .A1(n1628), .A2(n1797), .B1(n1629), .B2(n1804), .ZN(n1826)
         );
  XNOR2_X1 U1488 ( .A(n1546), .B(n1827), .ZN(n812) );
  AOI221_X1 U1489 ( .B1(n1801), .B2(B[14]), .C1(n1800), .C2(B[13]), .A(n1828), 
        .ZN(n1827) );
  OAI22_X1 U1490 ( .A1(n1632), .A2(n1797), .B1(n1633), .B2(n1804), .ZN(n1828)
         );
  XNOR2_X1 U1491 ( .A(n1546), .B(n1829), .ZN(n811) );
  AOI221_X1 U1492 ( .B1(n1801), .B2(B[15]), .C1(n1800), .C2(B[14]), .A(n1830), 
        .ZN(n1829) );
  OAI22_X1 U1493 ( .A1(n1636), .A2(n1797), .B1(n1637), .B2(n1804), .ZN(n1830)
         );
  XNOR2_X1 U1494 ( .A(n1546), .B(n1831), .ZN(n810) );
  AOI221_X1 U1495 ( .B1(n1801), .B2(B[16]), .C1(n1800), .C2(B[15]), .A(n1832), 
        .ZN(n1831) );
  OAI22_X1 U1496 ( .A1(n1640), .A2(n1797), .B1(n1641), .B2(n1804), .ZN(n1832)
         );
  XNOR2_X1 U1497 ( .A(n1546), .B(n1833), .ZN(n809) );
  AOI221_X1 U1498 ( .B1(n1801), .B2(B[17]), .C1(n1800), .C2(B[16]), .A(n1834), 
        .ZN(n1833) );
  OAI22_X1 U1499 ( .A1(n1644), .A2(n1797), .B1(n1645), .B2(n1804), .ZN(n1834)
         );
  XNOR2_X1 U1500 ( .A(n1546), .B(n1835), .ZN(n808) );
  AOI221_X1 U1501 ( .B1(n1801), .B2(B[18]), .C1(n1800), .C2(B[17]), .A(n1836), 
        .ZN(n1835) );
  OAI22_X1 U1502 ( .A1(n1648), .A2(n1797), .B1(n1649), .B2(n1804), .ZN(n1836)
         );
  XNOR2_X1 U1503 ( .A(n1546), .B(n1837), .ZN(n807) );
  AOI221_X1 U1504 ( .B1(n1801), .B2(B[19]), .C1(n1800), .C2(B[18]), .A(n1838), 
        .ZN(n1837) );
  OAI22_X1 U1505 ( .A1(n1652), .A2(n1797), .B1(n1653), .B2(n1804), .ZN(n1838)
         );
  XNOR2_X1 U1506 ( .A(n1546), .B(n1839), .ZN(n806) );
  AOI221_X1 U1507 ( .B1(n1801), .B2(B[20]), .C1(n1800), .C2(B[19]), .A(n1840), 
        .ZN(n1839) );
  OAI22_X1 U1508 ( .A1(n1656), .A2(n1797), .B1(n1657), .B2(n1804), .ZN(n1840)
         );
  XNOR2_X1 U1509 ( .A(A[14]), .B(n1841), .ZN(n805) );
  AOI221_X1 U1510 ( .B1(n1801), .B2(B[21]), .C1(n1800), .C2(B[20]), .A(n1842), 
        .ZN(n1841) );
  OAI22_X1 U1511 ( .A1(n1660), .A2(n1797), .B1(n1661), .B2(n1804), .ZN(n1842)
         );
  XNOR2_X1 U1512 ( .A(A[14]), .B(n1843), .ZN(n804) );
  AOI221_X1 U1513 ( .B1(n1801), .B2(B[22]), .C1(n1800), .C2(B[21]), .A(n1844), 
        .ZN(n1843) );
  OAI22_X1 U1514 ( .A1(n1562), .A2(n1797), .B1(n1564), .B2(n1804), .ZN(n1844)
         );
  XNOR2_X1 U1515 ( .A(A[14]), .B(n1845), .ZN(n803) );
  AOI221_X1 U1516 ( .B1(n1801), .B2(B[23]), .C1(n1800), .C2(B[22]), .A(n1846), 
        .ZN(n1845) );
  OAI22_X1 U1517 ( .A1(n1567), .A2(n1797), .B1(n1568), .B2(n1804), .ZN(n1846)
         );
  XNOR2_X1 U1518 ( .A(A[14]), .B(n1847), .ZN(n802) );
  AOI221_X1 U1519 ( .B1(n1801), .B2(B[23]), .C1(n1800), .C2(n1554), .A(n1848), 
        .ZN(n1847) );
  OAI22_X1 U1520 ( .A1(n1571), .A2(n1797), .B1(n1572), .B2(n1804), .ZN(n1848)
         );
  XNOR2_X1 U1521 ( .A(A[14]), .B(n1849), .ZN(n801) );
  OAI221_X1 U1522 ( .B1(n1556), .B2(n1804), .C1(n1556), .C2(n1797), .A(n1850), 
        .ZN(n1849) );
  OAI21_X1 U1523 ( .B1(n1801), .B2(n1800), .A(n1554), .ZN(n1850) );
  INV_X1 U1524 ( .A(n1854), .ZN(n1851) );
  XNOR2_X1 U1525 ( .A(A[12]), .B(A[13]), .ZN(n1852) );
  XNOR2_X1 U1526 ( .A(A[13]), .B(n1547), .ZN(n1853) );
  XOR2_X1 U1527 ( .A(A[12]), .B(n1549), .Z(n1854) );
  XNOR2_X1 U1528 ( .A(n1855), .B(n1545), .ZN(n800) );
  OAI22_X1 U1529 ( .A1(n1574), .A2(n1856), .B1(n1574), .B2(n1857), .ZN(n1855)
         );
  XNOR2_X1 U1530 ( .A(n1858), .B(n1545), .ZN(n799) );
  OAI222_X1 U1531 ( .A1(n1578), .A2(n1856), .B1(n1574), .B2(n1859), .C1(n1580), 
        .C2(n1857), .ZN(n1858) );
  INV_X1 U1532 ( .A(n1860), .ZN(n1859) );
  INV_X1 U1533 ( .A(n1861), .ZN(n1856) );
  XNOR2_X1 U1534 ( .A(n1544), .B(n1862), .ZN(n798) );
  AOI221_X1 U1535 ( .B1(n1861), .B2(B[2]), .C1(n1860), .C2(B[1]), .A(n1863), 
        .ZN(n1862) );
  OAI22_X1 U1536 ( .A1(n1585), .A2(n1857), .B1(n1574), .B2(n1864), .ZN(n1863)
         );
  XNOR2_X1 U1537 ( .A(n1544), .B(n1865), .ZN(n797) );
  AOI221_X1 U1538 ( .B1(n1861), .B2(B[3]), .C1(n1860), .C2(B[2]), .A(n1866), 
        .ZN(n1865) );
  OAI22_X1 U1539 ( .A1(n1589), .A2(n1857), .B1(n1578), .B2(n1864), .ZN(n1866)
         );
  XNOR2_X1 U1540 ( .A(n1544), .B(n1867), .ZN(n796) );
  AOI221_X1 U1541 ( .B1(n1861), .B2(B[4]), .C1(n1860), .C2(B[3]), .A(n1868), 
        .ZN(n1867) );
  OAI22_X1 U1542 ( .A1(n1592), .A2(n1857), .B1(n1593), .B2(n1864), .ZN(n1868)
         );
  XNOR2_X1 U1543 ( .A(n1544), .B(n1869), .ZN(n795) );
  AOI221_X1 U1544 ( .B1(n1861), .B2(B[5]), .C1(n1860), .C2(B[4]), .A(n1870), 
        .ZN(n1869) );
  OAI22_X1 U1545 ( .A1(n1596), .A2(n1857), .B1(n1597), .B2(n1864), .ZN(n1870)
         );
  XNOR2_X1 U1546 ( .A(n1544), .B(n1871), .ZN(n794) );
  AOI221_X1 U1547 ( .B1(n1861), .B2(B[6]), .C1(n1860), .C2(B[5]), .A(n1872), 
        .ZN(n1871) );
  OAI22_X1 U1548 ( .A1(n1600), .A2(n1857), .B1(n1601), .B2(n1864), .ZN(n1872)
         );
  XNOR2_X1 U1549 ( .A(n1544), .B(n1873), .ZN(n793) );
  AOI221_X1 U1550 ( .B1(n1861), .B2(B[7]), .C1(n1860), .C2(B[6]), .A(n1874), 
        .ZN(n1873) );
  OAI22_X1 U1551 ( .A1(n1604), .A2(n1857), .B1(n1605), .B2(n1864), .ZN(n1874)
         );
  XNOR2_X1 U1552 ( .A(n1544), .B(n1875), .ZN(n792) );
  AOI221_X1 U1553 ( .B1(n1861), .B2(B[8]), .C1(n1860), .C2(B[7]), .A(n1876), 
        .ZN(n1875) );
  OAI22_X1 U1554 ( .A1(n1608), .A2(n1857), .B1(n1609), .B2(n1864), .ZN(n1876)
         );
  XNOR2_X1 U1555 ( .A(n1544), .B(n1877), .ZN(n791) );
  AOI221_X1 U1556 ( .B1(n1861), .B2(B[9]), .C1(n1860), .C2(B[8]), .A(n1878), 
        .ZN(n1877) );
  OAI22_X1 U1557 ( .A1(n1612), .A2(n1857), .B1(n1613), .B2(n1864), .ZN(n1878)
         );
  XNOR2_X1 U1558 ( .A(n1544), .B(n1879), .ZN(n790) );
  AOI221_X1 U1559 ( .B1(n1861), .B2(B[10]), .C1(n1860), .C2(B[9]), .A(n1880), 
        .ZN(n1879) );
  OAI22_X1 U1560 ( .A1(n1616), .A2(n1857), .B1(n1617), .B2(n1864), .ZN(n1880)
         );
  XNOR2_X1 U1561 ( .A(n1544), .B(n1881), .ZN(n789) );
  AOI221_X1 U1562 ( .B1(n1861), .B2(B[11]), .C1(n1860), .C2(B[10]), .A(n1882), 
        .ZN(n1881) );
  OAI22_X1 U1563 ( .A1(n1620), .A2(n1857), .B1(n1621), .B2(n1864), .ZN(n1882)
         );
  XNOR2_X1 U1564 ( .A(n1544), .B(n1883), .ZN(n788) );
  AOI221_X1 U1565 ( .B1(n1861), .B2(B[12]), .C1(n1860), .C2(B[11]), .A(n1884), 
        .ZN(n1883) );
  OAI22_X1 U1566 ( .A1(n1624), .A2(n1857), .B1(n1625), .B2(n1864), .ZN(n1884)
         );
  XNOR2_X1 U1567 ( .A(n1544), .B(n1885), .ZN(n787) );
  AOI221_X1 U1568 ( .B1(n1861), .B2(B[13]), .C1(n1860), .C2(B[12]), .A(n1886), 
        .ZN(n1885) );
  OAI22_X1 U1569 ( .A1(n1628), .A2(n1857), .B1(n1629), .B2(n1864), .ZN(n1886)
         );
  XNOR2_X1 U1570 ( .A(n1544), .B(n1887), .ZN(n786) );
  AOI221_X1 U1571 ( .B1(n1861), .B2(B[14]), .C1(n1860), .C2(B[13]), .A(n1888), 
        .ZN(n1887) );
  OAI22_X1 U1572 ( .A1(n1632), .A2(n1857), .B1(n1633), .B2(n1864), .ZN(n1888)
         );
  XNOR2_X1 U1573 ( .A(n1544), .B(n1889), .ZN(n785) );
  AOI221_X1 U1574 ( .B1(n1861), .B2(B[15]), .C1(n1860), .C2(B[14]), .A(n1890), 
        .ZN(n1889) );
  OAI22_X1 U1575 ( .A1(n1636), .A2(n1857), .B1(n1637), .B2(n1864), .ZN(n1890)
         );
  XNOR2_X1 U1576 ( .A(n1544), .B(n1891), .ZN(n784) );
  AOI221_X1 U1577 ( .B1(n1861), .B2(B[16]), .C1(n1860), .C2(B[15]), .A(n1892), 
        .ZN(n1891) );
  OAI22_X1 U1578 ( .A1(n1640), .A2(n1857), .B1(n1641), .B2(n1864), .ZN(n1892)
         );
  XNOR2_X1 U1579 ( .A(n1544), .B(n1893), .ZN(n783) );
  AOI221_X1 U1580 ( .B1(n1861), .B2(B[17]), .C1(n1860), .C2(B[16]), .A(n1894), 
        .ZN(n1893) );
  OAI22_X1 U1581 ( .A1(n1644), .A2(n1857), .B1(n1645), .B2(n1864), .ZN(n1894)
         );
  XNOR2_X1 U1582 ( .A(n1544), .B(n1895), .ZN(n782) );
  AOI221_X1 U1583 ( .B1(n1861), .B2(B[18]), .C1(n1860), .C2(B[17]), .A(n1896), 
        .ZN(n1895) );
  OAI22_X1 U1584 ( .A1(n1648), .A2(n1857), .B1(n1649), .B2(n1864), .ZN(n1896)
         );
  XNOR2_X1 U1585 ( .A(n1544), .B(n1897), .ZN(n781) );
  AOI221_X1 U1586 ( .B1(n1861), .B2(B[19]), .C1(n1860), .C2(B[18]), .A(n1898), 
        .ZN(n1897) );
  OAI22_X1 U1587 ( .A1(n1652), .A2(n1857), .B1(n1653), .B2(n1864), .ZN(n1898)
         );
  XNOR2_X1 U1588 ( .A(n1544), .B(n1899), .ZN(n780) );
  AOI221_X1 U1589 ( .B1(n1861), .B2(B[20]), .C1(n1860), .C2(B[19]), .A(n1900), 
        .ZN(n1899) );
  OAI22_X1 U1590 ( .A1(n1656), .A2(n1857), .B1(n1657), .B2(n1864), .ZN(n1900)
         );
  XNOR2_X1 U1591 ( .A(A[17]), .B(n1901), .ZN(n779) );
  AOI221_X1 U1592 ( .B1(n1861), .B2(B[21]), .C1(n1860), .C2(B[20]), .A(n1902), 
        .ZN(n1901) );
  OAI22_X1 U1593 ( .A1(n1660), .A2(n1857), .B1(n1661), .B2(n1864), .ZN(n1902)
         );
  XNOR2_X1 U1594 ( .A(A[17]), .B(n1903), .ZN(n778) );
  AOI221_X1 U1595 ( .B1(n1861), .B2(B[22]), .C1(n1860), .C2(B[21]), .A(n1904), 
        .ZN(n1903) );
  OAI22_X1 U1596 ( .A1(n1562), .A2(n1857), .B1(n1564), .B2(n1864), .ZN(n1904)
         );
  XNOR2_X1 U1597 ( .A(A[17]), .B(n1905), .ZN(n777) );
  AOI221_X1 U1598 ( .B1(n1861), .B2(B[23]), .C1(n1860), .C2(B[22]), .A(n1906), 
        .ZN(n1905) );
  OAI22_X1 U1599 ( .A1(n1567), .A2(n1857), .B1(n1568), .B2(n1864), .ZN(n1906)
         );
  XNOR2_X1 U1600 ( .A(A[17]), .B(n1907), .ZN(n776) );
  AOI221_X1 U1601 ( .B1(n1861), .B2(B[23]), .C1(n1860), .C2(n1554), .A(n1908), 
        .ZN(n1907) );
  OAI22_X1 U1602 ( .A1(n1571), .A2(n1857), .B1(n1572), .B2(n1864), .ZN(n1908)
         );
  XNOR2_X1 U1603 ( .A(A[17]), .B(n1909), .ZN(n775) );
  OAI221_X1 U1604 ( .B1(n1556), .B2(n1864), .C1(n1556), .C2(n1857), .A(n1910), 
        .ZN(n1909) );
  OAI21_X1 U1605 ( .B1(n1861), .B2(n1860), .A(n1554), .ZN(n1910) );
  INV_X1 U1606 ( .A(n1914), .ZN(n1911) );
  XNOR2_X1 U1607 ( .A(A[15]), .B(A[16]), .ZN(n1912) );
  XNOR2_X1 U1608 ( .A(A[16]), .B(n1545), .ZN(n1913) );
  XOR2_X1 U1609 ( .A(A[15]), .B(n1547), .Z(n1914) );
  XNOR2_X1 U1610 ( .A(n1915), .B(n1543), .ZN(n774) );
  OAI22_X1 U1611 ( .A1(n1574), .A2(n1916), .B1(n1574), .B2(n1917), .ZN(n1915)
         );
  XNOR2_X1 U1612 ( .A(n1918), .B(n1543), .ZN(n773) );
  OAI222_X1 U1613 ( .A1(n1578), .A2(n1916), .B1(n1574), .B2(n1919), .C1(n1580), 
        .C2(n1917), .ZN(n1918) );
  INV_X1 U1614 ( .A(n1920), .ZN(n1919) );
  INV_X1 U1615 ( .A(n1921), .ZN(n1916) );
  XNOR2_X1 U1616 ( .A(n1542), .B(n1922), .ZN(n772) );
  AOI221_X1 U1617 ( .B1(n1921), .B2(B[2]), .C1(n1920), .C2(B[1]), .A(n1923), 
        .ZN(n1922) );
  OAI22_X1 U1618 ( .A1(n1585), .A2(n1917), .B1(n1574), .B2(n1924), .ZN(n1923)
         );
  XNOR2_X1 U1619 ( .A(n1542), .B(n1925), .ZN(n771) );
  AOI221_X1 U1620 ( .B1(n1921), .B2(B[3]), .C1(n1920), .C2(B[2]), .A(n1926), 
        .ZN(n1925) );
  OAI22_X1 U1621 ( .A1(n1589), .A2(n1917), .B1(n1578), .B2(n1924), .ZN(n1926)
         );
  XNOR2_X1 U1622 ( .A(n1542), .B(n1927), .ZN(n770) );
  AOI221_X1 U1623 ( .B1(n1921), .B2(B[4]), .C1(n1920), .C2(B[3]), .A(n1928), 
        .ZN(n1927) );
  OAI22_X1 U1624 ( .A1(n1592), .A2(n1917), .B1(n1593), .B2(n1924), .ZN(n1928)
         );
  XNOR2_X1 U1625 ( .A(n1542), .B(n1929), .ZN(n769) );
  AOI221_X1 U1626 ( .B1(n1921), .B2(B[5]), .C1(n1920), .C2(B[4]), .A(n1930), 
        .ZN(n1929) );
  OAI22_X1 U1627 ( .A1(n1596), .A2(n1917), .B1(n1597), .B2(n1924), .ZN(n1930)
         );
  XNOR2_X1 U1628 ( .A(n1542), .B(n1931), .ZN(n768) );
  AOI221_X1 U1629 ( .B1(n1921), .B2(B[6]), .C1(n1920), .C2(B[5]), .A(n1932), 
        .ZN(n1931) );
  OAI22_X1 U1630 ( .A1(n1600), .A2(n1917), .B1(n1601), .B2(n1924), .ZN(n1932)
         );
  XNOR2_X1 U1631 ( .A(n1542), .B(n1933), .ZN(n767) );
  AOI221_X1 U1632 ( .B1(n1921), .B2(B[7]), .C1(n1920), .C2(B[6]), .A(n1934), 
        .ZN(n1933) );
  OAI22_X1 U1633 ( .A1(n1604), .A2(n1917), .B1(n1605), .B2(n1924), .ZN(n1934)
         );
  XNOR2_X1 U1634 ( .A(n1542), .B(n1935), .ZN(n766) );
  AOI221_X1 U1635 ( .B1(n1921), .B2(B[8]), .C1(n1920), .C2(B[7]), .A(n1936), 
        .ZN(n1935) );
  OAI22_X1 U1636 ( .A1(n1608), .A2(n1917), .B1(n1609), .B2(n1924), .ZN(n1936)
         );
  XNOR2_X1 U1637 ( .A(n1542), .B(n1937), .ZN(n765) );
  AOI221_X1 U1638 ( .B1(n1921), .B2(B[9]), .C1(n1920), .C2(B[8]), .A(n1938), 
        .ZN(n1937) );
  OAI22_X1 U1639 ( .A1(n1612), .A2(n1917), .B1(n1613), .B2(n1924), .ZN(n1938)
         );
  XNOR2_X1 U1640 ( .A(n1542), .B(n1939), .ZN(n764) );
  AOI221_X1 U1641 ( .B1(n1921), .B2(B[10]), .C1(n1920), .C2(B[9]), .A(n1940), 
        .ZN(n1939) );
  OAI22_X1 U1642 ( .A1(n1616), .A2(n1917), .B1(n1617), .B2(n1924), .ZN(n1940)
         );
  XNOR2_X1 U1643 ( .A(n1542), .B(n1941), .ZN(n763) );
  AOI221_X1 U1644 ( .B1(n1921), .B2(B[11]), .C1(n1920), .C2(B[10]), .A(n1942), 
        .ZN(n1941) );
  OAI22_X1 U1645 ( .A1(n1620), .A2(n1917), .B1(n1621), .B2(n1924), .ZN(n1942)
         );
  XNOR2_X1 U1646 ( .A(n1542), .B(n1943), .ZN(n762) );
  AOI221_X1 U1647 ( .B1(n1921), .B2(B[12]), .C1(n1920), .C2(B[11]), .A(n1944), 
        .ZN(n1943) );
  OAI22_X1 U1648 ( .A1(n1624), .A2(n1917), .B1(n1625), .B2(n1924), .ZN(n1944)
         );
  XNOR2_X1 U1649 ( .A(n1542), .B(n1945), .ZN(n761) );
  AOI221_X1 U1650 ( .B1(n1921), .B2(B[13]), .C1(n1920), .C2(B[12]), .A(n1946), 
        .ZN(n1945) );
  OAI22_X1 U1651 ( .A1(n1628), .A2(n1917), .B1(n1629), .B2(n1924), .ZN(n1946)
         );
  XNOR2_X1 U1652 ( .A(n1542), .B(n1947), .ZN(n760) );
  AOI221_X1 U1653 ( .B1(n1921), .B2(B[14]), .C1(n1920), .C2(B[13]), .A(n1948), 
        .ZN(n1947) );
  OAI22_X1 U1654 ( .A1(n1632), .A2(n1917), .B1(n1633), .B2(n1924), .ZN(n1948)
         );
  XNOR2_X1 U1655 ( .A(n1542), .B(n1949), .ZN(n759) );
  AOI221_X1 U1656 ( .B1(n1921), .B2(B[15]), .C1(n1920), .C2(B[14]), .A(n1950), 
        .ZN(n1949) );
  OAI22_X1 U1657 ( .A1(n1636), .A2(n1917), .B1(n1637), .B2(n1924), .ZN(n1950)
         );
  XNOR2_X1 U1658 ( .A(n1542), .B(n1951), .ZN(n758) );
  AOI221_X1 U1659 ( .B1(n1921), .B2(B[16]), .C1(n1920), .C2(B[15]), .A(n1952), 
        .ZN(n1951) );
  OAI22_X1 U1660 ( .A1(n1640), .A2(n1917), .B1(n1641), .B2(n1924), .ZN(n1952)
         );
  XNOR2_X1 U1661 ( .A(n1542), .B(n1953), .ZN(n757) );
  AOI221_X1 U1662 ( .B1(n1921), .B2(B[17]), .C1(n1920), .C2(B[16]), .A(n1954), 
        .ZN(n1953) );
  OAI22_X1 U1663 ( .A1(n1644), .A2(n1917), .B1(n1645), .B2(n1924), .ZN(n1954)
         );
  XNOR2_X1 U1664 ( .A(n1542), .B(n1955), .ZN(n756) );
  AOI221_X1 U1665 ( .B1(n1921), .B2(B[18]), .C1(n1920), .C2(B[17]), .A(n1956), 
        .ZN(n1955) );
  OAI22_X1 U1666 ( .A1(n1648), .A2(n1917), .B1(n1649), .B2(n1924), .ZN(n1956)
         );
  XNOR2_X1 U1667 ( .A(n1542), .B(n1957), .ZN(n755) );
  AOI221_X1 U1668 ( .B1(n1921), .B2(B[19]), .C1(n1920), .C2(B[18]), .A(n1958), 
        .ZN(n1957) );
  OAI22_X1 U1669 ( .A1(n1652), .A2(n1917), .B1(n1653), .B2(n1924), .ZN(n1958)
         );
  XNOR2_X1 U1670 ( .A(n1542), .B(n1959), .ZN(n754) );
  AOI221_X1 U1671 ( .B1(n1921), .B2(B[20]), .C1(n1920), .C2(B[19]), .A(n1960), 
        .ZN(n1959) );
  OAI22_X1 U1672 ( .A1(n1656), .A2(n1917), .B1(n1657), .B2(n1924), .ZN(n1960)
         );
  XNOR2_X1 U1673 ( .A(A[20]), .B(n1961), .ZN(n753) );
  AOI221_X1 U1674 ( .B1(n1921), .B2(B[21]), .C1(n1920), .C2(B[20]), .A(n1962), 
        .ZN(n1961) );
  OAI22_X1 U1675 ( .A1(n1660), .A2(n1917), .B1(n1661), .B2(n1924), .ZN(n1962)
         );
  XNOR2_X1 U1676 ( .A(A[20]), .B(n1963), .ZN(n752) );
  AOI221_X1 U1677 ( .B1(n1921), .B2(B[22]), .C1(n1920), .C2(B[21]), .A(n1964), 
        .ZN(n1963) );
  OAI22_X1 U1678 ( .A1(n1562), .A2(n1917), .B1(n1564), .B2(n1924), .ZN(n1964)
         );
  XNOR2_X1 U1679 ( .A(A[20]), .B(n1965), .ZN(n751) );
  AOI221_X1 U1680 ( .B1(n1921), .B2(n1554), .C1(n1920), .C2(B[22]), .A(n1966), 
        .ZN(n1965) );
  OAI22_X1 U1681 ( .A1(n1567), .A2(n1917), .B1(n1568), .B2(n1924), .ZN(n1966)
         );
  XNOR2_X1 U1682 ( .A(A[20]), .B(n1967), .ZN(n750) );
  AOI221_X1 U1683 ( .B1(n1921), .B2(B[23]), .C1(n1920), .C2(n1554), .A(n1968), 
        .ZN(n1967) );
  OAI22_X1 U1684 ( .A1(n1571), .A2(n1917), .B1(n1572), .B2(n1924), .ZN(n1968)
         );
  XNOR2_X1 U1685 ( .A(A[20]), .B(n1969), .ZN(n749) );
  OAI221_X1 U1686 ( .B1(n1556), .B2(n1924), .C1(n1556), .C2(n1917), .A(n1970), 
        .ZN(n1969) );
  OAI21_X1 U1687 ( .B1(n1921), .B2(n1920), .A(n1554), .ZN(n1970) );
  INV_X1 U1688 ( .A(n1974), .ZN(n1971) );
  XNOR2_X1 U1689 ( .A(A[18]), .B(A[19]), .ZN(n1972) );
  XNOR2_X1 U1690 ( .A(A[19]), .B(n1543), .ZN(n1973) );
  XOR2_X1 U1691 ( .A(A[18]), .B(n1545), .Z(n1974) );
  XNOR2_X1 U1692 ( .A(n1975), .B(n1541), .ZN(n748) );
  OAI22_X1 U1693 ( .A1(n1574), .A2(n1535), .B1(n1574), .B2(n1976), .ZN(n1975)
         );
  XNOR2_X1 U1694 ( .A(n1977), .B(n1541), .ZN(n747) );
  OAI222_X1 U1695 ( .A1(n1578), .A2(n1535), .B1(n1574), .B2(n1534), .C1(n1580), 
        .C2(n1976), .ZN(n1977) );
  INV_X1 U1696 ( .A(n1397), .ZN(n1580) );
  XNOR2_X1 U1697 ( .A(n1540), .B(n1978), .ZN(n746) );
  AOI221_X1 U1698 ( .B1(n1537), .B2(B[2]), .C1(n1536), .C2(B[1]), .A(n1979), 
        .ZN(n1978) );
  OAI22_X1 U1699 ( .A1(n1585), .A2(n1976), .B1(n1574), .B2(n1538), .ZN(n1979)
         );
  INV_X1 U1700 ( .A(n1396), .ZN(n1585) );
  XNOR2_X1 U1701 ( .A(n1540), .B(n1981), .ZN(n745) );
  AOI221_X1 U1702 ( .B1(n1537), .B2(B[3]), .C1(n1536), .C2(B[2]), .A(n1982), 
        .ZN(n1981) );
  OAI22_X1 U1703 ( .A1(n1589), .A2(n1976), .B1(n1578), .B2(n1539), .ZN(n1982)
         );
  XNOR2_X1 U1704 ( .A(n1540), .B(n1983), .ZN(n744) );
  AOI221_X1 U1705 ( .B1(n1537), .B2(B[4]), .C1(n1536), .C2(B[3]), .A(n1984), 
        .ZN(n1983) );
  OAI22_X1 U1706 ( .A1(n1592), .A2(n1976), .B1(n1593), .B2(n1539), .ZN(n1984)
         );
  XNOR2_X1 U1707 ( .A(n1540), .B(n1985), .ZN(n743) );
  AOI221_X1 U1708 ( .B1(n1537), .B2(B[5]), .C1(n1536), .C2(B[4]), .A(n1986), 
        .ZN(n1985) );
  OAI22_X1 U1709 ( .A1(n1596), .A2(n1976), .B1(n1597), .B2(n1539), .ZN(n1986)
         );
  XNOR2_X1 U1710 ( .A(n1540), .B(n1987), .ZN(n742) );
  AOI221_X1 U1711 ( .B1(n1537), .B2(B[6]), .C1(n1536), .C2(B[5]), .A(n1988), 
        .ZN(n1987) );
  OAI22_X1 U1712 ( .A1(n1600), .A2(n1976), .B1(n1601), .B2(n1539), .ZN(n1988)
         );
  XNOR2_X1 U1713 ( .A(n1540), .B(n1989), .ZN(n741) );
  AOI221_X1 U1714 ( .B1(n1537), .B2(B[7]), .C1(n1536), .C2(B[6]), .A(n1990), 
        .ZN(n1989) );
  OAI22_X1 U1715 ( .A1(n1604), .A2(n1976), .B1(n1605), .B2(n1539), .ZN(n1990)
         );
  XNOR2_X1 U1716 ( .A(n1540), .B(n1991), .ZN(n740) );
  AOI221_X1 U1717 ( .B1(n1537), .B2(B[9]), .C1(n1536), .C2(B[8]), .A(n1992), 
        .ZN(n1991) );
  OAI22_X1 U1718 ( .A1(n1612), .A2(n1976), .B1(n1613), .B2(n1539), .ZN(n1992)
         );
  XNOR2_X1 U1719 ( .A(n1540), .B(n1993), .ZN(n739) );
  AOI221_X1 U1720 ( .B1(n1537), .B2(B[10]), .C1(n1536), .C2(B[9]), .A(n1994), 
        .ZN(n1993) );
  OAI22_X1 U1721 ( .A1(n1616), .A2(n1976), .B1(n1617), .B2(n1539), .ZN(n1994)
         );
  XNOR2_X1 U1722 ( .A(n1540), .B(n1995), .ZN(n738) );
  AOI221_X1 U1723 ( .B1(n1537), .B2(B[12]), .C1(n1536), .C2(B[11]), .A(n1996), 
        .ZN(n1995) );
  OAI22_X1 U1724 ( .A1(n1624), .A2(n1976), .B1(n1625), .B2(n1539), .ZN(n1996)
         );
  XNOR2_X1 U1725 ( .A(n1540), .B(n1997), .ZN(n737) );
  AOI221_X1 U1726 ( .B1(n1537), .B2(B[13]), .C1(n1536), .C2(B[12]), .A(n1998), 
        .ZN(n1997) );
  OAI22_X1 U1727 ( .A1(n1628), .A2(n1976), .B1(n1629), .B2(n1539), .ZN(n1998)
         );
  XNOR2_X1 U1728 ( .A(n1540), .B(n1999), .ZN(n736) );
  AOI221_X1 U1729 ( .B1(n1537), .B2(B[14]), .C1(n1536), .C2(B[13]), .A(n2000), 
        .ZN(n1999) );
  OAI22_X1 U1730 ( .A1(n1632), .A2(n1976), .B1(n1633), .B2(n1539), .ZN(n2000)
         );
  XNOR2_X1 U1731 ( .A(n1540), .B(n2001), .ZN(n735) );
  AOI221_X1 U1732 ( .B1(n1537), .B2(B[15]), .C1(n1536), .C2(B[14]), .A(n2002), 
        .ZN(n2001) );
  OAI22_X1 U1733 ( .A1(n1636), .A2(n1976), .B1(n1637), .B2(n1539), .ZN(n2002)
         );
  XNOR2_X1 U1734 ( .A(n1540), .B(n2003), .ZN(n734) );
  AOI221_X1 U1735 ( .B1(n1537), .B2(B[16]), .C1(n1536), .C2(B[15]), .A(n2004), 
        .ZN(n2003) );
  OAI22_X1 U1736 ( .A1(n1640), .A2(n1976), .B1(n1641), .B2(n1538), .ZN(n2004)
         );
  XNOR2_X1 U1737 ( .A(n1540), .B(n2005), .ZN(n733) );
  AOI221_X1 U1738 ( .B1(n1537), .B2(B[18]), .C1(n1536), .C2(B[17]), .A(n2006), 
        .ZN(n2005) );
  OAI22_X1 U1739 ( .A1(n1648), .A2(n1976), .B1(n1649), .B2(n1538), .ZN(n2006)
         );
  XNOR2_X1 U1740 ( .A(n1540), .B(n2007), .ZN(n732) );
  AOI221_X1 U1741 ( .B1(n1537), .B2(B[19]), .C1(n1536), .C2(B[18]), .A(n2008), 
        .ZN(n2007) );
  OAI22_X1 U1742 ( .A1(n1652), .A2(n1976), .B1(n1653), .B2(n1538), .ZN(n2008)
         );
  XNOR2_X1 U1743 ( .A(n1540), .B(n2009), .ZN(n731) );
  AOI221_X1 U1744 ( .B1(n1537), .B2(B[20]), .C1(n1536), .C2(B[19]), .A(n2010), 
        .ZN(n2009) );
  OAI22_X1 U1745 ( .A1(n1656), .A2(n1976), .B1(n1657), .B2(n1538), .ZN(n2010)
         );
  XNOR2_X1 U1746 ( .A(A[23]), .B(n2011), .ZN(n730) );
  AOI221_X1 U1747 ( .B1(n1537), .B2(B[21]), .C1(n1536), .C2(B[20]), .A(n2012), 
        .ZN(n2011) );
  OAI22_X1 U1748 ( .A1(n1660), .A2(n1976), .B1(n1661), .B2(n1538), .ZN(n2012)
         );
  XNOR2_X1 U1749 ( .A(A[23]), .B(n2013), .ZN(n729) );
  AOI221_X1 U1750 ( .B1(n1537), .B2(B[22]), .C1(n1536), .C2(B[21]), .A(n2014), 
        .ZN(n2013) );
  OAI22_X1 U1751 ( .A1(n1562), .A2(n1976), .B1(n1564), .B2(n1538), .ZN(n2014)
         );
  INV_X1 U1752 ( .A(B[20]), .ZN(n1564) );
  INV_X1 U1753 ( .A(n1376), .ZN(n1562) );
  XNOR2_X1 U1754 ( .A(n519), .B(n2015), .ZN(n506) );
  INV_X1 U1755 ( .A(n493), .ZN(n479) );
  NOR2_X1 U1756 ( .A1(n2015), .A2(n519), .ZN(n493) );
  XOR2_X1 U1757 ( .A(n2016), .B(n1674), .Z(n2015) );
  OAI221_X1 U1758 ( .B1(n1563), .B2(n1556), .C1(n1561), .C2(n1556), .A(n2017), 
        .ZN(n2016) );
  OAI21_X1 U1759 ( .B1(n1558), .B2(n1559), .A(n1554), .ZN(n2017) );
  INV_X1 U1760 ( .A(n454), .ZN(n442) );
  XOR2_X1 U1761 ( .A(n1540), .B(n2018), .Z(n454) );
  AOI221_X1 U1762 ( .B1(n1537), .B2(B[8]), .C1(n1536), .C2(B[7]), .A(n2019), 
        .ZN(n2018) );
  OAI22_X1 U1763 ( .A1(n1608), .A2(n1976), .B1(n1609), .B2(n1538), .ZN(n2019)
         );
  INV_X1 U1764 ( .A(n421), .ZN(n411) );
  XOR2_X1 U1765 ( .A(n1540), .B(n2020), .Z(n421) );
  AOI221_X1 U1766 ( .B1(n1537), .B2(B[11]), .C1(n1536), .C2(B[10]), .A(n2021), 
        .ZN(n2020) );
  OAI22_X1 U1767 ( .A1(n1620), .A2(n1976), .B1(n1621), .B2(n1538), .ZN(n2021)
         );
  INV_X1 U1768 ( .A(n387), .ZN(n395) );
  INV_X1 U1769 ( .A(n374), .ZN(n368) );
  XOR2_X1 U1770 ( .A(n1540), .B(n2022), .Z(n374) );
  AOI221_X1 U1771 ( .B1(n1537), .B2(B[17]), .C1(n1536), .C2(B[16]), .A(n2023), 
        .ZN(n2022) );
  OAI22_X1 U1772 ( .A1(n1644), .A2(n1976), .B1(n1645), .B2(n1538), .ZN(n2023)
         );
  INV_X1 U1773 ( .A(n356), .ZN(n360) );
  INV_X1 U1774 ( .A(n2024), .ZN(n351) );
  OAI222_X1 U1775 ( .A1(n2025), .A2(n2026), .B1(n2025), .B2(n2027), .C1(n2027), 
        .C2(n2026), .ZN(n326) );
  INV_X1 U1776 ( .A(n550), .ZN(n2027) );
  XNOR2_X1 U1777 ( .A(n1674), .B(n2028), .ZN(n2026) );
  AOI221_X1 U1778 ( .B1(B[21]), .B2(n1558), .C1(B[20]), .C2(n1559), .A(n2029), 
        .ZN(n2028) );
  OAI22_X1 U1779 ( .A1(n1561), .A2(n1660), .B1(n1563), .B2(n1661), .ZN(n2029)
         );
  INV_X1 U1780 ( .A(B[19]), .ZN(n1661) );
  INV_X1 U1781 ( .A(n1377), .ZN(n1660) );
  AOI222_X1 U1782 ( .A1(n2030), .A2(n2031), .B1(n2030), .B2(n564), .C1(n564), 
        .C2(n2031), .ZN(n2025) );
  XNOR2_X1 U1783 ( .A(A[2]), .B(n2032), .ZN(n2031) );
  AOI221_X1 U1784 ( .B1(B[20]), .B2(n1558), .C1(B[19]), .C2(n1559), .A(n2033), 
        .ZN(n2032) );
  OAI22_X1 U1785 ( .A1(n1561), .A2(n1656), .B1(n1563), .B2(n1657), .ZN(n2033)
         );
  INV_X1 U1786 ( .A(B[18]), .ZN(n1657) );
  INV_X1 U1787 ( .A(n1378), .ZN(n1656) );
  INV_X1 U1788 ( .A(n2034), .ZN(n2030) );
  AOI222_X1 U1789 ( .A1(n2035), .A2(n2036), .B1(n2035), .B2(n576), .C1(n576), 
        .C2(n2036), .ZN(n2034) );
  XNOR2_X1 U1790 ( .A(A[2]), .B(n2037), .ZN(n2036) );
  AOI221_X1 U1791 ( .B1(B[19]), .B2(n1558), .C1(B[18]), .C2(n1559), .A(n2038), 
        .ZN(n2037) );
  OAI22_X1 U1792 ( .A1(n1561), .A2(n1652), .B1(n1563), .B2(n1653), .ZN(n2038)
         );
  INV_X1 U1793 ( .A(B[17]), .ZN(n1653) );
  INV_X1 U1794 ( .A(n1379), .ZN(n1652) );
  OAI222_X1 U1795 ( .A1(n2039), .A2(n2040), .B1(n2039), .B2(n2041), .C1(n2041), 
        .C2(n2040), .ZN(n2035) );
  INV_X1 U1796 ( .A(n588), .ZN(n2041) );
  XNOR2_X1 U1797 ( .A(n1674), .B(n2042), .ZN(n2040) );
  AOI221_X1 U1798 ( .B1(B[18]), .B2(n1558), .C1(B[17]), .C2(n1559), .A(n2043), 
        .ZN(n2042) );
  OAI22_X1 U1799 ( .A1(n1561), .A2(n1648), .B1(n1563), .B2(n1649), .ZN(n2043)
         );
  INV_X1 U1800 ( .A(B[16]), .ZN(n1649) );
  INV_X1 U1801 ( .A(n1380), .ZN(n1648) );
  AOI222_X1 U1802 ( .A1(n2044), .A2(n2045), .B1(n2044), .B2(n600), .C1(n600), 
        .C2(n2045), .ZN(n2039) );
  XNOR2_X1 U1803 ( .A(A[2]), .B(n2046), .ZN(n2045) );
  AOI221_X1 U1804 ( .B1(B[17]), .B2(n1558), .C1(B[16]), .C2(n1559), .A(n2047), 
        .ZN(n2046) );
  OAI22_X1 U1805 ( .A1(n1561), .A2(n1644), .B1(n1563), .B2(n1645), .ZN(n2047)
         );
  INV_X1 U1806 ( .A(B[15]), .ZN(n1645) );
  INV_X1 U1807 ( .A(n1381), .ZN(n1644) );
  OAI222_X1 U1808 ( .A1(n2048), .A2(n2049), .B1(n2048), .B2(n2050), .C1(n2050), 
        .C2(n2049), .ZN(n2044) );
  INV_X1 U1809 ( .A(n610), .ZN(n2050) );
  XNOR2_X1 U1810 ( .A(n1674), .B(n2051), .ZN(n2049) );
  AOI221_X1 U1811 ( .B1(B[16]), .B2(n1558), .C1(B[15]), .C2(n1559), .A(n2052), 
        .ZN(n2051) );
  OAI22_X1 U1812 ( .A1(n1561), .A2(n1640), .B1(n1563), .B2(n1641), .ZN(n2052)
         );
  INV_X1 U1813 ( .A(B[14]), .ZN(n1641) );
  INV_X1 U1814 ( .A(n1382), .ZN(n1640) );
  AOI222_X1 U1815 ( .A1(n2053), .A2(n2054), .B1(n2053), .B2(n620), .C1(n620), 
        .C2(n2054), .ZN(n2048) );
  XNOR2_X1 U1816 ( .A(A[2]), .B(n2055), .ZN(n2054) );
  AOI221_X1 U1817 ( .B1(B[15]), .B2(n1558), .C1(B[14]), .C2(n1559), .A(n2056), 
        .ZN(n2055) );
  OAI22_X1 U1818 ( .A1(n1561), .A2(n1636), .B1(n1563), .B2(n1637), .ZN(n2056)
         );
  INV_X1 U1819 ( .A(B[13]), .ZN(n1637) );
  INV_X1 U1820 ( .A(n1383), .ZN(n1636) );
  OAI222_X1 U1821 ( .A1(n2057), .A2(n2058), .B1(n2057), .B2(n2059), .C1(n2059), 
        .C2(n2058), .ZN(n2053) );
  INV_X1 U1822 ( .A(n630), .ZN(n2059) );
  XNOR2_X1 U1823 ( .A(n1674), .B(n2060), .ZN(n2058) );
  AOI221_X1 U1824 ( .B1(B[14]), .B2(n1558), .C1(B[13]), .C2(n1559), .A(n2061), 
        .ZN(n2060) );
  OAI22_X1 U1825 ( .A1(n1561), .A2(n1632), .B1(n1563), .B2(n1633), .ZN(n2061)
         );
  INV_X1 U1826 ( .A(B[12]), .ZN(n1633) );
  INV_X1 U1827 ( .A(n1384), .ZN(n1632) );
  AOI222_X1 U1828 ( .A1(n2062), .A2(n2063), .B1(n2062), .B2(n638), .C1(n638), 
        .C2(n2063), .ZN(n2057) );
  XNOR2_X1 U1829 ( .A(A[2]), .B(n2064), .ZN(n2063) );
  AOI221_X1 U1830 ( .B1(B[13]), .B2(n1558), .C1(B[12]), .C2(n1559), .A(n2065), 
        .ZN(n2064) );
  OAI22_X1 U1831 ( .A1(n1561), .A2(n1628), .B1(n1563), .B2(n1629), .ZN(n2065)
         );
  INV_X1 U1832 ( .A(B[11]), .ZN(n1629) );
  INV_X1 U1833 ( .A(n1385), .ZN(n1628) );
  OAI222_X1 U1834 ( .A1(n2066), .A2(n2067), .B1(n2066), .B2(n2068), .C1(n2068), 
        .C2(n2067), .ZN(n2062) );
  INV_X1 U1835 ( .A(n646), .ZN(n2068) );
  XNOR2_X1 U1836 ( .A(n1674), .B(n2069), .ZN(n2067) );
  AOI221_X1 U1837 ( .B1(B[12]), .B2(n1558), .C1(B[11]), .C2(n1559), .A(n2070), 
        .ZN(n2069) );
  OAI22_X1 U1838 ( .A1(n1561), .A2(n1624), .B1(n1563), .B2(n1625), .ZN(n2070)
         );
  INV_X1 U1839 ( .A(B[10]), .ZN(n1625) );
  INV_X1 U1840 ( .A(n1386), .ZN(n1624) );
  AOI222_X1 U1841 ( .A1(n2071), .A2(n2072), .B1(n2071), .B2(n654), .C1(n654), 
        .C2(n2072), .ZN(n2066) );
  XNOR2_X1 U1842 ( .A(A[2]), .B(n2073), .ZN(n2072) );
  AOI221_X1 U1843 ( .B1(B[11]), .B2(n1558), .C1(B[10]), .C2(n1559), .A(n2074), 
        .ZN(n2073) );
  OAI22_X1 U1844 ( .A1(n1561), .A2(n1620), .B1(n1563), .B2(n1621), .ZN(n2074)
         );
  INV_X1 U1845 ( .A(B[9]), .ZN(n1621) );
  INV_X1 U1846 ( .A(n1387), .ZN(n1620) );
  OAI222_X1 U1847 ( .A1(n2075), .A2(n2076), .B1(n2075), .B2(n2077), .C1(n2077), 
        .C2(n2076), .ZN(n2071) );
  INV_X1 U1848 ( .A(n660), .ZN(n2077) );
  XNOR2_X1 U1849 ( .A(n1674), .B(n2078), .ZN(n2076) );
  AOI221_X1 U1850 ( .B1(B[10]), .B2(n1558), .C1(B[9]), .C2(n1559), .A(n2079), 
        .ZN(n2078) );
  OAI22_X1 U1851 ( .A1(n1561), .A2(n1616), .B1(n1563), .B2(n1617), .ZN(n2079)
         );
  INV_X1 U1852 ( .A(B[8]), .ZN(n1617) );
  INV_X1 U1853 ( .A(n1388), .ZN(n1616) );
  AOI222_X1 U1854 ( .A1(n2080), .A2(n2081), .B1(n2080), .B2(n666), .C1(n666), 
        .C2(n2081), .ZN(n2075) );
  XNOR2_X1 U1855 ( .A(A[2]), .B(n2082), .ZN(n2081) );
  AOI221_X1 U1856 ( .B1(B[9]), .B2(n1558), .C1(B[8]), .C2(n1559), .A(n2083), 
        .ZN(n2082) );
  OAI22_X1 U1857 ( .A1(n1561), .A2(n1612), .B1(n1563), .B2(n1613), .ZN(n2083)
         );
  INV_X1 U1858 ( .A(B[7]), .ZN(n1613) );
  INV_X1 U1859 ( .A(n1389), .ZN(n1612) );
  OAI222_X1 U1860 ( .A1(n2084), .A2(n2085), .B1(n2084), .B2(n2086), .C1(n2086), 
        .C2(n2085), .ZN(n2080) );
  INV_X1 U1861 ( .A(n672), .ZN(n2086) );
  XNOR2_X1 U1862 ( .A(n1674), .B(n2087), .ZN(n2085) );
  AOI221_X1 U1863 ( .B1(B[8]), .B2(n1558), .C1(B[7]), .C2(n1559), .A(n2088), 
        .ZN(n2087) );
  OAI22_X1 U1864 ( .A1(n1561), .A2(n1608), .B1(n1563), .B2(n1609), .ZN(n2088)
         );
  INV_X1 U1865 ( .A(B[6]), .ZN(n1609) );
  INV_X1 U1866 ( .A(n1390), .ZN(n1608) );
  AOI222_X1 U1867 ( .A1(n2089), .A2(n2090), .B1(n2089), .B2(n676), .C1(n676), 
        .C2(n2090), .ZN(n2084) );
  XNOR2_X1 U1868 ( .A(A[2]), .B(n2091), .ZN(n2090) );
  AOI221_X1 U1869 ( .B1(B[7]), .B2(n1558), .C1(B[6]), .C2(n1559), .A(n2092), 
        .ZN(n2091) );
  OAI22_X1 U1870 ( .A1(n1561), .A2(n1604), .B1(n1563), .B2(n1605), .ZN(n2092)
         );
  INV_X1 U1871 ( .A(B[5]), .ZN(n1605) );
  INV_X1 U1872 ( .A(n1391), .ZN(n1604) );
  OAI222_X1 U1873 ( .A1(n2093), .A2(n2094), .B1(n2093), .B2(n2095), .C1(n2095), 
        .C2(n2094), .ZN(n2089) );
  INV_X1 U1874 ( .A(n680), .ZN(n2095) );
  XNOR2_X1 U1875 ( .A(n1674), .B(n2096), .ZN(n2094) );
  AOI221_X1 U1876 ( .B1(B[6]), .B2(n1558), .C1(B[5]), .C2(n1559), .A(n2097), 
        .ZN(n2096) );
  OAI22_X1 U1877 ( .A1(n1561), .A2(n1600), .B1(n1563), .B2(n1601), .ZN(n2097)
         );
  INV_X1 U1878 ( .A(B[4]), .ZN(n1601) );
  INV_X1 U1879 ( .A(n1392), .ZN(n1600) );
  AOI222_X1 U1880 ( .A1(n2098), .A2(n2099), .B1(n2098), .B2(n684), .C1(n684), 
        .C2(n2099), .ZN(n2093) );
  XNOR2_X1 U1881 ( .A(A[2]), .B(n2100), .ZN(n2099) );
  AOI221_X1 U1882 ( .B1(B[5]), .B2(n1558), .C1(B[4]), .C2(n1559), .A(n2101), 
        .ZN(n2100) );
  OAI22_X1 U1883 ( .A1(n1561), .A2(n1596), .B1(n1563), .B2(n1597), .ZN(n2101)
         );
  INV_X1 U1884 ( .A(B[3]), .ZN(n1597) );
  INV_X1 U1885 ( .A(n1393), .ZN(n1596) );
  OAI222_X1 U1886 ( .A1(n2102), .A2(n2103), .B1(n2102), .B2(n2104), .C1(n2104), 
        .C2(n2103), .ZN(n2098) );
  INV_X1 U1887 ( .A(n686), .ZN(n2104) );
  XNOR2_X1 U1888 ( .A(n1674), .B(n2105), .ZN(n2103) );
  AOI221_X1 U1889 ( .B1(B[4]), .B2(n1558), .C1(B[3]), .C2(n1559), .A(n2106), 
        .ZN(n2105) );
  OAI22_X1 U1890 ( .A1(n1561), .A2(n1592), .B1(n1563), .B2(n1593), .ZN(n2106)
         );
  INV_X1 U1891 ( .A(B[2]), .ZN(n1593) );
  INV_X1 U1892 ( .A(n1394), .ZN(n1592) );
  AOI222_X1 U1893 ( .A1(n2107), .A2(n2108), .B1(n2107), .B2(n688), .C1(n688), 
        .C2(n2108), .ZN(n2102) );
  XNOR2_X1 U1894 ( .A(A[2]), .B(n2109), .ZN(n2108) );
  AOI221_X1 U1895 ( .B1(B[3]), .B2(n1558), .C1(B[2]), .C2(n1559), .A(n2110), 
        .ZN(n2109) );
  OAI22_X1 U1896 ( .A1(n1561), .A2(n1589), .B1(n1563), .B2(n1578), .ZN(n2110)
         );
  INV_X1 U1897 ( .A(B[1]), .ZN(n1578) );
  INV_X1 U1898 ( .A(n1395), .ZN(n1589) );
  AND2_X1 U1899 ( .A1(n2114), .A2(n2115), .ZN(n2107) );
  AOI211_X1 U1900 ( .C1(B[1]), .C2(n1558), .A(n2116), .B(B[0]), .ZN(n2115) );
  INV_X1 U1901 ( .A(n2117), .ZN(n2116) );
  AOI22_X1 U1902 ( .A1(n1558), .A2(B[2]), .B1(n2118), .B2(n1397), .ZN(n2117)
         );
  INV_X1 U1903 ( .A(A[0]), .ZN(n2112) );
  AOI221_X1 U1904 ( .B1(B[1]), .B2(n1559), .C1(n1396), .C2(n2118), .A(n1674), 
        .ZN(n2114) );
  INV_X1 U1905 ( .A(n1561), .ZN(n2118) );
  XNOR2_X1 U1906 ( .A(A[1]), .B(n1674), .ZN(n2111) );
  INV_X1 U1907 ( .A(A[2]), .ZN(n1674) );
  INV_X1 U1908 ( .A(A[1]), .ZN(n2113) );
  AOI21_X1 U1909 ( .B1(n2119), .B2(n2120), .A(n2121), .ZN(PRODUCT[47]) );
  OAI22_X1 U1910 ( .A1(n2122), .A2(n2123), .B1(n2122), .B2(n2124), .ZN(n2121)
         );
  INV_X1 U1911 ( .A(n2120), .ZN(n2124) );
  AOI222_X1 U1912 ( .A1(n2024), .A2(n303), .B1(n2123), .B2(n303), .C1(n2024), 
        .C2(n2123), .ZN(n2122) );
  XOR2_X1 U1913 ( .A(n1541), .B(n2125), .Z(n2024) );
  AOI221_X1 U1914 ( .B1(n1537), .B2(B[23]), .C1(n1536), .C2(B[22]), .A(n2126), 
        .ZN(n2125) );
  OAI22_X1 U1915 ( .A1(n1567), .A2(n1976), .B1(n1568), .B2(n1538), .ZN(n2126)
         );
  INV_X1 U1916 ( .A(B[21]), .ZN(n1568) );
  INV_X1 U1917 ( .A(n1375), .ZN(n1567) );
  XOR2_X1 U1918 ( .A(n2127), .B(n1541), .Z(n2120) );
  OAI221_X1 U1919 ( .B1(n1556), .B2(n1539), .C1(n1556), .C2(n1976), .A(n2128), 
        .ZN(n2127) );
  OAI21_X1 U1920 ( .B1(n1537), .B2(n1536), .A(n1554), .ZN(n2128) );
  INV_X1 U1921 ( .A(n2123), .ZN(n2119) );
  XOR2_X1 U1922 ( .A(A[23]), .B(n2129), .Z(n2123) );
  AOI221_X1 U1923 ( .B1(n1537), .B2(n1554), .C1(n1536), .C2(n1554), .A(n2130), 
        .ZN(n2129) );
  OAI22_X1 U1924 ( .A1(n1571), .A2(n1976), .B1(n1572), .B2(n1538), .ZN(n2130)
         );
  NAND3_X1 U1925 ( .A1(n2131), .A2(n2132), .A3(n2133), .ZN(n1980) );
  INV_X1 U1926 ( .A(B[22]), .ZN(n1572) );
  INV_X1 U1927 ( .A(n1374), .ZN(n1571) );
  XNOR2_X1 U1928 ( .A(A[21]), .B(A[22]), .ZN(n2133) );
  INV_X1 U1929 ( .A(n2131), .ZN(n2134) );
  XOR2_X1 U1930 ( .A(A[21]), .B(n1543), .Z(n2131) );
  XNOR2_X1 U1931 ( .A(A[22]), .B(n1541), .ZN(n2132) );
endmodule


module iir_filter_DW01_add_3 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   carry_23_, carry_22_, carry_21_, carry_20_, carry_19_, carry_18_,
         carry_17_, carry_16_, carry_15_, carry_14_, carry_13_, carry_12_,
         carry_11_, carry_10_, carry_9_, carry_8_, carry_7_, carry_6_,
         carry_5_, carry_4_, carry_3_, carry_2_, carry_1_;

  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry_23_), .S(SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry_22_), .CO(carry_23_), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry_21_), .CO(carry_22_), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry_20_), .CO(carry_21_), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry_19_), .CO(carry_20_), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry_18_), .CO(carry_19_), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry_17_), .CO(carry_18_), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry_16_), .CO(carry_17_), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry_15_), .CO(carry_16_), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry_14_), .CO(carry_15_), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry_13_), .CO(carry_14_), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry_12_), .CO(carry_13_), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry_11_), .CO(carry_12_), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry_10_), .CO(carry_11_), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry_9_), .CO(carry_10_), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry_8_), .CO(carry_9_), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry_7_), .CO(carry_8_), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry_6_), .CO(carry_7_), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry_5_), .CO(carry_6_), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry_4_), .CO(carry_5_), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry_3_), .CO(carry_4_), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry_2_), .CO(carry_3_), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry_1_), .CO(carry_2_), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(A[0]), .A2(B[0]), .ZN(carry_1_) );
  XOR2_X1 U2 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module iir_filter_DW01_add_2 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   carry_23_, carry_22_, carry_21_, carry_20_, carry_19_, carry_18_,
         carry_17_, carry_16_, carry_15_, carry_14_, carry_13_, carry_12_,
         carry_11_, carry_10_, carry_9_, carry_8_, carry_7_, carry_6_,
         carry_5_, carry_4_, carry_3_, carry_2_, carry_1_;

  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry_23_), .S(SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry_22_), .CO(carry_23_), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry_21_), .CO(carry_22_), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry_20_), .CO(carry_21_), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry_19_), .CO(carry_20_), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry_18_), .CO(carry_19_), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry_17_), .CO(carry_18_), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry_16_), .CO(carry_17_), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry_15_), .CO(carry_16_), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry_14_), .CO(carry_15_), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry_13_), .CO(carry_14_), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry_12_), .CO(carry_13_), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry_11_), .CO(carry_12_), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry_10_), .CO(carry_11_), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry_9_), .CO(carry_10_), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry_8_), .CO(carry_9_), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry_7_), .CO(carry_8_), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry_6_), .CO(carry_7_), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry_5_), .CO(carry_6_), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry_4_), .CO(carry_5_), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry_3_), .CO(carry_4_), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry_2_), .CO(carry_3_), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry_1_), .CO(carry_2_), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(A[0]), .A2(B[0]), .ZN(carry_1_) );
  XOR2_X1 U2 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module iir_filter_DW01_add_1 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   carry_23_, carry_22_, carry_21_, carry_20_, carry_19_, carry_18_,
         carry_17_, carry_16_, carry_15_, carry_14_, carry_13_, carry_12_,
         carry_11_, carry_10_, carry_9_, carry_8_, carry_7_, carry_6_,
         carry_5_, carry_4_, carry_3_, carry_2_, carry_1_;

  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry_23_), .S(SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry_22_), .CO(carry_23_), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry_21_), .CO(carry_22_), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry_20_), .CO(carry_21_), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry_19_), .CO(carry_20_), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry_18_), .CO(carry_19_), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry_17_), .CO(carry_18_), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry_16_), .CO(carry_17_), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry_15_), .CO(carry_16_), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry_14_), .CO(carry_15_), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry_13_), .CO(carry_14_), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry_12_), .CO(carry_13_), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry_11_), .CO(carry_12_), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry_10_), .CO(carry_11_), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry_9_), .CO(carry_10_), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry_8_), .CO(carry_9_), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry_7_), .CO(carry_8_), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry_6_), .CO(carry_7_), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry_5_), .CO(carry_6_), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry_4_), .CO(carry_5_), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry_3_), .CO(carry_4_), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry_2_), .CO(carry_3_), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry_1_), .CO(carry_2_), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(A[0]), .A2(B[0]), .ZN(carry_1_) );
  XOR2_X1 U2 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module iir_filter_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] DIFF;
  input CI;
  output CO;
  wire   B_0_, carry_23_, carry_22_, carry_21_, carry_20_, carry_19_,
         carry_18_, carry_17_, carry_16_, carry_15_, carry_14_, carry_13_,
         carry_12_, carry_11_, carry_10_, carry_9_, carry_8_, carry_7_,
         carry_6_, carry_5_, carry_4_, carry_3_, carry_2_, carry_1_, B_not_23_,
         B_not_22_, B_not_21_, B_not_20_, B_not_19_, B_not_18_, B_not_17_,
         B_not_16_, B_not_15_, B_not_14_, B_not_13_, B_not_12_, B_not_11_,
         B_not_10_, B_not_9_, B_not_8_, B_not_7_, B_not_6_, B_not_5_, B_not_4_,
         B_not_3_, B_not_2_, B_not_1_;
  assign DIFF[0] = B_0_;
  assign B_0_ = B[0];

  FA_X1 U2_23 ( .A(A[23]), .B(B_not_23_), .CI(carry_23_), .S(DIFF[23]) );
  FA_X1 U2_22 ( .A(A[22]), .B(B_not_22_), .CI(carry_22_), .CO(carry_23_), .S(
        DIFF[22]) );
  FA_X1 U2_21 ( .A(A[21]), .B(B_not_21_), .CI(carry_21_), .CO(carry_22_), .S(
        DIFF[21]) );
  FA_X1 U2_20 ( .A(A[20]), .B(B_not_20_), .CI(carry_20_), .CO(carry_21_), .S(
        DIFF[20]) );
  FA_X1 U2_19 ( .A(A[19]), .B(B_not_19_), .CI(carry_19_), .CO(carry_20_), .S(
        DIFF[19]) );
  FA_X1 U2_18 ( .A(A[18]), .B(B_not_18_), .CI(carry_18_), .CO(carry_19_), .S(
        DIFF[18]) );
  FA_X1 U2_17 ( .A(A[17]), .B(B_not_17_), .CI(carry_17_), .CO(carry_18_), .S(
        DIFF[17]) );
  FA_X1 U2_16 ( .A(A[16]), .B(B_not_16_), .CI(carry_16_), .CO(carry_17_), .S(
        DIFF[16]) );
  FA_X1 U2_15 ( .A(A[15]), .B(B_not_15_), .CI(carry_15_), .CO(carry_16_), .S(
        DIFF[15]) );
  FA_X1 U2_14 ( .A(A[14]), .B(B_not_14_), .CI(carry_14_), .CO(carry_15_), .S(
        DIFF[14]) );
  FA_X1 U2_13 ( .A(A[13]), .B(B_not_13_), .CI(carry_13_), .CO(carry_14_), .S(
        DIFF[13]) );
  FA_X1 U2_12 ( .A(A[12]), .B(B_not_12_), .CI(carry_12_), .CO(carry_13_), .S(
        DIFF[12]) );
  FA_X1 U2_11 ( .A(A[11]), .B(B_not_11_), .CI(carry_11_), .CO(carry_12_), .S(
        DIFF[11]) );
  AND2_X1 U1 ( .A1(carry_10_), .A2(B_not_10_), .ZN(carry_11_) );
  XOR2_X1 U2 ( .A(B_not_10_), .B(carry_10_), .Z(DIFF[10]) );
  AND2_X1 U3 ( .A1(carry_9_), .A2(B_not_9_), .ZN(carry_10_) );
  XOR2_X1 U4 ( .A(B_not_9_), .B(carry_9_), .Z(DIFF[9]) );
  AND2_X1 U5 ( .A1(carry_8_), .A2(B_not_8_), .ZN(carry_9_) );
  XOR2_X1 U6 ( .A(B_not_8_), .B(carry_8_), .Z(DIFF[8]) );
  AND2_X1 U7 ( .A1(carry_7_), .A2(B_not_7_), .ZN(carry_8_) );
  XOR2_X1 U8 ( .A(B_not_7_), .B(carry_7_), .Z(DIFF[7]) );
  AND2_X1 U9 ( .A1(carry_6_), .A2(B_not_6_), .ZN(carry_7_) );
  XOR2_X1 U10 ( .A(B_not_6_), .B(carry_6_), .Z(DIFF[6]) );
  AND2_X1 U11 ( .A1(carry_5_), .A2(B_not_5_), .ZN(carry_6_) );
  XOR2_X1 U12 ( .A(B_not_5_), .B(carry_5_), .Z(DIFF[5]) );
  AND2_X1 U13 ( .A1(carry_4_), .A2(B_not_4_), .ZN(carry_5_) );
  XOR2_X1 U14 ( .A(B_not_4_), .B(carry_4_), .Z(DIFF[4]) );
  AND2_X1 U15 ( .A1(carry_3_), .A2(B_not_3_), .ZN(carry_4_) );
  XOR2_X1 U16 ( .A(B_not_3_), .B(carry_3_), .Z(DIFF[3]) );
  AND2_X1 U17 ( .A1(carry_2_), .A2(B_not_2_), .ZN(carry_3_) );
  XOR2_X1 U18 ( .A(B_not_2_), .B(carry_2_), .Z(DIFF[2]) );
  AND2_X1 U19 ( .A1(carry_1_), .A2(B_not_1_), .ZN(carry_2_) );
  XOR2_X1 U20 ( .A(B_not_1_), .B(carry_1_), .Z(DIFF[1]) );
  INV_X1 U21 ( .A(B_0_), .ZN(carry_1_) );
  INV_X1 U22 ( .A(B[9]), .ZN(B_not_9_) );
  INV_X1 U23 ( .A(B[8]), .ZN(B_not_8_) );
  INV_X1 U24 ( .A(B[7]), .ZN(B_not_7_) );
  INV_X1 U25 ( .A(B[6]), .ZN(B_not_6_) );
  INV_X1 U26 ( .A(B[5]), .ZN(B_not_5_) );
  INV_X1 U27 ( .A(B[4]), .ZN(B_not_4_) );
  INV_X1 U28 ( .A(B[3]), .ZN(B_not_3_) );
  INV_X1 U29 ( .A(B[2]), .ZN(B_not_2_) );
  INV_X1 U30 ( .A(B[23]), .ZN(B_not_23_) );
  INV_X1 U31 ( .A(B[22]), .ZN(B_not_22_) );
  INV_X1 U32 ( .A(B[21]), .ZN(B_not_21_) );
  INV_X1 U33 ( .A(B[20]), .ZN(B_not_20_) );
  INV_X1 U34 ( .A(B[1]), .ZN(B_not_1_) );
  INV_X1 U35 ( .A(B[19]), .ZN(B_not_19_) );
  INV_X1 U36 ( .A(B[18]), .ZN(B_not_18_) );
  INV_X1 U37 ( .A(B[17]), .ZN(B_not_17_) );
  INV_X1 U38 ( .A(B[16]), .ZN(B_not_16_) );
  INV_X1 U39 ( .A(B[15]), .ZN(B_not_15_) );
  INV_X1 U40 ( .A(B[14]), .ZN(B_not_14_) );
  INV_X1 U41 ( .A(B[13]), .ZN(B_not_13_) );
  INV_X1 U42 ( .A(B[12]), .ZN(B_not_12_) );
  INV_X1 U43 ( .A(B[11]), .ZN(B_not_11_) );
  INV_X1 U44 ( .A(B[10]), .ZN(B_not_10_) );
endmodule


module iir_filter_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   carry_23_, carry_22_, carry_21_, carry_20_, carry_19_, carry_18_,
         carry_17_, carry_16_, carry_15_, carry_14_, carry_13_, carry_12_,
         carry_11_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37;

  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry_23_), .S(SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry_22_), .CO(carry_23_), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry_21_), .CO(carry_22_), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry_20_), .CO(carry_21_), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry_19_), .CO(carry_20_), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry_18_), .CO(carry_19_), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry_17_), .CO(carry_18_), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry_16_), .CO(carry_17_), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry_15_), .CO(carry_16_), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry_14_), .CO(carry_15_), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry_13_), .CO(carry_14_), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry_12_), .CO(carry_13_), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry_11_), .CO(carry_12_), .S(
        SUM[11]) );
  OAI21_X1 U1 ( .B1(n1), .B2(n2), .A(n3), .ZN(carry_11_) );
  OAI21_X1 U2 ( .B1(A[10]), .B2(n4), .A(B[10]), .ZN(n3) );
  INV_X1 U3 ( .A(n1), .ZN(n4) );
  INV_X1 U4 ( .A(A[10]), .ZN(n2) );
  AOI21_X1 U5 ( .B1(n5), .B2(A[9]), .A(n6), .ZN(n1) );
  INV_X1 U6 ( .A(n7), .ZN(n6) );
  OAI21_X1 U7 ( .B1(A[9]), .B2(n5), .A(B[9]), .ZN(n7) );
  OAI21_X1 U8 ( .B1(n8), .B2(n9), .A(n10), .ZN(n5) );
  OAI21_X1 U9 ( .B1(A[8]), .B2(n11), .A(B[8]), .ZN(n10) );
  INV_X1 U10 ( .A(n8), .ZN(n11) );
  INV_X1 U11 ( .A(A[8]), .ZN(n9) );
  AOI21_X1 U12 ( .B1(n12), .B2(A[7]), .A(n13), .ZN(n8) );
  INV_X1 U13 ( .A(n14), .ZN(n13) );
  OAI21_X1 U14 ( .B1(A[7]), .B2(n12), .A(B[7]), .ZN(n14) );
  OAI21_X1 U15 ( .B1(n15), .B2(n16), .A(n17), .ZN(n12) );
  OAI21_X1 U16 ( .B1(A[6]), .B2(n18), .A(B[6]), .ZN(n17) );
  INV_X1 U17 ( .A(A[6]), .ZN(n16) );
  INV_X1 U18 ( .A(n18), .ZN(n15) );
  OAI21_X1 U19 ( .B1(n19), .B2(n20), .A(n21), .ZN(n18) );
  OAI21_X1 U20 ( .B1(A[5]), .B2(n22), .A(B[5]), .ZN(n21) );
  INV_X1 U21 ( .A(A[5]), .ZN(n20) );
  INV_X1 U22 ( .A(n22), .ZN(n19) );
  OAI21_X1 U23 ( .B1(n23), .B2(n24), .A(n25), .ZN(n22) );
  OAI21_X1 U24 ( .B1(A[4]), .B2(n26), .A(B[4]), .ZN(n25) );
  INV_X1 U25 ( .A(A[4]), .ZN(n24) );
  INV_X1 U26 ( .A(n26), .ZN(n23) );
  OAI21_X1 U27 ( .B1(n27), .B2(n28), .A(n29), .ZN(n26) );
  OAI21_X1 U28 ( .B1(A[3]), .B2(n30), .A(B[3]), .ZN(n29) );
  INV_X1 U29 ( .A(A[3]), .ZN(n28) );
  INV_X1 U30 ( .A(n30), .ZN(n27) );
  OAI21_X1 U31 ( .B1(n31), .B2(n32), .A(n33), .ZN(n30) );
  OAI21_X1 U32 ( .B1(A[2]), .B2(n34), .A(B[2]), .ZN(n33) );
  INV_X1 U33 ( .A(A[2]), .ZN(n32) );
  INV_X1 U34 ( .A(n34), .ZN(n31) );
  OAI21_X1 U35 ( .B1(n35), .B2(n36), .A(n37), .ZN(n34) );
  OAI211_X1 U36 ( .C1(A[1]), .C2(B[1]), .A(A[0]), .B(B[0]), .ZN(n37) );
  INV_X1 U37 ( .A(B[1]), .ZN(n36) );
  INV_X1 U38 ( .A(A[1]), .ZN(n35) );
endmodule


module iir_filter ( clk, rst_n, vIn, dIn, coeffs_fb, coeffs_ff, dOut, vOut );
  input [11:0] dIn;
  input [47:0] coeffs_fb;
  input [95:0] coeffs_ff;
  output [11:0] dOut;
  input clk, rst_n, vIn;
  output vOut;
  wire   delayed_controls_0__1_, delayed_controls_1__0_,
         delayed_controls_1__1_, delayed_controls_2__0_, DP_N4, DP_N2, DP_y_0_,
         DP_y_1_, DP_y_2_, DP_y_3_, DP_y_4_, DP_y_5_, DP_y_6_, DP_y_7_,
         DP_y_8_, DP_y_9_, DP_y_10_, DP_y_11_, DP_y_23, DP_sw1_0_, DP_sw1_1_,
         DP_sw1_2_, DP_sw1_3_, DP_sw1_4_, DP_sw1_5_, DP_sw1_6_, DP_sw1_7_,
         DP_sw1_8_, DP_sw1_9_, DP_sw1_10_, DP_sw1_11_, DP_sw1_12_, DP_sw1_13_,
         DP_sw1_14_, DP_sw1_15_, DP_sw1_16_, DP_sw1_17_, DP_sw1_18_,
         DP_sw1_19_, DP_sw1_20_, DP_sw1_21_, DP_sw1_22_, DP_sw1_23_, DP_sw0_0_,
         DP_sw0_1_, DP_sw0_2_, DP_sw0_3_, DP_sw0_4_, DP_sw0_5_, DP_sw0_6_,
         DP_sw0_7_, DP_sw0_8_, DP_sw0_9_, DP_sw0_10_, DP_sw0_11_, DP_sw0_12_,
         DP_sw0_13_, DP_sw0_14_, DP_sw0_15_, DP_sw0_16_, DP_sw0_17_,
         DP_sw0_18_, DP_sw0_19_, DP_sw0_20_, DP_sw0_21_, DP_sw0_22_,
         DP_sw0_23_, DP_w_0_, DP_w_1_, DP_w_2_, DP_w_3_, DP_w_4_, DP_w_5_,
         DP_w_6_, DP_w_7_, DP_w_8_, DP_w_9_, DP_w_10_, DP_w_11_, DP_w_12_,
         DP_w_13_, DP_w_14_, DP_w_15_, DP_w_16_, DP_w_17_, DP_w_18_, DP_w_19_,
         DP_w_20_, DP_w_21_, DP_w_22_, DP_w_23_, CU_nextState_0_, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n72, n73, n74, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n560, n562, n564, n566, n568,
         n570, n572, n574, n576, n578, n580, n582, n584, n586, n588, n590,
         n592, n594, n596, n598, n600, n602, n604, n606, n706, n707, n711,
         n712, n716, n717, n721, n722, n726, n727, n731, n732, n736, n737,
         n741, n742, n746, n747, n751, n752, n756, n757, n761, n762, n766,
         n767, n771, n772, n776, n777, n781, n782, n786, n787, n791, n792,
         n796, n797, n801, n802, n806, n807, n811, n812, n816, n817, n820,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141;
  wire   [0:23] DP_ff;
  wire   [0:23] DP_ff_part;
  wire   [0:23] DP_fb;
  wire   [0:23] DP_pipe13;
  wire   [0:23] DP_pipe0_coeff_pipe03;
  wire   [0:23] DP_pipe12;
  wire   [0:23] DP_pipe0_coeff_pipe02;
  wire   [0:23] DP_pipe11;
  wire   [0:23] DP_pipe0_coeff_pipe01;
  wire   [0:23] DP_pipe10;
  wire   [0:23] DP_pipe0_coeff_pipe00;
  wire   [0:23] DP_pipe03;
  wire   [0:23] DP_pipe02;
  wire   [0:23] DP_pipe01;
  wire   [0:23] DP_pipe00;
  wire   [0:23] DP_ret1;
  wire   [0:23] DP_sw1_coeff_ret1;
  wire   [0:23] DP_ret0;
  wire   [0:23] DP_sw0_coeff_ret0;
  wire   [0:23] DP_sw2;
  wire   [95:0] DP_coeffs_ff_int;
  wire   [47:0] DP_coeffs_fb_int;
  wire   [0:11] DP_x;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154;

  DFFR_X1 DP_reg_in_Q_reg_0_ ( .D(n1002), .CK(clk), .RN(n1092), .Q(DP_x[0]), 
        .QN(n301) );
  DFFR_X1 DP_reg_in_Q_reg_1_ ( .D(n1001), .CK(clk), .RN(n1092), .Q(DP_x[1]), 
        .QN(n300) );
  DFFR_X1 DP_reg_in_Q_reg_2_ ( .D(n1000), .CK(clk), .RN(n1092), .Q(DP_x[2]), 
        .QN(n299) );
  DFFR_X1 DP_reg_in_Q_reg_3_ ( .D(n999), .CK(clk), .RN(n1092), .Q(DP_x[3]), 
        .QN(n298) );
  DFFR_X1 DP_reg_in_Q_reg_4_ ( .D(n998), .CK(clk), .RN(n1092), .Q(DP_x[4]), 
        .QN(n297) );
  DFFR_X1 DP_reg_in_Q_reg_5_ ( .D(n997), .CK(clk), .RN(n1092), .Q(DP_x[5]), 
        .QN(n296) );
  DFFR_X1 DP_reg_in_Q_reg_6_ ( .D(n996), .CK(clk), .RN(n1092), .Q(DP_x[6]), 
        .QN(n295) );
  DFFR_X1 DP_reg_in_Q_reg_7_ ( .D(n995), .CK(clk), .RN(n1092), .Q(DP_x[7]), 
        .QN(n294) );
  DFFR_X1 DP_reg_in_Q_reg_8_ ( .D(n994), .CK(clk), .RN(n1092), .Q(DP_x[8]), 
        .QN(n293) );
  DFFR_X1 DP_reg_in_Q_reg_9_ ( .D(n993), .CK(clk), .RN(n1092), .Q(DP_x[9]), 
        .QN(n292) );
  DFFR_X1 DP_reg_in_Q_reg_10_ ( .D(n992), .CK(clk), .RN(n1092), .Q(DP_x[10]), 
        .QN(n291) );
  DFFR_X1 DP_reg_in_Q_reg_11_ ( .D(n991), .CK(clk), .RN(n1092), .Q(DP_x[11]), 
        .QN(n290) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_0_ ( .D(n990), .CK(clk), .RN(n1093), .Q(
        DP_coeffs_fb_int[23]), .QN(n289) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_1_ ( .D(n989), .CK(clk), .RN(n1093), .Q(
        DP_coeffs_fb_int[22]), .QN(n288) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_2_ ( .D(n988), .CK(clk), .RN(n1093), .Q(
        DP_coeffs_fb_int[21]), .QN(n287) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_3_ ( .D(n987), .CK(clk), .RN(n1093), .Q(
        DP_coeffs_fb_int[20]), .QN(n286) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_4_ ( .D(n986), .CK(clk), .RN(n1093), .Q(
        DP_coeffs_fb_int[19]), .QN(n285) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_5_ ( .D(n985), .CK(clk), .RN(n1093), .Q(
        DP_coeffs_fb_int[18]), .QN(n284) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_6_ ( .D(n984), .CK(clk), .RN(n1093), .Q(
        DP_coeffs_fb_int[17]), .QN(n283) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_7_ ( .D(n983), .CK(clk), .RN(n1093), .Q(
        DP_coeffs_fb_int[16]), .QN(n282) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_8_ ( .D(n982), .CK(clk), .RN(n1093), .Q(
        DP_coeffs_fb_int[15]), .QN(n281) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_9_ ( .D(n981), .CK(clk), .RN(n1093), .Q(
        DP_coeffs_fb_int[14]), .QN(n280) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_10_ ( .D(n980), .CK(clk), .RN(n1093), .Q(
        DP_coeffs_fb_int[13]), .QN(n279) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_11_ ( .D(n979), .CK(clk), .RN(n1093), .Q(
        DP_coeffs_fb_int[12]), .QN(n278) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_12_ ( .D(n978), .CK(clk), .RN(n1094), .Q(
        DP_coeffs_fb_int[11]), .QN(n277) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_13_ ( .D(n977), .CK(clk), .RN(n1094), .Q(
        DP_coeffs_fb_int[10]), .QN(n519) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_14_ ( .D(n976), .CK(clk), .RN(n1094), .Q(
        DP_coeffs_fb_int[9]), .QN(n518) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_15_ ( .D(n975), .CK(clk), .RN(n1094), .Q(
        DP_coeffs_fb_int[8]), .QN(n517) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_16_ ( .D(n974), .CK(clk), .RN(n1094), .Q(
        DP_coeffs_fb_int[7]), .QN(n516) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_17_ ( .D(n973), .CK(clk), .RN(n1094), .Q(
        DP_coeffs_fb_int[6]), .QN(n515) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_18_ ( .D(n972), .CK(clk), .RN(n1094), .Q(
        DP_coeffs_fb_int[5]), .QN(n514) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_19_ ( .D(n971), .CK(clk), .RN(n1094), .Q(
        DP_coeffs_fb_int[4]), .QN(n513) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_20_ ( .D(n970), .CK(clk), .RN(n1094), .Q(
        DP_coeffs_fb_int[3]), .QN(n512) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_21_ ( .D(n969), .CK(clk), .RN(n1094), .Q(
        DP_coeffs_fb_int[2]), .QN(n511) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_22_ ( .D(n968), .CK(clk), .RN(n1094), .Q(
        DP_coeffs_fb_int[1]), .QN(n510) );
  DFFR_X1 DP_reg_coeff_fb_i_1_Q_reg_23_ ( .D(n967), .CK(clk), .RN(n1094), .Q(
        DP_coeffs_fb_int[0]), .QN(n509) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_0_ ( .D(n966), .CK(clk), .RN(n1095), .Q(
        DP_coeffs_fb_int[47]), .QN(n508) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_1_ ( .D(n965), .CK(clk), .RN(n1095), .Q(
        DP_coeffs_fb_int[46]), .QN(n507) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_2_ ( .D(n964), .CK(clk), .RN(n1095), .Q(
        DP_coeffs_fb_int[45]), .QN(n506) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_3_ ( .D(n963), .CK(clk), .RN(n1095), .Q(
        DP_coeffs_fb_int[44]), .QN(n505) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_4_ ( .D(n962), .CK(clk), .RN(n1095), .Q(
        DP_coeffs_fb_int[43]), .QN(n504) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_5_ ( .D(n961), .CK(clk), .RN(n1095), .Q(
        DP_coeffs_fb_int[42]), .QN(n503) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_6_ ( .D(n960), .CK(clk), .RN(n1095), .Q(
        DP_coeffs_fb_int[41]), .QN(n502) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_7_ ( .D(n959), .CK(clk), .RN(n1095), .Q(
        DP_coeffs_fb_int[40]), .QN(n501) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_8_ ( .D(n958), .CK(clk), .RN(n1095), .Q(
        DP_coeffs_fb_int[39]), .QN(n500) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_9_ ( .D(n957), .CK(clk), .RN(n1095), .Q(
        DP_coeffs_fb_int[38]), .QN(n499) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_10_ ( .D(n956), .CK(clk), .RN(n1095), .Q(
        DP_coeffs_fb_int[37]), .QN(n498) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_11_ ( .D(n955), .CK(clk), .RN(n1095), .Q(
        DP_coeffs_fb_int[36]), .QN(n497) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_12_ ( .D(n954), .CK(clk), .RN(n1096), .Q(
        DP_coeffs_fb_int[35]), .QN(n496) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_13_ ( .D(n953), .CK(clk), .RN(n1096), .Q(
        DP_coeffs_fb_int[34]), .QN(n495) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_14_ ( .D(n952), .CK(clk), .RN(n1096), .Q(
        DP_coeffs_fb_int[33]), .QN(n494) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_15_ ( .D(n951), .CK(clk), .RN(n1096), .Q(
        DP_coeffs_fb_int[32]), .QN(n493) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_16_ ( .D(n950), .CK(clk), .RN(n1096), .Q(
        DP_coeffs_fb_int[31]), .QN(n492) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_17_ ( .D(n949), .CK(clk), .RN(n1096), .Q(
        DP_coeffs_fb_int[30]), .QN(n491) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_18_ ( .D(n948), .CK(clk), .RN(n1096), .Q(
        DP_coeffs_fb_int[29]), .QN(n490) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_19_ ( .D(n947), .CK(clk), .RN(n1096), .Q(
        DP_coeffs_fb_int[28]), .QN(n489) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_20_ ( .D(n946), .CK(clk), .RN(n1096), .Q(
        DP_coeffs_fb_int[27]), .QN(n488) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_21_ ( .D(n945), .CK(clk), .RN(n1096), .Q(
        DP_coeffs_fb_int[26]), .QN(n487) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_22_ ( .D(n944), .CK(clk), .RN(n1096), .Q(
        DP_coeffs_fb_int[25]), .QN(n486) );
  DFFR_X1 DP_reg_coeff_fb_i_2_Q_reg_23_ ( .D(n943), .CK(clk), .RN(n1096), .Q(
        DP_coeffs_fb_int[24]), .QN(n485) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_0_ ( .D(n942), .CK(clk), .RN(n1097), .Q(
        DP_coeffs_ff_int[23]), .QN(n484) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_1_ ( .D(n941), .CK(clk), .RN(n1097), .Q(
        DP_coeffs_ff_int[22]), .QN(n483) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_2_ ( .D(n940), .CK(clk), .RN(n1097), .Q(
        DP_coeffs_ff_int[21]), .QN(n482) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_3_ ( .D(n939), .CK(clk), .RN(n1097), .Q(
        DP_coeffs_ff_int[20]), .QN(n481) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_4_ ( .D(n938), .CK(clk), .RN(n1097), .Q(
        DP_coeffs_ff_int[19]), .QN(n480) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_5_ ( .D(n937), .CK(clk), .RN(n1097), .Q(
        DP_coeffs_ff_int[18]), .QN(n479) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_6_ ( .D(n936), .CK(clk), .RN(n1097), .Q(
        DP_coeffs_ff_int[17]), .QN(n478) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_7_ ( .D(n935), .CK(clk), .RN(n1097), .Q(
        DP_coeffs_ff_int[16]), .QN(n477) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_8_ ( .D(n934), .CK(clk), .RN(n1097), .Q(
        DP_coeffs_ff_int[15]), .QN(n476) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_9_ ( .D(n933), .CK(clk), .RN(n1097), .Q(
        DP_coeffs_ff_int[14]), .QN(n475) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_10_ ( .D(n932), .CK(clk), .RN(n1097), .Q(
        DP_coeffs_ff_int[13]), .QN(n474) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_11_ ( .D(n931), .CK(clk), .RN(n1097), .Q(
        DP_coeffs_ff_int[12]), .QN(n473) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_12_ ( .D(n930), .CK(clk), .RN(n1098), .Q(
        DP_coeffs_ff_int[11]), .QN(n472) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_13_ ( .D(n929), .CK(clk), .RN(n1098), .Q(
        DP_coeffs_ff_int[10]), .QN(n471) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_14_ ( .D(n928), .CK(clk), .RN(n1098), .Q(
        DP_coeffs_ff_int[9]), .QN(n470) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_15_ ( .D(n927), .CK(clk), .RN(n1098), .Q(
        DP_coeffs_ff_int[8]), .QN(n469) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_16_ ( .D(n926), .CK(clk), .RN(n1098), .Q(
        DP_coeffs_ff_int[7]), .QN(n468) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_17_ ( .D(n925), .CK(clk), .RN(n1098), .Q(
        DP_coeffs_ff_int[6]), .QN(n467) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_18_ ( .D(n924), .CK(clk), .RN(n1098), .Q(
        DP_coeffs_ff_int[5]), .QN(n466) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_19_ ( .D(n923), .CK(clk), .RN(n1098), .Q(
        DP_coeffs_ff_int[4]), .QN(n465) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_20_ ( .D(n922), .CK(clk), .RN(n1098), .Q(
        DP_coeffs_ff_int[3]), .QN(n464) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_21_ ( .D(n921), .CK(clk), .RN(n1098), .Q(
        DP_coeffs_ff_int[2]), .QN(n463) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_22_ ( .D(n920), .CK(clk), .RN(n1098), .Q(
        DP_coeffs_ff_int[1]), .QN(n462) );
  DFFR_X1 DP_reg_b_i_0_Q_reg_23_ ( .D(n919), .CK(clk), .RN(n1098), .Q(
        DP_coeffs_ff_int[0]), .QN(n461) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_0_ ( .D(n918), .CK(clk), .RN(n1099), .Q(
        DP_coeffs_ff_int[47]), .QN(n460) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_1_ ( .D(n917), .CK(clk), .RN(n1099), .Q(
        DP_coeffs_ff_int[46]), .QN(n459) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_2_ ( .D(n916), .CK(clk), .RN(n1099), .Q(
        DP_coeffs_ff_int[45]), .QN(n458) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_3_ ( .D(n915), .CK(clk), .RN(n1099), .Q(
        DP_coeffs_ff_int[44]), .QN(n457) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_4_ ( .D(n914), .CK(clk), .RN(n1099), .Q(
        DP_coeffs_ff_int[43]), .QN(n456) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_5_ ( .D(n913), .CK(clk), .RN(n1099), .Q(
        DP_coeffs_ff_int[42]), .QN(n455) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_6_ ( .D(n912), .CK(clk), .RN(n1099), .Q(
        DP_coeffs_ff_int[41]), .QN(n454) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_7_ ( .D(n911), .CK(clk), .RN(n1099), .Q(
        DP_coeffs_ff_int[40]), .QN(n453) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_8_ ( .D(n910), .CK(clk), .RN(n1099), .Q(
        DP_coeffs_ff_int[39]), .QN(n452) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_9_ ( .D(n909), .CK(clk), .RN(n1099), .Q(
        DP_coeffs_ff_int[38]), .QN(n451) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_10_ ( .D(n908), .CK(clk), .RN(n1099), .Q(
        DP_coeffs_ff_int[37]), .QN(n450) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_11_ ( .D(n907), .CK(clk), .RN(n1099), .Q(
        DP_coeffs_ff_int[36]), .QN(n449) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_12_ ( .D(n906), .CK(clk), .RN(n1100), .Q(
        DP_coeffs_ff_int[35]), .QN(n448) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_13_ ( .D(n905), .CK(clk), .RN(n1100), .Q(
        DP_coeffs_ff_int[34]), .QN(n447) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_14_ ( .D(n904), .CK(clk), .RN(n1100), .Q(
        DP_coeffs_ff_int[33]), .QN(n446) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_15_ ( .D(n903), .CK(clk), .RN(n1100), .Q(
        DP_coeffs_ff_int[32]), .QN(n445) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_16_ ( .D(n902), .CK(clk), .RN(n1100), .Q(
        DP_coeffs_ff_int[31]), .QN(n444) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_17_ ( .D(n901), .CK(clk), .RN(n1100), .Q(
        DP_coeffs_ff_int[30]), .QN(n443) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_18_ ( .D(n900), .CK(clk), .RN(n1100), .Q(
        DP_coeffs_ff_int[29]), .QN(n442) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_19_ ( .D(n899), .CK(clk), .RN(n1100), .Q(
        DP_coeffs_ff_int[28]), .QN(n441) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_20_ ( .D(n898), .CK(clk), .RN(n1100), .Q(
        DP_coeffs_ff_int[27]), .QN(n440) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_21_ ( .D(n897), .CK(clk), .RN(n1100), .Q(
        DP_coeffs_ff_int[26]), .QN(n439) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_22_ ( .D(n896), .CK(clk), .RN(n1100), .Q(
        DP_coeffs_ff_int[25]), .QN(n438) );
  DFFR_X1 DP_reg_b_i_1_Q_reg_23_ ( .D(n895), .CK(clk), .RN(n1100), .Q(
        DP_coeffs_ff_int[24]), .QN(n437) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_0_ ( .D(n894), .CK(clk), .RN(n1101), .Q(
        DP_coeffs_ff_int[71]), .QN(n436) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_1_ ( .D(n893), .CK(clk), .RN(n1101), .Q(
        DP_coeffs_ff_int[70]), .QN(n435) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_2_ ( .D(n892), .CK(clk), .RN(n1101), .Q(
        DP_coeffs_ff_int[69]), .QN(n434) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_3_ ( .D(n891), .CK(clk), .RN(n1101), .Q(
        DP_coeffs_ff_int[68]), .QN(n433) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_4_ ( .D(n890), .CK(clk), .RN(n1101), .Q(
        DP_coeffs_ff_int[67]), .QN(n432) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_5_ ( .D(n889), .CK(clk), .RN(n1101), .Q(
        DP_coeffs_ff_int[66]), .QN(n431) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_6_ ( .D(n888), .CK(clk), .RN(n1101), .Q(
        DP_coeffs_ff_int[65]), .QN(n430) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_7_ ( .D(n887), .CK(clk), .RN(n1101), .Q(
        DP_coeffs_ff_int[64]), .QN(n429) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_8_ ( .D(n886), .CK(clk), .RN(n1101), .Q(
        DP_coeffs_ff_int[63]), .QN(n428) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_9_ ( .D(n885), .CK(clk), .RN(n1101), .Q(
        DP_coeffs_ff_int[62]), .QN(n427) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_10_ ( .D(n884), .CK(clk), .RN(n1101), .Q(
        DP_coeffs_ff_int[61]), .QN(n426) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_11_ ( .D(n883), .CK(clk), .RN(n1101), .Q(
        DP_coeffs_ff_int[60]), .QN(n425) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_12_ ( .D(n882), .CK(clk), .RN(n1102), .Q(
        DP_coeffs_ff_int[59]), .QN(n424) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_13_ ( .D(n881), .CK(clk), .RN(n1102), .Q(
        DP_coeffs_ff_int[58]), .QN(n423) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_14_ ( .D(n880), .CK(clk), .RN(n1102), .Q(
        DP_coeffs_ff_int[57]), .QN(n422) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_15_ ( .D(n879), .CK(clk), .RN(n1102), .Q(
        DP_coeffs_ff_int[56]), .QN(n421) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_16_ ( .D(n878), .CK(clk), .RN(n1102), .Q(
        DP_coeffs_ff_int[55]), .QN(n420) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_17_ ( .D(n877), .CK(clk), .RN(n1102), .Q(
        DP_coeffs_ff_int[54]), .QN(n419) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_18_ ( .D(n876), .CK(clk), .RN(n1102), .Q(
        DP_coeffs_ff_int[53]), .QN(n418) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_19_ ( .D(n875), .CK(clk), .RN(n1102), .Q(
        DP_coeffs_ff_int[52]), .QN(n417) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_20_ ( .D(n874), .CK(clk), .RN(n1102), .Q(
        DP_coeffs_ff_int[51]), .QN(n416) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_21_ ( .D(n873), .CK(clk), .RN(n1102), .Q(
        DP_coeffs_ff_int[50]), .QN(n415) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_22_ ( .D(n872), .CK(clk), .RN(n1102), .Q(
        DP_coeffs_ff_int[49]), .QN(n414) );
  DFFR_X1 DP_reg_b_i_2_Q_reg_23_ ( .D(n871), .CK(clk), .RN(n1102), .Q(
        DP_coeffs_ff_int[48]), .QN(n413) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_0_ ( .D(n870), .CK(clk), .RN(n1103), .Q(
        DP_coeffs_ff_int[95]), .QN(n412) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_1_ ( .D(n869), .CK(clk), .RN(n1103), .Q(
        DP_coeffs_ff_int[94]), .QN(n411) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_2_ ( .D(n868), .CK(clk), .RN(n1103), .Q(
        DP_coeffs_ff_int[93]), .QN(n410) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_3_ ( .D(n867), .CK(clk), .RN(n1103), .Q(
        DP_coeffs_ff_int[92]), .QN(n409) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_4_ ( .D(n866), .CK(clk), .RN(n1103), .Q(
        DP_coeffs_ff_int[91]), .QN(n408) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_5_ ( .D(n865), .CK(clk), .RN(n1103), .Q(
        DP_coeffs_ff_int[90]), .QN(n407) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_6_ ( .D(n864), .CK(clk), .RN(n1103), .Q(
        DP_coeffs_ff_int[89]), .QN(n406) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_7_ ( .D(n863), .CK(clk), .RN(n1103), .Q(
        DP_coeffs_ff_int[88]), .QN(n405) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_8_ ( .D(n862), .CK(clk), .RN(n1103), .Q(
        DP_coeffs_ff_int[87]), .QN(n404) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_9_ ( .D(n861), .CK(clk), .RN(n1103), .Q(
        DP_coeffs_ff_int[86]), .QN(n403) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_10_ ( .D(n860), .CK(clk), .RN(n1103), .Q(
        DP_coeffs_ff_int[85]), .QN(n402) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_11_ ( .D(n859), .CK(clk), .RN(n1103), .Q(
        DP_coeffs_ff_int[84]), .QN(n401) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_12_ ( .D(n858), .CK(clk), .RN(n1104), .Q(
        DP_coeffs_ff_int[83]), .QN(n400) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_13_ ( .D(n857), .CK(clk), .RN(n1104), .Q(
        DP_coeffs_ff_int[82]), .QN(n399) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_14_ ( .D(n856), .CK(clk), .RN(n1104), .Q(
        DP_coeffs_ff_int[81]), .QN(n398) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_15_ ( .D(n855), .CK(clk), .RN(n1104), .Q(
        DP_coeffs_ff_int[80]), .QN(n397) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_16_ ( .D(n854), .CK(clk), .RN(n1104), .Q(
        DP_coeffs_ff_int[79]), .QN(n396) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_17_ ( .D(n853), .CK(clk), .RN(n1104), .Q(
        DP_coeffs_ff_int[78]), .QN(n395) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_18_ ( .D(n852), .CK(clk), .RN(n1104), .Q(
        DP_coeffs_ff_int[77]), .QN(n394) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_19_ ( .D(n851), .CK(clk), .RN(n1104), .Q(
        DP_coeffs_ff_int[76]), .QN(n393) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_20_ ( .D(n850), .CK(clk), .RN(n1104), .Q(
        DP_coeffs_ff_int[75]), .QN(n392) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_21_ ( .D(n849), .CK(clk), .RN(n1104), .Q(
        DP_coeffs_ff_int[74]), .QN(n391) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_22_ ( .D(n848), .CK(clk), .RN(n1104), .Q(
        DP_coeffs_ff_int[73]), .QN(n390) );
  DFFR_X1 DP_reg_b_i_3_Q_reg_23_ ( .D(n847), .CK(clk), .RN(n1104), .Q(
        DP_coeffs_ff_int[72]), .QN(n389) );
  DFFR_X1 CU_presentState_reg_1_ ( .D(n1033), .CK(clk), .RN(n1105), .Q(
        delayed_controls_0__1_) );
  DFFR_X1 DP_reg_sw1_Q_reg_0_ ( .D(n846), .CK(clk), .RN(n1105), .Q(DP_sw1_0_), 
        .QN(n1003) );
  DFFR_X1 DP_reg_pipe02_Q_reg_0_ ( .D(DP_sw1_0_), .CK(clk), .RN(n1105), .Q(
        DP_pipe02[0]) );
  DFFR_X1 DP_reg_ret1_Q_reg_0_ ( .D(DP_sw1_coeff_ret1[0]), .CK(clk), .RN(n1105), .Q(DP_ret1[0]) );
  DFFR_X1 DP_reg_ret1_Q_reg_1_ ( .D(DP_sw1_coeff_ret1[1]), .CK(clk), .RN(n1105), .Q(DP_ret1[1]) );
  DFFR_X1 DP_reg_ret1_Q_reg_2_ ( .D(DP_sw1_coeff_ret1[2]), .CK(clk), .RN(n1105), .Q(DP_ret1[2]) );
  DFFR_X1 DP_reg_ret1_Q_reg_3_ ( .D(DP_sw1_coeff_ret1[3]), .CK(clk), .RN(n1105), .Q(DP_ret1[3]) );
  DFFR_X1 DP_reg_ret1_Q_reg_4_ ( .D(DP_sw1_coeff_ret1[4]), .CK(clk), .RN(n1105), .Q(DP_ret1[4]) );
  DFFR_X1 DP_reg_ret1_Q_reg_5_ ( .D(DP_sw1_coeff_ret1[5]), .CK(clk), .RN(n1105), .Q(DP_ret1[5]) );
  DFFR_X1 DP_reg_ret1_Q_reg_6_ ( .D(DP_sw1_coeff_ret1[6]), .CK(clk), .RN(n1105), .Q(DP_ret1[6]) );
  DFFR_X1 DP_reg_ret1_Q_reg_7_ ( .D(DP_sw1_coeff_ret1[7]), .CK(clk), .RN(n1105), .Q(DP_ret1[7]) );
  DFFR_X1 DP_reg_ret1_Q_reg_8_ ( .D(DP_sw1_coeff_ret1[8]), .CK(clk), .RN(n1105), .Q(DP_ret1[8]) );
  DFFR_X1 DP_reg_ret1_Q_reg_9_ ( .D(DP_sw1_coeff_ret1[9]), .CK(clk), .RN(n1106), .Q(DP_ret1[9]) );
  DFFR_X1 DP_reg_ret1_Q_reg_10_ ( .D(DP_sw1_coeff_ret1[10]), .CK(clk), .RN(
        n1106), .Q(DP_ret1[10]) );
  DFFR_X1 DP_reg_ret1_Q_reg_11_ ( .D(DP_sw1_coeff_ret1[11]), .CK(clk), .RN(
        n1106), .Q(DP_ret1[11]) );
  DFFR_X1 DP_reg_ret1_Q_reg_12_ ( .D(DP_sw1_coeff_ret1[12]), .CK(clk), .RN(
        n1106), .Q(DP_ret1[12]) );
  DFFR_X1 DP_reg_ret1_Q_reg_13_ ( .D(DP_sw1_coeff_ret1[13]), .CK(clk), .RN(
        n1106), .Q(DP_ret1[13]) );
  DFFR_X1 DP_reg_ret1_Q_reg_14_ ( .D(DP_sw1_coeff_ret1[14]), .CK(clk), .RN(
        n1106), .Q(DP_ret1[14]) );
  DFFR_X1 DP_reg_ret1_Q_reg_15_ ( .D(DP_sw1_coeff_ret1[15]), .CK(clk), .RN(
        n1106), .Q(DP_ret1[15]) );
  DFFR_X1 DP_reg_ret1_Q_reg_16_ ( .D(DP_sw1_coeff_ret1[16]), .CK(clk), .RN(
        n1106), .Q(DP_ret1[16]) );
  DFFR_X1 DP_reg_ret1_Q_reg_17_ ( .D(DP_sw1_coeff_ret1[17]), .CK(clk), .RN(
        n1106), .Q(DP_ret1[17]) );
  DFFR_X1 DP_reg_ret1_Q_reg_18_ ( .D(DP_sw1_coeff_ret1[18]), .CK(clk), .RN(
        n1106), .Q(DP_ret1[18]) );
  DFFR_X1 DP_reg_ret1_Q_reg_19_ ( .D(DP_sw1_coeff_ret1[19]), .CK(clk), .RN(
        n1106), .Q(DP_ret1[19]) );
  DFFR_X1 DP_reg_ret1_Q_reg_20_ ( .D(DP_sw1_coeff_ret1[20]), .CK(clk), .RN(
        n1106), .Q(DP_ret1[20]) );
  DFFR_X1 DP_reg_ret1_Q_reg_21_ ( .D(DP_sw1_coeff_ret1[21]), .CK(clk), .RN(
        n1107), .Q(DP_ret1[21]) );
  DFFR_X1 DP_reg_ret1_Q_reg_22_ ( .D(DP_sw1_coeff_ret1[22]), .CK(clk), .RN(
        n1107), .Q(DP_ret1[22]) );
  DFFR_X1 DP_reg_ret1_Q_reg_23_ ( .D(DP_sw1_coeff_ret1[23]), .CK(clk), .RN(
        n1107), .Q(DP_ret1[23]) );
  DFFR_X1 DP_reg_sw0_Q_reg_0_ ( .D(n820), .CK(clk), .RN(n1107), .Q(DP_sw0_0_), 
        .QN(n1026) );
  DFFR_X1 DP_reg_pipe01_Q_reg_0_ ( .D(DP_sw0_0_), .CK(clk), .RN(n1107), .Q(
        DP_pipe01[0]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_0_ ( .D(DP_w_0_), .CK(clk), .RN(n1107), .Q(
        DP_pipe00[0]) );
  DFFR_X1 DP_reg_sw0_Q_reg_1_ ( .D(n817), .CK(clk), .RN(n1107), .Q(DP_sw0_1_)
         );
  DFFR_X1 DP_reg_sw1_Q_reg_1_ ( .D(n816), .CK(clk), .RN(n1107), .Q(DP_sw1_1_), 
        .QN(n1025) );
  DFFR_X1 DP_reg_pipe02_Q_reg_1_ ( .D(DP_sw1_1_), .CK(clk), .RN(n1107), .Q(
        DP_pipe02[1]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_1_ ( .D(DP_sw0_1_), .CK(clk), .RN(n1107), .Q(
        DP_pipe01[1]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_1_ ( .D(DP_w_1_), .CK(clk), .RN(n1107), .Q(
        DP_pipe00[1]) );
  DFFR_X1 DP_reg_sw0_Q_reg_2_ ( .D(n812), .CK(clk), .RN(n1107), .Q(DP_sw0_2_)
         );
  DFFR_X1 DP_reg_sw1_Q_reg_2_ ( .D(n811), .CK(clk), .RN(n1108), .Q(DP_sw1_2_), 
        .QN(n1007) );
  DFFR_X1 DP_reg_pipe02_Q_reg_2_ ( .D(DP_sw1_2_), .CK(clk), .RN(n1108), .Q(
        DP_pipe02[2]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_2_ ( .D(DP_sw0_2_), .CK(clk), .RN(n1108), .Q(
        DP_pipe01[2]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_2_ ( .D(DP_w_2_), .CK(clk), .RN(n1108), .Q(
        DP_pipe00[2]) );
  DFFR_X1 DP_reg_sw0_Q_reg_3_ ( .D(n807), .CK(clk), .RN(n1108), .Q(DP_sw0_3_)
         );
  DFFR_X1 DP_reg_sw1_Q_reg_3_ ( .D(n806), .CK(clk), .RN(n1108), .Q(DP_sw1_3_), 
        .QN(n1008) );
  DFFR_X1 DP_reg_pipe02_Q_reg_3_ ( .D(DP_sw1_3_), .CK(clk), .RN(n1108), .Q(
        DP_pipe02[3]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_3_ ( .D(DP_sw0_3_), .CK(clk), .RN(n1108), .Q(
        DP_pipe01[3]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_3_ ( .D(DP_w_3_), .CK(clk), .RN(n1108), .Q(
        DP_pipe00[3]) );
  DFFR_X1 DP_reg_sw0_Q_reg_4_ ( .D(n802), .CK(clk), .RN(n1108), .Q(DP_sw0_4_)
         );
  DFFR_X1 DP_reg_sw1_Q_reg_4_ ( .D(n801), .CK(clk), .RN(n1108), .Q(DP_sw1_4_), 
        .QN(n1009) );
  DFFR_X1 DP_reg_pipe02_Q_reg_4_ ( .D(DP_sw1_4_), .CK(clk), .RN(n1108), .Q(
        DP_pipe02[4]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_4_ ( .D(DP_sw0_4_), .CK(clk), .RN(n1109), .Q(
        DP_pipe01[4]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_4_ ( .D(DP_w_4_), .CK(clk), .RN(n1109), .Q(
        DP_pipe00[4]) );
  DFFR_X1 DP_reg_sw0_Q_reg_5_ ( .D(n797), .CK(clk), .RN(n1109), .Q(DP_sw0_5_)
         );
  DFFR_X1 DP_reg_sw1_Q_reg_5_ ( .D(n796), .CK(clk), .RN(n1109), .Q(DP_sw1_5_), 
        .QN(n1010) );
  DFFR_X1 DP_reg_pipe02_Q_reg_5_ ( .D(DP_sw1_5_), .CK(clk), .RN(n1109), .Q(
        DP_pipe02[5]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_5_ ( .D(DP_sw0_5_), .CK(clk), .RN(n1109), .Q(
        DP_pipe01[5]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_5_ ( .D(DP_w_5_), .CK(clk), .RN(n1109), .Q(
        DP_pipe00[5]) );
  DFFR_X1 DP_reg_sw0_Q_reg_6_ ( .D(n792), .CK(clk), .RN(n1109), .Q(DP_sw0_6_)
         );
  DFFR_X1 DP_reg_sw1_Q_reg_6_ ( .D(n791), .CK(clk), .RN(n1109), .Q(DP_sw1_6_), 
        .QN(n1011) );
  DFFR_X1 DP_reg_pipe02_Q_reg_6_ ( .D(DP_sw1_6_), .CK(clk), .RN(n1109), .Q(
        DP_pipe02[6]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_6_ ( .D(DP_sw0_6_), .CK(clk), .RN(n1109), .Q(
        DP_pipe01[6]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_6_ ( .D(DP_w_6_), .CK(clk), .RN(n1109), .Q(
        DP_pipe00[6]) );
  DFFR_X1 DP_reg_sw0_Q_reg_7_ ( .D(n787), .CK(clk), .RN(n1110), .Q(DP_sw0_7_)
         );
  DFFR_X1 DP_reg_sw1_Q_reg_7_ ( .D(n786), .CK(clk), .RN(n1110), .Q(DP_sw1_7_), 
        .QN(n1012) );
  DFFR_X1 DP_reg_pipe02_Q_reg_7_ ( .D(DP_sw1_7_), .CK(clk), .RN(n1110), .Q(
        DP_pipe02[7]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_7_ ( .D(DP_sw0_7_), .CK(clk), .RN(n1110), .Q(
        DP_pipe01[7]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_7_ ( .D(DP_w_7_), .CK(clk), .RN(n1110), .Q(
        DP_pipe00[7]) );
  DFFR_X1 DP_reg_sw0_Q_reg_8_ ( .D(n782), .CK(clk), .RN(n1110), .Q(DP_sw0_8_)
         );
  DFFR_X1 DP_reg_sw1_Q_reg_8_ ( .D(n781), .CK(clk), .RN(n1110), .Q(DP_sw1_8_), 
        .QN(n1013) );
  DFFR_X1 DP_reg_pipe02_Q_reg_8_ ( .D(DP_sw1_8_), .CK(clk), .RN(n1110), .Q(
        DP_pipe02[8]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_8_ ( .D(DP_sw0_8_), .CK(clk), .RN(n1110), .Q(
        DP_pipe01[8]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_8_ ( .D(DP_w_8_), .CK(clk), .RN(n1110), .Q(
        DP_pipe00[8]) );
  DFFR_X1 DP_reg_sw0_Q_reg_9_ ( .D(n777), .CK(clk), .RN(n1110), .Q(DP_sw0_9_)
         );
  DFFR_X1 DP_reg_sw1_Q_reg_9_ ( .D(n776), .CK(clk), .RN(n1110), .Q(DP_sw1_9_), 
        .QN(n1014) );
  DFFR_X1 DP_reg_pipe02_Q_reg_9_ ( .D(DP_sw1_9_), .CK(clk), .RN(n1111), .Q(
        DP_pipe02[9]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_9_ ( .D(DP_sw0_9_), .CK(clk), .RN(n1111), .Q(
        DP_pipe01[9]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_9_ ( .D(DP_w_9_), .CK(clk), .RN(n1111), .Q(
        DP_pipe00[9]) );
  DFFR_X1 DP_reg_sw0_Q_reg_10_ ( .D(n772), .CK(clk), .RN(n1111), .Q(DP_sw0_10_) );
  DFFR_X1 DP_reg_sw1_Q_reg_10_ ( .D(n771), .CK(clk), .RN(n1111), .Q(DP_sw1_10_), .QN(n1015) );
  DFFR_X1 DP_reg_pipe02_Q_reg_10_ ( .D(DP_sw1_10_), .CK(clk), .RN(n1111), .Q(
        DP_pipe02[10]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_10_ ( .D(DP_sw0_10_), .CK(clk), .RN(n1111), .Q(
        DP_pipe01[10]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_10_ ( .D(DP_w_10_), .CK(clk), .RN(n1111), .Q(
        DP_pipe00[10]) );
  DFFR_X1 DP_reg_sw0_Q_reg_11_ ( .D(n767), .CK(clk), .RN(n1111), .Q(DP_sw0_11_) );
  DFFR_X1 DP_reg_sw1_Q_reg_11_ ( .D(n766), .CK(clk), .RN(n1111), .Q(DP_sw1_11_), .QN(n1016) );
  DFFR_X1 DP_reg_pipe02_Q_reg_11_ ( .D(DP_sw1_11_), .CK(clk), .RN(n1111), .Q(
        DP_pipe02[11]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_11_ ( .D(DP_sw0_11_), .CK(clk), .RN(n1111), .Q(
        DP_pipe01[11]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_11_ ( .D(DP_w_11_), .CK(clk), .RN(n1112), .Q(
        DP_pipe00[11]) );
  DFFR_X1 DP_reg_sw0_Q_reg_12_ ( .D(n762), .CK(clk), .RN(n1112), .Q(DP_sw0_12_) );
  DFFR_X1 DP_reg_sw1_Q_reg_12_ ( .D(n761), .CK(clk), .RN(n1112), .Q(DP_sw1_12_), .QN(n1017) );
  DFFR_X1 DP_reg_pipe02_Q_reg_12_ ( .D(DP_sw1_12_), .CK(clk), .RN(n1112), .Q(
        DP_pipe02[12]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_12_ ( .D(DP_sw0_12_), .CK(clk), .RN(n1112), .Q(
        DP_pipe01[12]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_12_ ( .D(DP_w_12_), .CK(clk), .RN(n1112), .Q(
        DP_pipe00[12]) );
  DFFR_X1 DP_reg_sw0_Q_reg_13_ ( .D(n757), .CK(clk), .RN(n1112), .Q(DP_sw0_13_) );
  DFFR_X1 DP_reg_sw1_Q_reg_13_ ( .D(n756), .CK(clk), .RN(n1112), .Q(DP_sw1_13_), .QN(n1018) );
  DFFR_X1 DP_reg_pipe02_Q_reg_13_ ( .D(DP_sw1_13_), .CK(clk), .RN(n1112), .Q(
        DP_pipe02[13]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_13_ ( .D(DP_sw0_13_), .CK(clk), .RN(n1112), .Q(
        DP_pipe01[13]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_13_ ( .D(DP_w_13_), .CK(clk), .RN(n1112), .Q(
        DP_pipe00[13]) );
  DFFR_X1 DP_reg_sw0_Q_reg_14_ ( .D(n752), .CK(clk), .RN(n1112), .Q(DP_sw0_14_) );
  DFFR_X1 DP_reg_sw1_Q_reg_14_ ( .D(n751), .CK(clk), .RN(n1113), .Q(DP_sw1_14_), .QN(n1019) );
  DFFR_X1 DP_reg_pipe02_Q_reg_14_ ( .D(DP_sw1_14_), .CK(clk), .RN(n1113), .Q(
        DP_pipe02[14]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_14_ ( .D(DP_sw0_14_), .CK(clk), .RN(n1113), .Q(
        DP_pipe01[14]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_14_ ( .D(DP_w_14_), .CK(clk), .RN(n1113), .Q(
        DP_pipe00[14]) );
  DFFR_X1 DP_reg_sw0_Q_reg_15_ ( .D(n747), .CK(clk), .RN(n1113), .Q(DP_sw0_15_) );
  DFFR_X1 DP_reg_sw1_Q_reg_15_ ( .D(n746), .CK(clk), .RN(n1113), .Q(DP_sw1_15_), .QN(n1020) );
  DFFR_X1 DP_reg_pipe02_Q_reg_15_ ( .D(DP_sw1_15_), .CK(clk), .RN(n1113), .Q(
        DP_pipe02[15]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_15_ ( .D(DP_sw0_15_), .CK(clk), .RN(n1113), .Q(
        DP_pipe01[15]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_15_ ( .D(DP_w_15_), .CK(clk), .RN(n1113), .Q(
        DP_pipe00[15]) );
  DFFR_X1 DP_reg_sw0_Q_reg_16_ ( .D(n742), .CK(clk), .RN(n1113), .Q(DP_sw0_16_) );
  DFFR_X1 DP_reg_sw1_Q_reg_16_ ( .D(n741), .CK(clk), .RN(n1113), .Q(DP_sw1_16_), .QN(n1021) );
  DFFR_X1 DP_reg_pipe02_Q_reg_16_ ( .D(DP_sw1_16_), .CK(clk), .RN(n1113), .Q(
        DP_pipe02[16]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_16_ ( .D(DP_sw0_16_), .CK(clk), .RN(n1114), .Q(
        DP_pipe01[16]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_16_ ( .D(DP_w_16_), .CK(clk), .RN(n1114), .Q(
        DP_pipe00[16]) );
  DFFR_X1 DP_reg_sw0_Q_reg_17_ ( .D(n737), .CK(clk), .RN(n1114), .Q(DP_sw0_17_) );
  DFFR_X1 DP_reg_sw1_Q_reg_17_ ( .D(n736), .CK(clk), .RN(n1114), .Q(DP_sw1_17_), .QN(n1022) );
  DFFR_X1 DP_reg_pipe02_Q_reg_17_ ( .D(DP_sw1_17_), .CK(clk), .RN(n1114), .Q(
        DP_pipe02[17]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_17_ ( .D(DP_sw0_17_), .CK(clk), .RN(n1114), .Q(
        DP_pipe01[17]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_17_ ( .D(DP_w_17_), .CK(clk), .RN(n1114), .Q(
        DP_pipe00[17]) );
  DFFR_X1 DP_reg_sw0_Q_reg_18_ ( .D(n732), .CK(clk), .RN(n1114), .Q(DP_sw0_18_) );
  DFFR_X1 DP_reg_sw1_Q_reg_18_ ( .D(n731), .CK(clk), .RN(n1114), .Q(DP_sw1_18_), .QN(n1023) );
  DFFR_X1 DP_reg_pipe02_Q_reg_18_ ( .D(DP_sw1_18_), .CK(clk), .RN(n1114), .Q(
        DP_pipe02[18]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_18_ ( .D(DP_sw0_18_), .CK(clk), .RN(n1114), .Q(
        DP_pipe01[18]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_18_ ( .D(DP_w_18_), .CK(clk), .RN(n1114), .Q(
        DP_pipe00[18]) );
  DFFR_X1 DP_reg_sw0_Q_reg_19_ ( .D(n727), .CK(clk), .RN(n1115), .Q(DP_sw0_19_) );
  DFFR_X1 DP_reg_sw1_Q_reg_19_ ( .D(n726), .CK(clk), .RN(n1115), .Q(DP_sw1_19_), .QN(n1024) );
  DFFR_X1 DP_reg_pipe02_Q_reg_19_ ( .D(DP_sw1_19_), .CK(clk), .RN(n1115), .Q(
        DP_pipe02[19]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_19_ ( .D(DP_sw0_19_), .CK(clk), .RN(n1115), .Q(
        DP_pipe01[19]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_19_ ( .D(DP_w_19_), .CK(clk), .RN(n1115), .Q(
        DP_pipe00[19]) );
  DFFR_X1 DP_reg_sw0_Q_reg_20_ ( .D(n722), .CK(clk), .RN(n1115), .Q(DP_sw0_20_) );
  DFFR_X1 DP_reg_sw1_Q_reg_20_ ( .D(n721), .CK(clk), .RN(n1115), .Q(DP_sw1_20_), .QN(n1005) );
  DFFR_X1 DP_reg_pipe02_Q_reg_20_ ( .D(DP_sw1_20_), .CK(clk), .RN(n1115), .Q(
        DP_pipe02[20]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_20_ ( .D(DP_sw0_20_), .CK(clk), .RN(n1115), .Q(
        DP_pipe01[20]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_20_ ( .D(DP_w_20_), .CK(clk), .RN(n1115), .Q(
        DP_pipe00[20]) );
  DFFR_X1 DP_reg_sw0_Q_reg_21_ ( .D(n717), .CK(clk), .RN(n1115), .Q(DP_sw0_21_) );
  DFFR_X1 DP_reg_sw1_Q_reg_21_ ( .D(n716), .CK(clk), .RN(n1115), .Q(DP_sw1_21_), .QN(n1006) );
  DFFR_X1 DP_reg_pipe02_Q_reg_21_ ( .D(DP_sw1_21_), .CK(clk), .RN(n1116), .Q(
        DP_pipe02[21]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_21_ ( .D(DP_sw0_21_), .CK(clk), .RN(n1116), .Q(
        DP_pipe01[21]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_21_ ( .D(DP_w_21_), .CK(clk), .RN(n1116), .Q(
        DP_pipe00[21]) );
  DFFR_X1 DP_reg_sw0_Q_reg_22_ ( .D(n712), .CK(clk), .RN(n1116), .Q(DP_sw0_22_) );
  DFFR_X1 DP_reg_sw1_Q_reg_22_ ( .D(n711), .CK(clk), .RN(n1116), .Q(DP_sw1_22_), .QN(n1004) );
  DFFR_X1 DP_reg_pipe02_Q_reg_22_ ( .D(DP_sw1_22_), .CK(clk), .RN(n1116), .Q(
        DP_pipe02[22]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_22_ ( .D(DP_sw0_22_), .CK(clk), .RN(n1116), .Q(
        DP_pipe01[22]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_22_ ( .D(DP_w_22_), .CK(clk), .RN(n1116), .Q(
        DP_pipe00[22]) );
  DFFR_X1 DP_reg_sw0_Q_reg_23_ ( .D(n707), .CK(clk), .RN(n1116), .Q(DP_sw0_23_) );
  DFFR_X1 DP_reg_sw1_Q_reg_23_ ( .D(n706), .CK(clk), .RN(n1116), .Q(DP_sw1_23_) );
  DFFR_X1 DP_reg_pipe02_Q_reg_23_ ( .D(n1058), .CK(clk), .RN(n1116), .Q(
        DP_pipe02[23]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_0_ ( .D(DP_pipe0_coeff_pipe02[0]), .CK(clk), 
        .RN(n1116), .Q(DP_pipe12[0]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_1_ ( .D(DP_pipe0_coeff_pipe02[1]), .CK(clk), 
        .RN(n1117), .Q(DP_pipe12[1]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_2_ ( .D(DP_pipe0_coeff_pipe02[2]), .CK(clk), 
        .RN(n1117), .Q(DP_pipe12[2]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_3_ ( .D(DP_pipe0_coeff_pipe02[3]), .CK(clk), 
        .RN(n1117), .Q(DP_pipe12[3]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_4_ ( .D(DP_pipe0_coeff_pipe02[4]), .CK(clk), 
        .RN(n1117), .Q(DP_pipe12[4]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_5_ ( .D(DP_pipe0_coeff_pipe02[5]), .CK(clk), 
        .RN(n1117), .Q(DP_pipe12[5]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_6_ ( .D(DP_pipe0_coeff_pipe02[6]), .CK(clk), 
        .RN(n1117), .Q(DP_pipe12[6]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_7_ ( .D(DP_pipe0_coeff_pipe02[7]), .CK(clk), 
        .RN(n1117), .Q(DP_pipe12[7]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_8_ ( .D(DP_pipe0_coeff_pipe02[8]), .CK(clk), 
        .RN(n1117), .Q(DP_pipe12[8]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_9_ ( .D(DP_pipe0_coeff_pipe02[9]), .CK(clk), 
        .RN(n1117), .Q(DP_pipe12[9]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_10_ ( .D(DP_pipe0_coeff_pipe02[10]), .CK(clk), 
        .RN(n1117), .Q(DP_pipe12[10]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_11_ ( .D(DP_pipe0_coeff_pipe02[11]), .CK(clk), 
        .RN(n1117), .Q(DP_pipe12[11]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_12_ ( .D(DP_pipe0_coeff_pipe02[12]), .CK(clk), 
        .RN(n1117), .Q(DP_pipe12[12]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_13_ ( .D(DP_pipe0_coeff_pipe02[13]), .CK(clk), 
        .RN(n1118), .Q(DP_pipe12[13]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_14_ ( .D(DP_pipe0_coeff_pipe02[14]), .CK(clk), 
        .RN(n1118), .Q(DP_pipe12[14]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_15_ ( .D(DP_pipe0_coeff_pipe02[15]), .CK(clk), 
        .RN(n1118), .Q(DP_pipe12[15]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_16_ ( .D(DP_pipe0_coeff_pipe02[16]), .CK(clk), 
        .RN(n1118), .Q(DP_pipe12[16]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_17_ ( .D(DP_pipe0_coeff_pipe02[17]), .CK(clk), 
        .RN(n1118), .Q(DP_pipe12[17]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_18_ ( .D(DP_pipe0_coeff_pipe02[18]), .CK(clk), 
        .RN(n1118), .Q(DP_pipe12[18]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_19_ ( .D(DP_pipe0_coeff_pipe02[19]), .CK(clk), 
        .RN(n1118), .Q(DP_pipe12[19]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_20_ ( .D(DP_pipe0_coeff_pipe02[20]), .CK(clk), 
        .RN(n1118), .Q(DP_pipe12[20]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_21_ ( .D(DP_pipe0_coeff_pipe02[21]), .CK(clk), 
        .RN(n1118), .Q(DP_pipe12[21]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_22_ ( .D(DP_pipe0_coeff_pipe02[22]), .CK(clk), 
        .RN(n1118), .Q(DP_pipe12[22]) );
  DFFR_X1 DP_reg_pipe12_Q_reg_23_ ( .D(DP_pipe0_coeff_pipe02[23]), .CK(clk), 
        .RN(n1118), .Q(DP_pipe12[23]) );
  DFFR_X1 DP_reg_pipe01_Q_reg_23_ ( .D(DP_sw0_23_), .CK(clk), .RN(n1118), .Q(
        DP_pipe01[23]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_0_ ( .D(DP_pipe0_coeff_pipe01[0]), .CK(clk), 
        .RN(n1119), .Q(DP_pipe11[0]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_1_ ( .D(DP_pipe0_coeff_pipe01[1]), .CK(clk), 
        .RN(n1119), .Q(DP_pipe11[1]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_2_ ( .D(DP_pipe0_coeff_pipe01[2]), .CK(clk), 
        .RN(n1119), .Q(DP_pipe11[2]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_3_ ( .D(DP_pipe0_coeff_pipe01[3]), .CK(clk), 
        .RN(n1119), .Q(DP_pipe11[3]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_4_ ( .D(DP_pipe0_coeff_pipe01[4]), .CK(clk), 
        .RN(n1119), .Q(DP_pipe11[4]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_5_ ( .D(DP_pipe0_coeff_pipe01[5]), .CK(clk), 
        .RN(n1119), .Q(DP_pipe11[5]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_6_ ( .D(DP_pipe0_coeff_pipe01[6]), .CK(clk), 
        .RN(n1119), .Q(DP_pipe11[6]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_7_ ( .D(DP_pipe0_coeff_pipe01[7]), .CK(clk), 
        .RN(n1119), .Q(DP_pipe11[7]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_8_ ( .D(DP_pipe0_coeff_pipe01[8]), .CK(clk), 
        .RN(n1119), .Q(DP_pipe11[8]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_9_ ( .D(DP_pipe0_coeff_pipe01[9]), .CK(clk), 
        .RN(n1119), .Q(DP_pipe11[9]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_10_ ( .D(DP_pipe0_coeff_pipe01[10]), .CK(clk), 
        .RN(n1119), .Q(DP_pipe11[10]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_11_ ( .D(DP_pipe0_coeff_pipe01[11]), .CK(clk), 
        .RN(n1119), .Q(DP_pipe11[11]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_12_ ( .D(DP_pipe0_coeff_pipe01[12]), .CK(clk), 
        .RN(n1120), .Q(DP_pipe11[12]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_13_ ( .D(DP_pipe0_coeff_pipe01[13]), .CK(clk), 
        .RN(n1120), .Q(DP_pipe11[13]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_14_ ( .D(DP_pipe0_coeff_pipe01[14]), .CK(clk), 
        .RN(n1120), .Q(DP_pipe11[14]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_15_ ( .D(DP_pipe0_coeff_pipe01[15]), .CK(clk), 
        .RN(n1120), .Q(DP_pipe11[15]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_16_ ( .D(DP_pipe0_coeff_pipe01[16]), .CK(clk), 
        .RN(n1120), .Q(DP_pipe11[16]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_17_ ( .D(DP_pipe0_coeff_pipe01[17]), .CK(clk), 
        .RN(n1120), .Q(DP_pipe11[17]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_18_ ( .D(DP_pipe0_coeff_pipe01[18]), .CK(clk), 
        .RN(n1120), .Q(DP_pipe11[18]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_19_ ( .D(DP_pipe0_coeff_pipe01[19]), .CK(clk), 
        .RN(n1120), .Q(DP_pipe11[19]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_20_ ( .D(DP_pipe0_coeff_pipe01[20]), .CK(clk), 
        .RN(n1120), .Q(DP_pipe11[20]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_21_ ( .D(DP_pipe0_coeff_pipe01[21]), .CK(clk), 
        .RN(n1120), .Q(DP_pipe11[21]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_22_ ( .D(DP_pipe0_coeff_pipe01[22]), .CK(clk), 
        .RN(n1120), .Q(DP_pipe11[22]) );
  DFFR_X1 DP_reg_pipe11_Q_reg_23_ ( .D(DP_pipe0_coeff_pipe01[23]), .CK(clk), 
        .RN(n1120), .Q(DP_pipe11[23]) );
  DFFR_X1 DP_reg_ret0_Q_reg_0_ ( .D(DP_sw0_coeff_ret0[0]), .CK(clk), .RN(n1121), .Q(DP_ret0[0]) );
  DFFR_X1 DP_reg_ret0_Q_reg_1_ ( .D(DP_sw0_coeff_ret0[1]), .CK(clk), .RN(n1121), .Q(DP_ret0[1]) );
  DFFR_X1 DP_reg_ret0_Q_reg_2_ ( .D(DP_sw0_coeff_ret0[2]), .CK(clk), .RN(n1121), .Q(DP_ret0[2]) );
  DFFR_X1 DP_reg_ret0_Q_reg_3_ ( .D(DP_sw0_coeff_ret0[3]), .CK(clk), .RN(n1121), .Q(DP_ret0[3]) );
  DFFR_X1 DP_reg_ret0_Q_reg_4_ ( .D(DP_sw0_coeff_ret0[4]), .CK(clk), .RN(n1121), .Q(DP_ret0[4]) );
  DFFR_X1 DP_reg_ret0_Q_reg_5_ ( .D(DP_sw0_coeff_ret0[5]), .CK(clk), .RN(n1121), .Q(DP_ret0[5]) );
  DFFR_X1 DP_reg_ret0_Q_reg_6_ ( .D(DP_sw0_coeff_ret0[6]), .CK(clk), .RN(n1121), .Q(DP_ret0[6]) );
  DFFR_X1 DP_reg_ret0_Q_reg_7_ ( .D(DP_sw0_coeff_ret0[7]), .CK(clk), .RN(n1121), .Q(DP_ret0[7]) );
  DFFR_X1 DP_reg_ret0_Q_reg_8_ ( .D(DP_sw0_coeff_ret0[8]), .CK(clk), .RN(n1121), .Q(DP_ret0[8]) );
  DFFR_X1 DP_reg_ret0_Q_reg_9_ ( .D(DP_sw0_coeff_ret0[9]), .CK(clk), .RN(n1121), .Q(DP_ret0[9]) );
  DFFR_X1 DP_reg_ret0_Q_reg_10_ ( .D(DP_sw0_coeff_ret0[10]), .CK(clk), .RN(
        n1121), .Q(DP_ret0[10]) );
  DFFR_X1 DP_reg_ret0_Q_reg_11_ ( .D(DP_sw0_coeff_ret0[11]), .CK(clk), .RN(
        n1121), .Q(DP_ret0[11]) );
  DFFR_X1 DP_reg_ret0_Q_reg_12_ ( .D(DP_sw0_coeff_ret0[12]), .CK(clk), .RN(
        n1122), .Q(DP_ret0[12]) );
  DFFR_X1 DP_reg_ret0_Q_reg_13_ ( .D(DP_sw0_coeff_ret0[13]), .CK(clk), .RN(
        n1122), .Q(DP_ret0[13]) );
  DFFR_X1 DP_reg_ret0_Q_reg_14_ ( .D(DP_sw0_coeff_ret0[14]), .CK(clk), .RN(
        n1122), .Q(DP_ret0[14]) );
  DFFR_X1 DP_reg_ret0_Q_reg_15_ ( .D(DP_sw0_coeff_ret0[15]), .CK(clk), .RN(
        n1122), .Q(DP_ret0[15]) );
  DFFR_X1 DP_reg_ret0_Q_reg_16_ ( .D(DP_sw0_coeff_ret0[16]), .CK(clk), .RN(
        n1122), .Q(DP_ret0[16]) );
  DFFR_X1 DP_reg_ret0_Q_reg_17_ ( .D(DP_sw0_coeff_ret0[17]), .CK(clk), .RN(
        n1122), .Q(DP_ret0[17]) );
  DFFR_X1 DP_reg_ret0_Q_reg_18_ ( .D(DP_sw0_coeff_ret0[18]), .CK(clk), .RN(
        n1122), .Q(DP_ret0[18]) );
  DFFR_X1 DP_reg_ret0_Q_reg_19_ ( .D(DP_sw0_coeff_ret0[19]), .CK(clk), .RN(
        n1122), .Q(DP_ret0[19]) );
  DFFR_X1 DP_reg_ret0_Q_reg_20_ ( .D(DP_sw0_coeff_ret0[20]), .CK(clk), .RN(
        n1122), .Q(DP_ret0[20]) );
  DFFR_X1 DP_reg_ret0_Q_reg_21_ ( .D(DP_sw0_coeff_ret0[21]), .CK(clk), .RN(
        n1122), .Q(DP_ret0[21]) );
  DFFR_X1 DP_reg_ret0_Q_reg_22_ ( .D(DP_sw0_coeff_ret0[22]), .CK(clk), .RN(
        n1122), .Q(DP_ret0[22]) );
  DFFR_X1 DP_reg_ret0_Q_reg_23_ ( .D(DP_sw0_coeff_ret0[23]), .CK(clk), .RN(
        n1122), .Q(DP_ret0[23]) );
  DFFR_X1 DP_reg_pipe00_Q_reg_23_ ( .D(DP_w_23_), .CK(clk), .RN(n1123), .Q(
        DP_pipe00[23]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_0_ ( .D(DP_pipe0_coeff_pipe00[0]), .CK(clk), 
        .RN(n1123), .Q(DP_pipe10[0]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_1_ ( .D(DP_pipe0_coeff_pipe00[1]), .CK(clk), 
        .RN(n1123), .Q(DP_pipe10[1]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_2_ ( .D(DP_pipe0_coeff_pipe00[2]), .CK(clk), 
        .RN(n1123), .Q(DP_pipe10[2]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_3_ ( .D(DP_pipe0_coeff_pipe00[3]), .CK(clk), 
        .RN(n1123), .Q(DP_pipe10[3]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_4_ ( .D(DP_pipe0_coeff_pipe00[4]), .CK(clk), 
        .RN(n1123), .Q(DP_pipe10[4]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_5_ ( .D(DP_pipe0_coeff_pipe00[5]), .CK(clk), 
        .RN(n1123), .Q(DP_pipe10[5]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_6_ ( .D(DP_pipe0_coeff_pipe00[6]), .CK(clk), 
        .RN(n1123), .Q(DP_pipe10[6]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_7_ ( .D(DP_pipe0_coeff_pipe00[7]), .CK(clk), 
        .RN(n1123), .Q(DP_pipe10[7]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_8_ ( .D(DP_pipe0_coeff_pipe00[8]), .CK(clk), 
        .RN(n1123), .Q(DP_pipe10[8]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_9_ ( .D(DP_pipe0_coeff_pipe00[9]), .CK(clk), 
        .RN(n1123), .Q(DP_pipe10[9]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_10_ ( .D(DP_pipe0_coeff_pipe00[10]), .CK(clk), 
        .RN(n1123), .Q(DP_pipe10[10]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_11_ ( .D(DP_pipe0_coeff_pipe00[11]), .CK(clk), 
        .RN(n1124), .Q(DP_pipe10[11]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_12_ ( .D(DP_pipe0_coeff_pipe00[12]), .CK(clk), 
        .RN(n1124), .Q(DP_pipe10[12]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_13_ ( .D(DP_pipe0_coeff_pipe00[13]), .CK(clk), 
        .RN(n1124), .Q(DP_pipe10[13]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_14_ ( .D(DP_pipe0_coeff_pipe00[14]), .CK(clk), 
        .RN(n1124), .Q(DP_pipe10[14]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_15_ ( .D(DP_pipe0_coeff_pipe00[15]), .CK(clk), 
        .RN(n1124), .Q(DP_pipe10[15]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_16_ ( .D(DP_pipe0_coeff_pipe00[16]), .CK(clk), 
        .RN(n1124), .Q(DP_pipe10[16]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_17_ ( .D(DP_pipe0_coeff_pipe00[17]), .CK(clk), 
        .RN(n1124), .Q(DP_pipe10[17]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_18_ ( .D(DP_pipe0_coeff_pipe00[18]), .CK(clk), 
        .RN(n1124), .Q(DP_pipe10[18]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_19_ ( .D(DP_pipe0_coeff_pipe00[19]), .CK(clk), 
        .RN(n1124), .Q(DP_pipe10[19]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_20_ ( .D(DP_pipe0_coeff_pipe00[20]), .CK(clk), 
        .RN(n1124), .Q(DP_pipe10[20]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_21_ ( .D(DP_pipe0_coeff_pipe00[21]), .CK(clk), 
        .RN(n1124), .Q(DP_pipe10[21]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_22_ ( .D(DP_pipe0_coeff_pipe00[22]), .CK(clk), 
        .RN(n1124), .Q(DP_pipe10[22]) );
  DFFR_X1 DP_reg_pipe10_Q_reg_23_ ( .D(DP_pipe0_coeff_pipe00[23]), .CK(clk), 
        .RN(n1125), .Q(DP_pipe10[23]) );
  DFFR_X1 DP_reg_sw2_Q_reg_23_ ( .D(n606), .CK(clk), .RN(n1125), .Q(DP_sw2[23]), .QN(n339) );
  DFFR_X1 DP_reg_pipe03_Q_reg_23_ ( .D(DP_sw2[23]), .CK(clk), .RN(n1125), .Q(
        DP_pipe03[23]) );
  DFFR_X1 DP_reg_sw2_Q_reg_22_ ( .D(n604), .CK(clk), .RN(n1125), .Q(DP_sw2[22]), .QN(n338) );
  DFFR_X1 DP_reg_pipe03_Q_reg_22_ ( .D(DP_sw2[22]), .CK(clk), .RN(n1125), .Q(
        DP_pipe03[22]) );
  DFFR_X1 DP_reg_sw2_Q_reg_21_ ( .D(n602), .CK(clk), .RN(n1125), .Q(DP_sw2[21]), .QN(n337) );
  DFFR_X1 DP_reg_pipe03_Q_reg_21_ ( .D(DP_sw2[21]), .CK(clk), .RN(n1125), .Q(
        DP_pipe03[21]) );
  DFFR_X1 DP_reg_sw2_Q_reg_20_ ( .D(n600), .CK(clk), .RN(n1125), .Q(DP_sw2[20]), .QN(n336) );
  DFFR_X1 DP_reg_pipe03_Q_reg_20_ ( .D(DP_sw2[20]), .CK(clk), .RN(n1125), .Q(
        DP_pipe03[20]) );
  DFFR_X1 DP_reg_sw2_Q_reg_19_ ( .D(n598), .CK(clk), .RN(n1125), .Q(DP_sw2[19]), .QN(n335) );
  DFFR_X1 DP_reg_pipe03_Q_reg_19_ ( .D(DP_sw2[19]), .CK(clk), .RN(n1125), .Q(
        DP_pipe03[19]) );
  DFFR_X1 DP_reg_sw2_Q_reg_18_ ( .D(n596), .CK(clk), .RN(n1125), .Q(DP_sw2[18]), .QN(n334) );
  DFFR_X1 DP_reg_pipe03_Q_reg_18_ ( .D(DP_sw2[18]), .CK(clk), .RN(n1126), .Q(
        DP_pipe03[18]) );
  DFFR_X1 DP_reg_sw2_Q_reg_17_ ( .D(n594), .CK(clk), .RN(n1126), .Q(DP_sw2[17]), .QN(n333) );
  DFFR_X1 DP_reg_pipe03_Q_reg_17_ ( .D(DP_sw2[17]), .CK(clk), .RN(n1126), .Q(
        DP_pipe03[17]) );
  DFFR_X1 DP_reg_sw2_Q_reg_16_ ( .D(n592), .CK(clk), .RN(n1126), .Q(DP_sw2[16]), .QN(n332) );
  DFFR_X1 DP_reg_pipe03_Q_reg_16_ ( .D(DP_sw2[16]), .CK(clk), .RN(n1126), .Q(
        DP_pipe03[16]) );
  DFFR_X1 DP_reg_sw2_Q_reg_15_ ( .D(n590), .CK(clk), .RN(n1126), .Q(DP_sw2[15]), .QN(n331) );
  DFFR_X1 DP_reg_pipe03_Q_reg_15_ ( .D(DP_sw2[15]), .CK(clk), .RN(n1126), .Q(
        DP_pipe03[15]) );
  DFFR_X1 DP_reg_sw2_Q_reg_14_ ( .D(n588), .CK(clk), .RN(n1126), .Q(DP_sw2[14]), .QN(n330) );
  DFFR_X1 DP_reg_pipe03_Q_reg_14_ ( .D(DP_sw2[14]), .CK(clk), .RN(n1126), .Q(
        DP_pipe03[14]) );
  DFFR_X1 DP_reg_sw2_Q_reg_13_ ( .D(n586), .CK(clk), .RN(n1126), .Q(DP_sw2[13]), .QN(n329) );
  DFFR_X1 DP_reg_pipe03_Q_reg_13_ ( .D(DP_sw2[13]), .CK(clk), .RN(n1126), .Q(
        DP_pipe03[13]) );
  DFFR_X1 DP_reg_sw2_Q_reg_12_ ( .D(n584), .CK(clk), .RN(n1126), .Q(DP_sw2[12]), .QN(n328) );
  DFFR_X1 DP_reg_pipe03_Q_reg_12_ ( .D(DP_sw2[12]), .CK(clk), .RN(n1127), .Q(
        DP_pipe03[12]) );
  DFFR_X1 DP_reg_sw2_Q_reg_11_ ( .D(n582), .CK(clk), .RN(n1127), .Q(DP_sw2[11]), .QN(n327) );
  DFFR_X1 DP_reg_pipe03_Q_reg_11_ ( .D(DP_sw2[11]), .CK(clk), .RN(n1127), .Q(
        DP_pipe03[11]) );
  DFFR_X1 DP_reg_sw2_Q_reg_10_ ( .D(n580), .CK(clk), .RN(n1127), .Q(DP_sw2[10]), .QN(n326) );
  DFFR_X1 DP_reg_pipe03_Q_reg_10_ ( .D(DP_sw2[10]), .CK(clk), .RN(n1127), .Q(
        DP_pipe03[10]) );
  DFFR_X1 DP_reg_sw2_Q_reg_9_ ( .D(n578), .CK(clk), .RN(n1127), .Q(DP_sw2[9]), 
        .QN(n325) );
  DFFR_X1 DP_reg_pipe03_Q_reg_9_ ( .D(DP_sw2[9]), .CK(clk), .RN(n1127), .Q(
        DP_pipe03[9]) );
  DFFR_X1 DP_reg_sw2_Q_reg_8_ ( .D(n576), .CK(clk), .RN(n1127), .Q(DP_sw2[8]), 
        .QN(n324) );
  DFFR_X1 DP_reg_pipe03_Q_reg_8_ ( .D(DP_sw2[8]), .CK(clk), .RN(n1127), .Q(
        DP_pipe03[8]) );
  DFFR_X1 DP_reg_sw2_Q_reg_7_ ( .D(n574), .CK(clk), .RN(n1127), .Q(DP_sw2[7]), 
        .QN(n323) );
  DFFR_X1 DP_reg_pipe03_Q_reg_7_ ( .D(DP_sw2[7]), .CK(clk), .RN(n1127), .Q(
        DP_pipe03[7]) );
  DFFR_X1 DP_reg_sw2_Q_reg_6_ ( .D(n572), .CK(clk), .RN(n1127), .Q(DP_sw2[6]), 
        .QN(n322) );
  DFFR_X1 DP_reg_pipe03_Q_reg_6_ ( .D(DP_sw2[6]), .CK(clk), .RN(n1128), .Q(
        DP_pipe03[6]) );
  DFFR_X1 DP_reg_sw2_Q_reg_5_ ( .D(n570), .CK(clk), .RN(n1128), .Q(DP_sw2[5]), 
        .QN(n321) );
  DFFR_X1 DP_reg_pipe03_Q_reg_5_ ( .D(DP_sw2[5]), .CK(clk), .RN(n1128), .Q(
        DP_pipe03[5]) );
  DFFR_X1 DP_reg_sw2_Q_reg_4_ ( .D(n568), .CK(clk), .RN(n1128), .Q(DP_sw2[4]), 
        .QN(n320) );
  DFFR_X1 DP_reg_pipe03_Q_reg_4_ ( .D(DP_sw2[4]), .CK(clk), .RN(n1128), .Q(
        DP_pipe03[4]) );
  DFFR_X1 DP_reg_sw2_Q_reg_3_ ( .D(n566), .CK(clk), .RN(n1128), .Q(DP_sw2[3]), 
        .QN(n319) );
  DFFR_X1 DP_reg_pipe03_Q_reg_3_ ( .D(DP_sw2[3]), .CK(clk), .RN(n1128), .Q(
        DP_pipe03[3]) );
  DFFR_X1 DP_reg_sw2_Q_reg_2_ ( .D(n564), .CK(clk), .RN(n1128), .Q(DP_sw2[2]), 
        .QN(n318) );
  DFFR_X1 DP_reg_pipe03_Q_reg_2_ ( .D(DP_sw2[2]), .CK(clk), .RN(n1128), .Q(
        DP_pipe03[2]) );
  DFFR_X1 DP_reg_sw2_Q_reg_1_ ( .D(n562), .CK(clk), .RN(n1128), .Q(DP_sw2[1]), 
        .QN(n317) );
  DFFR_X1 DP_reg_pipe03_Q_reg_1_ ( .D(DP_sw2[1]), .CK(clk), .RN(n1128), .Q(
        DP_pipe03[1]) );
  DFFR_X1 DP_reg_sw2_Q_reg_0_ ( .D(n560), .CK(clk), .RN(n1128), .Q(DP_sw2[0]), 
        .QN(n316) );
  DFFR_X1 DP_reg_pipe03_Q_reg_0_ ( .D(DP_sw2[0]), .CK(clk), .RN(n1129), .Q(
        DP_pipe03[0]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_0_ ( .D(DP_pipe0_coeff_pipe03[0]), .CK(clk), 
        .RN(n1129), .Q(DP_pipe13[0]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_1_ ( .D(DP_pipe0_coeff_pipe03[1]), .CK(clk), 
        .RN(n1129), .Q(DP_pipe13[1]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_2_ ( .D(DP_pipe0_coeff_pipe03[2]), .CK(clk), 
        .RN(n1129), .Q(DP_pipe13[2]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_3_ ( .D(DP_pipe0_coeff_pipe03[3]), .CK(clk), 
        .RN(n1129), .Q(DP_pipe13[3]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_4_ ( .D(DP_pipe0_coeff_pipe03[4]), .CK(clk), 
        .RN(n1129), .Q(DP_pipe13[4]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_5_ ( .D(DP_pipe0_coeff_pipe03[5]), .CK(clk), 
        .RN(n1129), .Q(DP_pipe13[5]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_6_ ( .D(DP_pipe0_coeff_pipe03[6]), .CK(clk), 
        .RN(n1129), .Q(DP_pipe13[6]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_7_ ( .D(DP_pipe0_coeff_pipe03[7]), .CK(clk), 
        .RN(n1129), .Q(DP_pipe13[7]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_8_ ( .D(DP_pipe0_coeff_pipe03[8]), .CK(clk), 
        .RN(n1129), .Q(DP_pipe13[8]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_9_ ( .D(DP_pipe0_coeff_pipe03[9]), .CK(clk), 
        .RN(n1129), .Q(DP_pipe13[9]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_10_ ( .D(DP_pipe0_coeff_pipe03[10]), .CK(clk), 
        .RN(n1129), .Q(DP_pipe13[10]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_11_ ( .D(DP_pipe0_coeff_pipe03[11]), .CK(clk), 
        .RN(n1130), .Q(DP_pipe13[11]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_12_ ( .D(DP_pipe0_coeff_pipe03[12]), .CK(clk), 
        .RN(n1130), .Q(DP_pipe13[12]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_13_ ( .D(DP_pipe0_coeff_pipe03[13]), .CK(clk), 
        .RN(n1130), .Q(DP_pipe13[13]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_14_ ( .D(DP_pipe0_coeff_pipe03[14]), .CK(clk), 
        .RN(n1130), .Q(DP_pipe13[14]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_15_ ( .D(DP_pipe0_coeff_pipe03[15]), .CK(clk), 
        .RN(n1130), .Q(DP_pipe13[15]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_16_ ( .D(DP_pipe0_coeff_pipe03[16]), .CK(clk), 
        .RN(n1130), .Q(DP_pipe13[16]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_17_ ( .D(DP_pipe0_coeff_pipe03[17]), .CK(clk), 
        .RN(n1130), .Q(DP_pipe13[17]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_18_ ( .D(DP_pipe0_coeff_pipe03[18]), .CK(clk), 
        .RN(n1130), .Q(DP_pipe13[18]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_19_ ( .D(DP_pipe0_coeff_pipe03[19]), .CK(clk), 
        .RN(n1130), .Q(DP_pipe13[19]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_20_ ( .D(DP_pipe0_coeff_pipe03[20]), .CK(clk), 
        .RN(n1130), .Q(DP_pipe13[20]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_21_ ( .D(DP_pipe0_coeff_pipe03[21]), .CK(clk), 
        .RN(n1130), .Q(DP_pipe13[21]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_22_ ( .D(DP_pipe0_coeff_pipe03[22]), .CK(clk), 
        .RN(n1130), .Q(DP_pipe13[22]) );
  DFFR_X1 DP_reg_pipe13_Q_reg_23_ ( .D(DP_pipe0_coeff_pipe03[23]), .CK(clk), 
        .RN(n1131), .Q(DP_pipe13[23]) );
  DFFR_X1 CU_presentState_reg_0_ ( .D(CU_nextState_0_), .CK(clk), .RN(n1131), 
        .QN(n315) );
  DFFR_X1 reg_delay_0_Q_reg_0_ ( .D(delayed_controls_0__1_), .CK(clk), .RN(
        n1131), .Q(delayed_controls_1__1_) );
  DFFR_X1 reg_delay_0_Q_reg_1_ ( .D(n1033), .CK(clk), .RN(n1131), .Q(
        delayed_controls_1__0_) );
  DFFR_X1 reg_delay_1_Q_reg_0_ ( .D(delayed_controls_1__1_), .CK(clk), .RN(
        n1131), .Q(vOut) );
  DFFR_X1 reg_delay_1_Q_reg_1_ ( .D(delayed_controls_1__0_), .CK(clk), .RN(
        n1131), .Q(delayed_controls_2__0_), .QN(n1027) );
  DFFR_X1 DP_reg_out_Q_reg_11_ ( .D(n531), .CK(clk), .RN(n1131), .Q(dOut[11]), 
        .QN(n313) );
  DFFR_X1 DP_reg_out_Q_reg_10_ ( .D(n530), .CK(clk), .RN(n1131), .Q(dOut[10]), 
        .QN(n312) );
  DFFR_X1 DP_reg_out_Q_reg_9_ ( .D(n529), .CK(clk), .RN(n1131), .Q(dOut[9]), 
        .QN(n311) );
  DFFR_X1 DP_reg_out_Q_reg_8_ ( .D(n528), .CK(clk), .RN(n1131), .Q(dOut[8]), 
        .QN(n310) );
  DFFR_X1 DP_reg_out_Q_reg_7_ ( .D(n527), .CK(clk), .RN(n1131), .Q(dOut[7]), 
        .QN(n309) );
  DFFR_X1 DP_reg_out_Q_reg_6_ ( .D(n526), .CK(clk), .RN(n1131), .Q(dOut[6]), 
        .QN(n308) );
  DFFR_X1 DP_reg_out_Q_reg_5_ ( .D(n525), .CK(clk), .RN(n1132), .Q(dOut[5]), 
        .QN(n307) );
  DFFR_X1 DP_reg_out_Q_reg_4_ ( .D(n524), .CK(clk), .RN(n1132), .Q(dOut[4]), 
        .QN(n306) );
  DFFR_X1 DP_reg_out_Q_reg_3_ ( .D(n523), .CK(clk), .RN(n1132), .Q(dOut[3]), 
        .QN(n305) );
  DFFR_X1 DP_reg_out_Q_reg_2_ ( .D(n522), .CK(clk), .RN(n1132), .Q(dOut[2]), 
        .QN(n304) );
  DFFR_X1 DP_reg_out_Q_reg_1_ ( .D(n521), .CK(clk), .RN(n1132), .Q(dOut[1]), 
        .QN(n303) );
  DFFR_X1 DP_reg_out_Q_reg_0_ ( .D(n520), .CK(clk), .RN(n1132), .Q(dOut[0]), 
        .QN(n302) );
  XOR2_X1 U501 ( .A(n1086), .B(n1033), .Z(CU_nextState_0_) );
  XOR2_X1 U503 ( .A(n315), .B(delayed_controls_0__1_), .Z(n74) );
  iir_filter_DW01_add_0 DP_add_223 ( .A({DP_pipe10[23], DP_pipe10[22], 
        DP_pipe10[21], DP_pipe10[20], DP_pipe10[19], DP_pipe10[18], 
        DP_pipe10[17], DP_pipe10[16], DP_pipe10[15], DP_pipe10[14], 
        DP_pipe10[13], DP_pipe10[12], DP_pipe10[11], DP_pipe10[10], 
        DP_pipe10[9], DP_pipe10[8], DP_pipe10[7], DP_pipe10[6], DP_pipe10[5], 
        DP_pipe10[4], DP_pipe10[3], DP_pipe10[2], DP_pipe10[1], DP_pipe10[0]}), 
        .B({DP_ff[23], DP_ff[22], DP_ff[21], DP_ff[20], DP_ff[19], DP_ff[18], 
        DP_ff[17], DP_ff[16], DP_ff[15], DP_ff[14], DP_ff[13], DP_ff[12], 
        DP_ff[11], DP_ff[10], DP_ff[9], DP_ff[8], DP_ff[7], DP_ff[6], DP_ff[5], 
        DP_ff[4], DP_ff[3], DP_ff[2], DP_ff[1], DP_ff[0]}), .CI(1'b0), .SUM({
        DP_y_23, DP_y_11_, DP_y_10_, DP_y_9_, DP_y_8_, DP_y_7_, DP_y_6_, 
        DP_y_5_, DP_y_4_, DP_y_3_, DP_y_2_, DP_y_1_, DP_y_0_, 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10}) );
  iir_filter_DW01_sub_0 DP_sub_217 ( .A({DP_x[11], DP_x[11], DP_x[10], DP_x[9], 
        DP_x[8], DP_x[7], DP_x[6], DP_x[5], DP_x[4], DP_x[3], DP_x[2], DP_x[1], 
        DP_x[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({DP_fb[23], DP_fb[22], DP_fb[21], DP_fb[20], DP_fb[19], 
        DP_fb[18], DP_fb[17], DP_fb[16], DP_fb[15], DP_fb[14], DP_fb[13], 
        DP_fb[12], DP_fb[11], DP_fb[10], DP_fb[9], DP_fb[8], DP_fb[7], 
        DP_fb[6], DP_fb[5], DP_fb[4], DP_fb[3], DP_fb[2], DP_fb[1], DP_fb[0]}), 
        .CI(1'b0), .DIFF({DP_w_23_, DP_w_22_, DP_w_21_, DP_w_20_, DP_w_19_, 
        DP_w_18_, DP_w_17_, DP_w_16_, DP_w_15_, DP_w_14_, DP_w_13_, DP_w_12_, 
        DP_w_11_, DP_w_10_, DP_w_9_, DP_w_8_, DP_w_7_, DP_w_6_, DP_w_5_, 
        DP_w_4_, DP_w_3_, DP_w_2_, DP_w_1_, DP_w_0_}) );
  iir_filter_DW01_add_1 DP_add_216 ( .A({DP_pipe11[23], DP_pipe11[22], 
        DP_pipe11[21], DP_pipe11[20], DP_pipe11[19], DP_pipe11[18], 
        DP_pipe11[17], DP_pipe11[16], DP_pipe11[15], DP_pipe11[14], 
        DP_pipe11[13], DP_pipe11[12], DP_pipe11[11], DP_pipe11[10], 
        DP_pipe11[9], DP_pipe11[8], DP_pipe11[7], DP_pipe11[6], DP_pipe11[5], 
        DP_pipe11[4], DP_pipe11[3], DP_pipe11[2], DP_pipe11[1], DP_pipe11[0]}), 
        .B({DP_ff_part[23], DP_ff_part[22], DP_ff_part[21], DP_ff_part[20], 
        DP_ff_part[19], DP_ff_part[18], DP_ff_part[17], DP_ff_part[16], 
        DP_ff_part[15], DP_ff_part[14], DP_ff_part[13], DP_ff_part[12], 
        DP_ff_part[11], DP_ff_part[10], DP_ff_part[9], DP_ff_part[8], 
        DP_ff_part[7], DP_ff_part[6], DP_ff_part[5], DP_ff_part[4], 
        DP_ff_part[3], DP_ff_part[2], DP_ff_part[1], DP_ff_part[0]}), .CI(1'b0), .SUM({DP_ff[23], DP_ff[22], DP_ff[21], DP_ff[20], DP_ff[19], DP_ff[18], 
        DP_ff[17], DP_ff[16], DP_ff[15], DP_ff[14], DP_ff[13], DP_ff[12], 
        DP_ff[11], DP_ff[10], DP_ff[9], DP_ff[8], DP_ff[7], DP_ff[6], DP_ff[5], 
        DP_ff[4], DP_ff[3], DP_ff[2], DP_ff[1], DP_ff[0]}) );
  iir_filter_DW01_add_2 DP_add_215 ( .A({DP_pipe12[23], DP_pipe12[22], 
        DP_pipe12[21], DP_pipe12[20], DP_pipe12[19], DP_pipe12[18], 
        DP_pipe12[17], DP_pipe12[16], DP_pipe12[15], DP_pipe12[14], 
        DP_pipe12[13], DP_pipe12[12], DP_pipe12[11], DP_pipe12[10], 
        DP_pipe12[9], DP_pipe12[8], DP_pipe12[7], DP_pipe12[6], DP_pipe12[5], 
        DP_pipe12[4], DP_pipe12[3], DP_pipe12[2], DP_pipe12[1], DP_pipe12[0]}), 
        .B({DP_pipe13[23], DP_pipe13[22], DP_pipe13[21], DP_pipe13[20], 
        DP_pipe13[19], DP_pipe13[18], DP_pipe13[17], DP_pipe13[16], 
        DP_pipe13[15], DP_pipe13[14], DP_pipe13[13], DP_pipe13[12], 
        DP_pipe13[11], DP_pipe13[10], DP_pipe13[9], DP_pipe13[8], DP_pipe13[7], 
        DP_pipe13[6], DP_pipe13[5], DP_pipe13[4], DP_pipe13[3], DP_pipe13[2], 
        DP_pipe13[1], DP_pipe13[0]}), .CI(1'b0), .SUM({DP_ff_part[23], 
        DP_ff_part[22], DP_ff_part[21], DP_ff_part[20], DP_ff_part[19], 
        DP_ff_part[18], DP_ff_part[17], DP_ff_part[16], DP_ff_part[15], 
        DP_ff_part[14], DP_ff_part[13], DP_ff_part[12], DP_ff_part[11], 
        DP_ff_part[10], DP_ff_part[9], DP_ff_part[8], DP_ff_part[7], 
        DP_ff_part[6], DP_ff_part[5], DP_ff_part[4], DP_ff_part[3], 
        DP_ff_part[2], DP_ff_part[1], DP_ff_part[0]}) );
  iir_filter_DW01_add_3 DP_add_214 ( .A({DP_ret0[23], DP_ret0[22], DP_ret0[21], 
        DP_ret0[20], DP_ret0[19], DP_ret0[18], DP_ret0[17], DP_ret0[16], 
        DP_ret0[15], DP_ret0[14], DP_ret0[13], DP_ret0[12], DP_ret0[11], 
        DP_ret0[10], DP_ret0[9], DP_ret0[8], DP_ret0[7], DP_ret0[6], 
        DP_ret0[5], DP_ret0[4], DP_ret0[3], DP_ret0[2], DP_ret0[1], DP_ret0[0]}), .B({DP_ret1[23], DP_ret1[22], DP_ret1[21], DP_ret1[20], DP_ret1[19], 
        DP_ret1[18], DP_ret1[17], DP_ret1[16], DP_ret1[15], DP_ret1[14], 
        DP_ret1[13], DP_ret1[12], DP_ret1[11], DP_ret1[10], DP_ret1[9], 
        DP_ret1[8], DP_ret1[7], DP_ret1[6], DP_ret1[5], DP_ret1[4], DP_ret1[3], 
        DP_ret1[2], DP_ret1[1], DP_ret1[0]}), .CI(1'b0), .SUM({DP_fb[23], 
        DP_fb[22], DP_fb[21], DP_fb[20], DP_fb[19], DP_fb[18], DP_fb[17], 
        DP_fb[16], DP_fb[15], DP_fb[14], DP_fb[13], DP_fb[12], DP_fb[11], 
        DP_fb[10], DP_fb[9], DP_fb[8], DP_fb[7], DP_fb[6], DP_fb[5], DP_fb[4], 
        DP_fb[3], DP_fb[2], DP_fb[1], DP_fb[0]}) );
  iir_filter_DW02_mult_0 DP_mult_209 ( .A({DP_coeffs_ff_int[72], 
        DP_coeffs_ff_int[73], DP_coeffs_ff_int[74], DP_coeffs_ff_int[75], 
        DP_coeffs_ff_int[76], DP_coeffs_ff_int[77], DP_coeffs_ff_int[78], 
        DP_coeffs_ff_int[79], DP_coeffs_ff_int[80], DP_coeffs_ff_int[81], 
        DP_coeffs_ff_int[82], DP_coeffs_ff_int[83], DP_coeffs_ff_int[84], 
        DP_coeffs_ff_int[85], DP_coeffs_ff_int[86], DP_coeffs_ff_int[87], 
        DP_coeffs_ff_int[88], DP_coeffs_ff_int[89], DP_coeffs_ff_int[90], 
        DP_coeffs_ff_int[91], DP_coeffs_ff_int[92], DP_coeffs_ff_int[93], 
        DP_coeffs_ff_int[94], DP_coeffs_ff_int[95]}), .B({DP_pipe03[23], 
        DP_pipe03[22], DP_pipe03[21], DP_pipe03[20], DP_pipe03[19], 
        DP_pipe03[18], DP_pipe03[17], DP_pipe03[16], DP_pipe03[15], 
        DP_pipe03[14], DP_pipe03[13], DP_pipe03[12], DP_pipe03[11], 
        DP_pipe03[10], DP_pipe03[9], DP_pipe03[8], DP_pipe03[7], DP_pipe03[6], 
        DP_pipe03[5], DP_pipe03[4], DP_pipe03[3], DP_pipe03[2], DP_pipe03[1], 
        DP_pipe03[0]}), .PRODUCT({DP_pipe0_coeff_pipe03[23], 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        DP_pipe0_coeff_pipe03[22], DP_pipe0_coeff_pipe03[21], 
        DP_pipe0_coeff_pipe03[20], DP_pipe0_coeff_pipe03[19], 
        DP_pipe0_coeff_pipe03[18], DP_pipe0_coeff_pipe03[17], 
        DP_pipe0_coeff_pipe03[16], DP_pipe0_coeff_pipe03[15], 
        DP_pipe0_coeff_pipe03[14], DP_pipe0_coeff_pipe03[13], 
        DP_pipe0_coeff_pipe03[12], DP_pipe0_coeff_pipe03[11], 
        DP_pipe0_coeff_pipe03[10], DP_pipe0_coeff_pipe03[9], 
        DP_pipe0_coeff_pipe03[8], DP_pipe0_coeff_pipe03[7], 
        DP_pipe0_coeff_pipe03[6], DP_pipe0_coeff_pipe03[5], 
        DP_pipe0_coeff_pipe03[4], DP_pipe0_coeff_pipe03[3], 
        DP_pipe0_coeff_pipe03[2], DP_pipe0_coeff_pipe03[1], 
        DP_pipe0_coeff_pipe03[0], SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34}), .TC(1'b1) );
  iir_filter_DW02_mult_1 DP_mult_208 ( .A({DP_coeffs_ff_int[48], 
        DP_coeffs_ff_int[49], DP_coeffs_ff_int[50], DP_coeffs_ff_int[51], 
        DP_coeffs_ff_int[52], DP_coeffs_ff_int[53], DP_coeffs_ff_int[54], 
        DP_coeffs_ff_int[55], DP_coeffs_ff_int[56], DP_coeffs_ff_int[57], 
        DP_coeffs_ff_int[58], DP_coeffs_ff_int[59], DP_coeffs_ff_int[60], 
        DP_coeffs_ff_int[61], DP_coeffs_ff_int[62], DP_coeffs_ff_int[63], 
        DP_coeffs_ff_int[64], DP_coeffs_ff_int[65], DP_coeffs_ff_int[66], 
        DP_coeffs_ff_int[67], DP_coeffs_ff_int[68], DP_coeffs_ff_int[69], 
        DP_coeffs_ff_int[70], DP_coeffs_ff_int[71]}), .B({DP_pipe02[23], 
        DP_pipe02[22], DP_pipe02[21], DP_pipe02[20], DP_pipe02[19], 
        DP_pipe02[18], DP_pipe02[17], DP_pipe02[16], DP_pipe02[15], 
        DP_pipe02[14], DP_pipe02[13], DP_pipe02[12], DP_pipe02[11], 
        DP_pipe02[10], DP_pipe02[9], DP_pipe02[8], DP_pipe02[7], DP_pipe02[6], 
        DP_pipe02[5], DP_pipe02[4], DP_pipe02[3], DP_pipe02[2], DP_pipe02[1], 
        DP_pipe02[0]}), .PRODUCT({DP_pipe0_coeff_pipe02[23], 
        SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, 
        DP_pipe0_coeff_pipe02[22], DP_pipe0_coeff_pipe02[21], 
        DP_pipe0_coeff_pipe02[20], DP_pipe0_coeff_pipe02[19], 
        DP_pipe0_coeff_pipe02[18], DP_pipe0_coeff_pipe02[17], 
        DP_pipe0_coeff_pipe02[16], DP_pipe0_coeff_pipe02[15], 
        DP_pipe0_coeff_pipe02[14], DP_pipe0_coeff_pipe02[13], 
        DP_pipe0_coeff_pipe02[12], DP_pipe0_coeff_pipe02[11], 
        DP_pipe0_coeff_pipe02[10], DP_pipe0_coeff_pipe02[9], 
        DP_pipe0_coeff_pipe02[8], DP_pipe0_coeff_pipe02[7], 
        DP_pipe0_coeff_pipe02[6], DP_pipe0_coeff_pipe02[5], 
        DP_pipe0_coeff_pipe02[4], DP_pipe0_coeff_pipe02[3], 
        DP_pipe0_coeff_pipe02[2], DP_pipe0_coeff_pipe02[1], 
        DP_pipe0_coeff_pipe02[0], SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58}), .TC(1'b1) );
  iir_filter_DW02_mult_2 DP_mult_207 ( .A({DP_coeffs_ff_int[24], 
        DP_coeffs_ff_int[25], DP_coeffs_ff_int[26], DP_coeffs_ff_int[27], 
        DP_coeffs_ff_int[28], DP_coeffs_ff_int[29], DP_coeffs_ff_int[30], 
        DP_coeffs_ff_int[31], DP_coeffs_ff_int[32], DP_coeffs_ff_int[33], 
        DP_coeffs_ff_int[34], DP_coeffs_ff_int[35], DP_coeffs_ff_int[36], 
        DP_coeffs_ff_int[37], DP_coeffs_ff_int[38], DP_coeffs_ff_int[39], 
        DP_coeffs_ff_int[40], DP_coeffs_ff_int[41], DP_coeffs_ff_int[42], 
        DP_coeffs_ff_int[43], DP_coeffs_ff_int[44], DP_coeffs_ff_int[45], 
        DP_coeffs_ff_int[46], DP_coeffs_ff_int[47]}), .B({DP_pipe01[23], 
        DP_pipe01[22], DP_pipe01[21], DP_pipe01[20], DP_pipe01[19], 
        DP_pipe01[18], DP_pipe01[17], DP_pipe01[16], DP_pipe01[15], 
        DP_pipe01[14], DP_pipe01[13], DP_pipe01[12], DP_pipe01[11], 
        DP_pipe01[10], DP_pipe01[9], DP_pipe01[8], DP_pipe01[7], DP_pipe01[6], 
        DP_pipe01[5], DP_pipe01[4], DP_pipe01[3], DP_pipe01[2], DP_pipe01[1], 
        DP_pipe01[0]}), .PRODUCT({DP_pipe0_coeff_pipe01[23], 
        SYNOPSYS_UNCONNECTED__59, SYNOPSYS_UNCONNECTED__60, 
        DP_pipe0_coeff_pipe01[22], DP_pipe0_coeff_pipe01[21], 
        DP_pipe0_coeff_pipe01[20], DP_pipe0_coeff_pipe01[19], 
        DP_pipe0_coeff_pipe01[18], DP_pipe0_coeff_pipe01[17], 
        DP_pipe0_coeff_pipe01[16], DP_pipe0_coeff_pipe01[15], 
        DP_pipe0_coeff_pipe01[14], DP_pipe0_coeff_pipe01[13], 
        DP_pipe0_coeff_pipe01[12], DP_pipe0_coeff_pipe01[11], 
        DP_pipe0_coeff_pipe01[10], DP_pipe0_coeff_pipe01[9], 
        DP_pipe0_coeff_pipe01[8], DP_pipe0_coeff_pipe01[7], 
        DP_pipe0_coeff_pipe01[6], DP_pipe0_coeff_pipe01[5], 
        DP_pipe0_coeff_pipe01[4], DP_pipe0_coeff_pipe01[3], 
        DP_pipe0_coeff_pipe01[2], DP_pipe0_coeff_pipe01[1], 
        DP_pipe0_coeff_pipe01[0], SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82}), .TC(1'b1) );
  iir_filter_DW02_mult_3 DP_mult_206 ( .A({DP_coeffs_ff_int[0], 
        DP_coeffs_ff_int[1], DP_coeffs_ff_int[2], DP_coeffs_ff_int[3], 
        DP_coeffs_ff_int[4], DP_coeffs_ff_int[5], DP_coeffs_ff_int[6], 
        DP_coeffs_ff_int[7], DP_coeffs_ff_int[8], DP_coeffs_ff_int[9], 
        DP_coeffs_ff_int[10], DP_coeffs_ff_int[11], DP_coeffs_ff_int[12], 
        DP_coeffs_ff_int[13], DP_coeffs_ff_int[14], DP_coeffs_ff_int[15], 
        DP_coeffs_ff_int[16], DP_coeffs_ff_int[17], DP_coeffs_ff_int[18], 
        DP_coeffs_ff_int[19], DP_coeffs_ff_int[20], DP_coeffs_ff_int[21], 
        DP_coeffs_ff_int[22], DP_coeffs_ff_int[23]}), .B({DP_pipe00[23], 
        DP_pipe00[22], DP_pipe00[21], DP_pipe00[20], DP_pipe00[19], 
        DP_pipe00[18], DP_pipe00[17], DP_pipe00[16], DP_pipe00[15], 
        DP_pipe00[14], DP_pipe00[13], DP_pipe00[12], DP_pipe00[11], 
        DP_pipe00[10], DP_pipe00[9], DP_pipe00[8], DP_pipe00[7], DP_pipe00[6], 
        DP_pipe00[5], DP_pipe00[4], DP_pipe00[3], DP_pipe00[2], DP_pipe00[1], 
        DP_pipe00[0]}), .PRODUCT({DP_pipe0_coeff_pipe00[23], 
        SYNOPSYS_UNCONNECTED__83, SYNOPSYS_UNCONNECTED__84, 
        DP_pipe0_coeff_pipe00[22], DP_pipe0_coeff_pipe00[21], 
        DP_pipe0_coeff_pipe00[20], DP_pipe0_coeff_pipe00[19], 
        DP_pipe0_coeff_pipe00[18], DP_pipe0_coeff_pipe00[17], 
        DP_pipe0_coeff_pipe00[16], DP_pipe0_coeff_pipe00[15], 
        DP_pipe0_coeff_pipe00[14], DP_pipe0_coeff_pipe00[13], 
        DP_pipe0_coeff_pipe00[12], DP_pipe0_coeff_pipe00[11], 
        DP_pipe0_coeff_pipe00[10], DP_pipe0_coeff_pipe00[9], 
        DP_pipe0_coeff_pipe00[8], DP_pipe0_coeff_pipe00[7], 
        DP_pipe0_coeff_pipe00[6], DP_pipe0_coeff_pipe00[5], 
        DP_pipe0_coeff_pipe00[4], DP_pipe0_coeff_pipe00[3], 
        DP_pipe0_coeff_pipe00[2], DP_pipe0_coeff_pipe00[1], 
        DP_pipe0_coeff_pipe00[0], SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106}), .TC(1'b1) );
  iir_filter_DW02_mult_4 DP_mult_205 ( .A({DP_coeffs_fb_int[24], 
        DP_coeffs_fb_int[25], DP_coeffs_fb_int[26], DP_coeffs_fb_int[27], 
        DP_coeffs_fb_int[28], DP_coeffs_fb_int[29], DP_coeffs_fb_int[30], 
        DP_coeffs_fb_int[31], DP_coeffs_fb_int[32], DP_coeffs_fb_int[33], 
        DP_coeffs_fb_int[34], DP_coeffs_fb_int[35], DP_coeffs_fb_int[36], 
        DP_coeffs_fb_int[37], DP_coeffs_fb_int[38], DP_coeffs_fb_int[39], 
        DP_coeffs_fb_int[40], DP_coeffs_fb_int[41], DP_coeffs_fb_int[42], 
        DP_coeffs_fb_int[43], DP_coeffs_fb_int[44], DP_coeffs_fb_int[45], 
        DP_coeffs_fb_int[46], DP_coeffs_fb_int[47]}), .B({n1058, DP_sw1_22_, 
        DP_sw1_21_, DP_sw1_20_, DP_sw1_19_, DP_sw1_18_, DP_sw1_17_, DP_sw1_16_, 
        DP_sw1_15_, DP_sw1_14_, DP_sw1_13_, DP_sw1_12_, DP_sw1_11_, DP_sw1_10_, 
        DP_sw1_9_, DP_sw1_8_, DP_sw1_7_, DP_sw1_6_, DP_sw1_5_, DP_sw1_4_, 
        DP_sw1_3_, DP_sw1_2_, DP_sw1_1_, DP_sw1_0_}), .PRODUCT({
        DP_sw1_coeff_ret1[23], SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, DP_sw1_coeff_ret1[22], 
        DP_sw1_coeff_ret1[21], DP_sw1_coeff_ret1[20], DP_sw1_coeff_ret1[19], 
        DP_sw1_coeff_ret1[18], DP_sw1_coeff_ret1[17], DP_sw1_coeff_ret1[16], 
        DP_sw1_coeff_ret1[15], DP_sw1_coeff_ret1[14], DP_sw1_coeff_ret1[13], 
        DP_sw1_coeff_ret1[12], DP_sw1_coeff_ret1[11], DP_sw1_coeff_ret1[10], 
        DP_sw1_coeff_ret1[9], DP_sw1_coeff_ret1[8], DP_sw1_coeff_ret1[7], 
        DP_sw1_coeff_ret1[6], DP_sw1_coeff_ret1[5], DP_sw1_coeff_ret1[4], 
        DP_sw1_coeff_ret1[3], DP_sw1_coeff_ret1[2], DP_sw1_coeff_ret1[1], 
        DP_sw1_coeff_ret1[0], SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130}), .TC(1'b1) );
  iir_filter_DW02_mult_5 DP_mult_204 ( .A({DP_coeffs_fb_int[0], 
        DP_coeffs_fb_int[1], DP_coeffs_fb_int[2], DP_coeffs_fb_int[3], 
        DP_coeffs_fb_int[4], DP_coeffs_fb_int[5], DP_coeffs_fb_int[6], 
        DP_coeffs_fb_int[7], DP_coeffs_fb_int[8], DP_coeffs_fb_int[9], 
        DP_coeffs_fb_int[10], DP_coeffs_fb_int[11], DP_coeffs_fb_int[12], 
        DP_coeffs_fb_int[13], DP_coeffs_fb_int[14], DP_coeffs_fb_int[15], 
        DP_coeffs_fb_int[16], DP_coeffs_fb_int[17], DP_coeffs_fb_int[18], 
        DP_coeffs_fb_int[19], DP_coeffs_fb_int[20], DP_coeffs_fb_int[21], 
        DP_coeffs_fb_int[22], DP_coeffs_fb_int[23]}), .B({DP_sw0_23_, 
        DP_sw0_22_, DP_sw0_21_, DP_sw0_20_, DP_sw0_19_, DP_sw0_18_, DP_sw0_17_, 
        DP_sw0_16_, DP_sw0_15_, DP_sw0_14_, DP_sw0_13_, DP_sw0_12_, DP_sw0_11_, 
        DP_sw0_10_, DP_sw0_9_, DP_sw0_8_, DP_sw0_7_, DP_sw0_6_, DP_sw0_5_, 
        DP_sw0_4_, DP_sw0_3_, DP_sw0_2_, DP_sw0_1_, DP_sw0_0_}), .PRODUCT({
        DP_sw0_coeff_ret0[23], SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, DP_sw0_coeff_ret0[22], 
        DP_sw0_coeff_ret0[21], DP_sw0_coeff_ret0[20], DP_sw0_coeff_ret0[19], 
        DP_sw0_coeff_ret0[18], DP_sw0_coeff_ret0[17], DP_sw0_coeff_ret0[16], 
        DP_sw0_coeff_ret0[15], DP_sw0_coeff_ret0[14], DP_sw0_coeff_ret0[13], 
        DP_sw0_coeff_ret0[12], DP_sw0_coeff_ret0[11], DP_sw0_coeff_ret0[10], 
        DP_sw0_coeff_ret0[9], DP_sw0_coeff_ret0[8], DP_sw0_coeff_ret0[7], 
        DP_sw0_coeff_ret0[6], DP_sw0_coeff_ret0[5], DP_sw0_coeff_ret0[4], 
        DP_sw0_coeff_ret0[3], DP_sw0_coeff_ret0[2], DP_sw0_coeff_ret0[1], 
        DP_sw0_coeff_ret0[0], SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154}), .TC(1'b1) );
  INV_X1 U504 ( .A(n1048), .ZN(n1032) );
  BUF_X1 U505 ( .A(n1050), .Z(n1048) );
  BUF_X1 U506 ( .A(n1057), .Z(n1035) );
  BUF_X1 U507 ( .A(n1056), .Z(n1036) );
  BUF_X1 U508 ( .A(n1057), .Z(n1034) );
  BUF_X1 U509 ( .A(n1056), .Z(n1037) );
  BUF_X1 U510 ( .A(n1055), .Z(n1038) );
  BUF_X1 U511 ( .A(n1051), .Z(n1047) );
  BUF_X1 U512 ( .A(n1051), .Z(n1046) );
  BUF_X1 U513 ( .A(n1052), .Z(n1045) );
  BUF_X1 U514 ( .A(n1053), .Z(n1043) );
  BUF_X1 U515 ( .A(n1052), .Z(n1044) );
  BUF_X1 U516 ( .A(n1053), .Z(n1042) );
  BUF_X1 U517 ( .A(n1054), .Z(n1041) );
  BUF_X1 U518 ( .A(n1055), .Z(n1039) );
  BUF_X1 U519 ( .A(n1054), .Z(n1040) );
  BUF_X1 U520 ( .A(n1050), .Z(n1049) );
  BUF_X1 U521 ( .A(n1088), .Z(n1062) );
  BUF_X1 U522 ( .A(n1088), .Z(n1063) );
  BUF_X1 U523 ( .A(n1088), .Z(n1064) );
  BUF_X1 U524 ( .A(n1088), .Z(n1065) );
  BUF_X1 U525 ( .A(n1087), .Z(n1068) );
  BUF_X1 U526 ( .A(n1087), .Z(n1069) );
  BUF_X1 U527 ( .A(n1087), .Z(n1071) );
  BUF_X1 U528 ( .A(n1087), .Z(n1070) );
  BUF_X1 U529 ( .A(n1088), .Z(n1067) );
  BUF_X1 U530 ( .A(n1088), .Z(n1066) );
  BUF_X1 U531 ( .A(n1089), .Z(n1060) );
  BUF_X1 U532 ( .A(n1089), .Z(n1061) );
  BUF_X1 U533 ( .A(n1086), .Z(n1079) );
  BUF_X1 U534 ( .A(n1086), .Z(n1078) );
  BUF_X1 U535 ( .A(n1086), .Z(n1077) );
  BUF_X1 U536 ( .A(n1086), .Z(n1074) );
  BUF_X1 U537 ( .A(n1087), .Z(n1073) );
  BUF_X1 U538 ( .A(n1086), .Z(n1075) );
  BUF_X1 U539 ( .A(n1086), .Z(n1076) );
  BUF_X1 U540 ( .A(n1085), .Z(n1083) );
  BUF_X1 U541 ( .A(n1085), .Z(n1082) );
  BUF_X1 U542 ( .A(n1085), .Z(n1081) );
  BUF_X1 U543 ( .A(n1085), .Z(n1080) );
  BUF_X1 U544 ( .A(n1085), .Z(n1084) );
  BUF_X1 U545 ( .A(n1087), .Z(n1072) );
  BUF_X1 U546 ( .A(n1028), .Z(n1050) );
  BUF_X1 U547 ( .A(n1028), .Z(n1051) );
  BUF_X1 U548 ( .A(n1028), .Z(n1052) );
  BUF_X1 U549 ( .A(n1029), .Z(n1053) );
  BUF_X1 U550 ( .A(n1029), .Z(n1055) );
  BUF_X1 U551 ( .A(n1029), .Z(n1054) );
  BUF_X1 U552 ( .A(n1030), .Z(n1057) );
  BUF_X1 U553 ( .A(n1030), .Z(n1056) );
  BUF_X1 U554 ( .A(n1090), .Z(n1087) );
  BUF_X1 U555 ( .A(n1090), .Z(n1088) );
  BUF_X1 U556 ( .A(n1091), .Z(n1086) );
  BUF_X1 U557 ( .A(n1091), .Z(n1085) );
  BUF_X1 U558 ( .A(n1090), .Z(n1089) );
  BUF_X1 U559 ( .A(n74), .Z(n1028) );
  BUF_X1 U560 ( .A(n74), .Z(n1029) );
  BUF_X1 U561 ( .A(n74), .Z(n1030) );
  NAND2_X1 U562 ( .A1(delayed_controls_2__0_), .A2(DP_N2), .ZN(n60) );
  OR2_X1 U563 ( .A1(n1027), .A2(DP_N4), .ZN(n58) );
  OAI221_X1 U564 ( .B1(n58), .B2(n59), .C1(delayed_controls_2__0_), .C2(n302), 
        .A(n60), .ZN(n520) );
  INV_X1 U565 ( .A(DP_y_0_), .ZN(n59) );
  OAI221_X1 U566 ( .B1(n58), .B2(n61), .C1(delayed_controls_2__0_), .C2(n303), 
        .A(n60), .ZN(n521) );
  INV_X1 U567 ( .A(DP_y_1_), .ZN(n61) );
  OAI221_X1 U568 ( .B1(n58), .B2(n62), .C1(delayed_controls_2__0_), .C2(n304), 
        .A(n60), .ZN(n522) );
  INV_X1 U569 ( .A(DP_y_2_), .ZN(n62) );
  OAI221_X1 U570 ( .B1(n58), .B2(n63), .C1(delayed_controls_2__0_), .C2(n305), 
        .A(n60), .ZN(n523) );
  INV_X1 U571 ( .A(DP_y_3_), .ZN(n63) );
  OAI221_X1 U572 ( .B1(n58), .B2(n64), .C1(delayed_controls_2__0_), .C2(n306), 
        .A(n60), .ZN(n524) );
  INV_X1 U573 ( .A(DP_y_4_), .ZN(n64) );
  OAI221_X1 U574 ( .B1(n58), .B2(n65), .C1(delayed_controls_2__0_), .C2(n307), 
        .A(n60), .ZN(n525) );
  INV_X1 U575 ( .A(DP_y_5_), .ZN(n65) );
  OAI221_X1 U576 ( .B1(n58), .B2(n66), .C1(delayed_controls_2__0_), .C2(n308), 
        .A(n60), .ZN(n526) );
  INV_X1 U577 ( .A(DP_y_6_), .ZN(n66) );
  OAI221_X1 U578 ( .B1(n58), .B2(n67), .C1(delayed_controls_2__0_), .C2(n309), 
        .A(n60), .ZN(n527) );
  INV_X1 U579 ( .A(DP_y_7_), .ZN(n67) );
  OAI221_X1 U580 ( .B1(n58), .B2(n68), .C1(delayed_controls_2__0_), .C2(n310), 
        .A(n60), .ZN(n528) );
  INV_X1 U581 ( .A(DP_y_8_), .ZN(n68) );
  OAI221_X1 U582 ( .B1(n58), .B2(n69), .C1(delayed_controls_2__0_), .C2(n311), 
        .A(n60), .ZN(n529) );
  INV_X1 U583 ( .A(DP_y_9_), .ZN(n69) );
  OAI221_X1 U584 ( .B1(n58), .B2(n70), .C1(delayed_controls_2__0_), .C2(n312), 
        .A(n60), .ZN(n530) );
  INV_X1 U585 ( .A(DP_y_10_), .ZN(n70) );
  INV_X1 U586 ( .A(n102), .ZN(n712) );
  AOI22_X1 U587 ( .A1(n1033), .A2(DP_w_22_), .B1(n1047), .B2(DP_sw0_22_), .ZN(
        n102) );
  INV_X1 U588 ( .A(n104), .ZN(n717) );
  AOI22_X1 U589 ( .A1(n1032), .A2(DP_w_21_), .B1(n1047), .B2(DP_sw0_21_), .ZN(
        n104) );
  INV_X1 U590 ( .A(n106), .ZN(n722) );
  AOI22_X1 U591 ( .A1(n1032), .A2(DP_w_20_), .B1(n1046), .B2(DP_sw0_20_), .ZN(
        n106) );
  INV_X1 U592 ( .A(n100), .ZN(n707) );
  AOI22_X1 U593 ( .A1(n1032), .A2(DP_w_23_), .B1(n1048), .B2(DP_sw0_23_), .ZN(
        n100) );
  OAI21_X1 U594 ( .B1(delayed_controls_2__0_), .B2(n313), .A(n72), .ZN(n531)
         );
  OAI211_X1 U595 ( .C1(DP_N4), .C2(DP_y_23), .A(n73), .B(
        delayed_controls_2__0_), .ZN(n72) );
  INV_X1 U596 ( .A(DP_N2), .ZN(n73) );
  INV_X1 U597 ( .A(n110), .ZN(n732) );
  AOI22_X1 U598 ( .A1(n1033), .A2(DP_w_18_), .B1(n1046), .B2(DP_sw0_18_), .ZN(
        n110) );
  INV_X1 U599 ( .A(n112), .ZN(n737) );
  AOI22_X1 U600 ( .A1(n1031), .A2(DP_w_17_), .B1(n1045), .B2(DP_sw0_17_), .ZN(
        n112) );
  INV_X1 U601 ( .A(n118), .ZN(n752) );
  AOI22_X1 U602 ( .A1(n1032), .A2(DP_w_14_), .B1(n1044), .B2(DP_sw0_14_), .ZN(
        n118) );
  INV_X1 U603 ( .A(n108), .ZN(n727) );
  AOI22_X1 U604 ( .A1(n1031), .A2(DP_w_19_), .B1(n1046), .B2(DP_sw0_19_), .ZN(
        n108) );
  INV_X1 U605 ( .A(n114), .ZN(n742) );
  AOI22_X1 U606 ( .A1(n1033), .A2(DP_w_16_), .B1(n1045), .B2(DP_sw0_16_), .ZN(
        n114) );
  INV_X1 U607 ( .A(n116), .ZN(n747) );
  AOI22_X1 U608 ( .A1(n1031), .A2(DP_w_15_), .B1(n1044), .B2(DP_sw0_15_), .ZN(
        n116) );
  INV_X1 U609 ( .A(n120), .ZN(n757) );
  AOI22_X1 U610 ( .A1(n1032), .A2(DP_w_13_), .B1(n1043), .B2(DP_sw0_13_), .ZN(
        n120) );
  INV_X1 U611 ( .A(n122), .ZN(n762) );
  AOI22_X1 U612 ( .A1(n1033), .A2(DP_w_12_), .B1(n1043), .B2(DP_sw0_12_), .ZN(
        n122) );
  INV_X1 U613 ( .A(n124), .ZN(n767) );
  AOI22_X1 U614 ( .A1(n1033), .A2(DP_w_11_), .B1(n1043), .B2(DP_sw0_11_), .ZN(
        n124) );
  INV_X1 U615 ( .A(n126), .ZN(n772) );
  AOI22_X1 U616 ( .A1(n1032), .A2(DP_w_10_), .B1(n1042), .B2(DP_sw0_10_), .ZN(
        n126) );
  INV_X1 U617 ( .A(n128), .ZN(n777) );
  AOI22_X1 U618 ( .A1(n1032), .A2(DP_w_9_), .B1(n1044), .B2(DP_sw0_9_), .ZN(
        n128) );
  INV_X1 U619 ( .A(n101), .ZN(n711) );
  AOI22_X1 U620 ( .A1(n1032), .A2(DP_sw0_22_), .B1(n1047), .B2(DP_sw1_22_), 
        .ZN(n101) );
  INV_X1 U621 ( .A(n103), .ZN(n716) );
  AOI22_X1 U622 ( .A1(n1031), .A2(DP_sw0_21_), .B1(n1047), .B2(DP_sw1_21_), 
        .ZN(n103) );
  INV_X1 U623 ( .A(n105), .ZN(n721) );
  AOI22_X1 U624 ( .A1(n1032), .A2(DP_sw0_20_), .B1(n1047), .B2(DP_sw1_20_), 
        .ZN(n105) );
  INV_X1 U625 ( .A(n107), .ZN(n726) );
  AOI22_X1 U626 ( .A1(n1032), .A2(DP_sw0_19_), .B1(n1046), .B2(DP_sw1_19_), 
        .ZN(n107) );
  INV_X1 U627 ( .A(n109), .ZN(n731) );
  AOI22_X1 U628 ( .A1(n1031), .A2(DP_sw0_18_), .B1(n1046), .B2(DP_sw1_18_), 
        .ZN(n109) );
  INV_X1 U629 ( .A(n111), .ZN(n736) );
  AOI22_X1 U630 ( .A1(n1033), .A2(DP_sw0_17_), .B1(n1045), .B2(DP_sw1_17_), 
        .ZN(n111) );
  INV_X1 U631 ( .A(n113), .ZN(n741) );
  AOI22_X1 U632 ( .A1(n1032), .A2(DP_sw0_16_), .B1(n1045), .B2(DP_sw1_16_), 
        .ZN(n113) );
  INV_X1 U633 ( .A(n115), .ZN(n746) );
  AOI22_X1 U634 ( .A1(n1033), .A2(DP_sw0_15_), .B1(n1045), .B2(DP_sw1_15_), 
        .ZN(n115) );
  INV_X1 U635 ( .A(n117), .ZN(n751) );
  AOI22_X1 U636 ( .A1(n1032), .A2(DP_sw0_14_), .B1(n1044), .B2(DP_sw1_14_), 
        .ZN(n117) );
  INV_X1 U637 ( .A(n119), .ZN(n756) );
  AOI22_X1 U638 ( .A1(n1032), .A2(DP_sw0_13_), .B1(n1044), .B2(DP_sw1_13_), 
        .ZN(n119) );
  INV_X1 U639 ( .A(n121), .ZN(n761) );
  AOI22_X1 U640 ( .A1(n1033), .A2(DP_sw0_12_), .B1(n1043), .B2(DP_sw1_12_), 
        .ZN(n121) );
  INV_X1 U641 ( .A(n125), .ZN(n771) );
  AOI22_X1 U642 ( .A1(n1032), .A2(DP_sw0_10_), .B1(n1042), .B2(DP_sw1_10_), 
        .ZN(n125) );
  INV_X1 U643 ( .A(n127), .ZN(n776) );
  AOI22_X1 U644 ( .A1(n1032), .A2(DP_sw0_9_), .B1(n1042), .B2(DP_sw1_9_), .ZN(
        n127) );
  INV_X1 U645 ( .A(n129), .ZN(n781) );
  AOI22_X1 U646 ( .A1(n1032), .A2(DP_sw0_8_), .B1(n1042), .B2(DP_sw1_8_), .ZN(
        n129) );
  INV_X1 U647 ( .A(n131), .ZN(n786) );
  AOI22_X1 U648 ( .A1(n1031), .A2(DP_sw0_7_), .B1(n1041), .B2(DP_sw1_7_), .ZN(
        n131) );
  INV_X1 U649 ( .A(n133), .ZN(n791) );
  AOI22_X1 U650 ( .A1(n1032), .A2(DP_sw0_6_), .B1(n1041), .B2(DP_sw1_6_), .ZN(
        n133) );
  INV_X1 U651 ( .A(n135), .ZN(n796) );
  AOI22_X1 U652 ( .A1(n1032), .A2(DP_sw0_5_), .B1(n1041), .B2(DP_sw1_5_), .ZN(
        n135) );
  OAI22_X1 U653 ( .A1(n1034), .A2(n1003), .B1(n1031), .B2(n316), .ZN(n560) );
  OAI22_X1 U654 ( .A1(n1034), .A2(n1025), .B1(n1031), .B2(n317), .ZN(n562) );
  OAI22_X1 U655 ( .A1(n1035), .A2(n1007), .B1(n1031), .B2(n318), .ZN(n564) );
  OAI22_X1 U656 ( .A1(n1034), .A2(n1008), .B1(n1031), .B2(n319), .ZN(n566) );
  OAI22_X1 U657 ( .A1(n1035), .A2(n1009), .B1(n1031), .B2(n320), .ZN(n568) );
  OAI22_X1 U658 ( .A1(n1035), .A2(n1010), .B1(n1031), .B2(n321), .ZN(n570) );
  OAI22_X1 U659 ( .A1(n1035), .A2(n1011), .B1(n1031), .B2(n322), .ZN(n572) );
  OAI22_X1 U660 ( .A1(n1035), .A2(n1012), .B1(n1031), .B2(n323), .ZN(n574) );
  OAI22_X1 U661 ( .A1(n1036), .A2(n1013), .B1(n1031), .B2(n324), .ZN(n576) );
  OAI22_X1 U662 ( .A1(n1036), .A2(n1014), .B1(n1031), .B2(n325), .ZN(n578) );
  OAI22_X1 U663 ( .A1(n1036), .A2(n1015), .B1(n1031), .B2(n326), .ZN(n580) );
  OAI22_X1 U664 ( .A1(n1036), .A2(n1016), .B1(n1031), .B2(n327), .ZN(n582) );
  INV_X1 U665 ( .A(n134), .ZN(n792) );
  AOI22_X1 U666 ( .A1(n1032), .A2(DP_w_6_), .B1(n1041), .B2(DP_sw0_6_), .ZN(
        n134) );
  INV_X1 U667 ( .A(n136), .ZN(n797) );
  AOI22_X1 U668 ( .A1(n1032), .A2(DP_w_5_), .B1(n1040), .B2(DP_sw0_5_), .ZN(
        n136) );
  INV_X1 U669 ( .A(n138), .ZN(n802) );
  AOI22_X1 U670 ( .A1(n1033), .A2(DP_w_4_), .B1(n1040), .B2(DP_sw0_4_), .ZN(
        n138) );
  OAI22_X1 U671 ( .A1(n1037), .A2(n1017), .B1(n1032), .B2(n328), .ZN(n584) );
  OAI22_X1 U672 ( .A1(n1034), .A2(n1018), .B1(n1031), .B2(n329), .ZN(n586) );
  OAI22_X1 U673 ( .A1(n1037), .A2(n1019), .B1(n1031), .B2(n330), .ZN(n588) );
  OAI22_X1 U674 ( .A1(n1036), .A2(n1020), .B1(n1033), .B2(n331), .ZN(n590) );
  OAI22_X1 U675 ( .A1(n1037), .A2(n1021), .B1(n1033), .B2(n332), .ZN(n592) );
  OAI22_X1 U676 ( .A1(n1038), .A2(n1022), .B1(n1032), .B2(n333), .ZN(n594) );
  OAI22_X1 U677 ( .A1(n1038), .A2(n1023), .B1(n1033), .B2(n334), .ZN(n596) );
  OAI22_X1 U678 ( .A1(n1037), .A2(n1024), .B1(n1031), .B2(n335), .ZN(n598) );
  OAI22_X1 U679 ( .A1(n1038), .A2(n1005), .B1(n1031), .B2(n336), .ZN(n600) );
  OAI22_X1 U680 ( .A1(n1034), .A2(n1006), .B1(n1031), .B2(n337), .ZN(n602) );
  OAI22_X1 U681 ( .A1(n1038), .A2(n1004), .B1(n1031), .B2(n338), .ZN(n604) );
  OAI22_X1 U682 ( .A1(n1037), .A2(n1059), .B1(n1032), .B2(n339), .ZN(n606) );
  OAI22_X1 U683 ( .A1(n1038), .A2(n1026), .B1(n1031), .B2(n1003), .ZN(n846) );
  OAI21_X1 U684 ( .B1(n1075), .B2(n389), .A(n147), .ZN(n847) );
  NAND2_X1 U685 ( .A1(coeffs_ff[23]), .A2(n1066), .ZN(n147) );
  OAI21_X1 U686 ( .B1(n1075), .B2(n390), .A(n148), .ZN(n848) );
  NAND2_X1 U687 ( .A1(coeffs_ff[22]), .A2(n1066), .ZN(n148) );
  OAI21_X1 U688 ( .B1(n1074), .B2(n391), .A(n149), .ZN(n849) );
  NAND2_X1 U689 ( .A1(coeffs_ff[21]), .A2(n1065), .ZN(n149) );
  OAI21_X1 U690 ( .B1(n1074), .B2(n392), .A(n150), .ZN(n850) );
  NAND2_X1 U691 ( .A1(coeffs_ff[20]), .A2(n1065), .ZN(n150) );
  OAI21_X1 U692 ( .B1(n1074), .B2(n393), .A(n151), .ZN(n851) );
  NAND2_X1 U693 ( .A1(coeffs_ff[19]), .A2(n1065), .ZN(n151) );
  OAI21_X1 U694 ( .B1(n1073), .B2(n394), .A(n152), .ZN(n852) );
  NAND2_X1 U695 ( .A1(coeffs_ff[18]), .A2(n1065), .ZN(n152) );
  OAI21_X1 U696 ( .B1(n1073), .B2(n395), .A(n153), .ZN(n853) );
  NAND2_X1 U697 ( .A1(coeffs_ff[17]), .A2(n1064), .ZN(n153) );
  OAI21_X1 U698 ( .B1(n1073), .B2(n396), .A(n154), .ZN(n854) );
  NAND2_X1 U699 ( .A1(coeffs_ff[16]), .A2(n1064), .ZN(n154) );
  OAI21_X1 U700 ( .B1(n1073), .B2(n397), .A(n155), .ZN(n855) );
  NAND2_X1 U701 ( .A1(coeffs_ff[15]), .A2(n1064), .ZN(n155) );
  OAI21_X1 U702 ( .B1(n1073), .B2(n398), .A(n156), .ZN(n856) );
  NAND2_X1 U703 ( .A1(coeffs_ff[14]), .A2(n1064), .ZN(n156) );
  OAI21_X1 U704 ( .B1(n1074), .B2(n399), .A(n157), .ZN(n857) );
  NAND2_X1 U705 ( .A1(coeffs_ff[13]), .A2(n1063), .ZN(n157) );
  OAI21_X1 U706 ( .B1(n1073), .B2(n400), .A(n158), .ZN(n858) );
  NAND2_X1 U707 ( .A1(coeffs_ff[12]), .A2(n1063), .ZN(n158) );
  OAI21_X1 U708 ( .B1(n1073), .B2(n401), .A(n159), .ZN(n859) );
  NAND2_X1 U709 ( .A1(coeffs_ff[11]), .A2(n1063), .ZN(n159) );
  OAI21_X1 U710 ( .B1(n1074), .B2(n402), .A(n160), .ZN(n860) );
  NAND2_X1 U711 ( .A1(coeffs_ff[10]), .A2(n1063), .ZN(n160) );
  OAI21_X1 U712 ( .B1(n1074), .B2(n403), .A(n161), .ZN(n861) );
  NAND2_X1 U713 ( .A1(coeffs_ff[9]), .A2(n1062), .ZN(n161) );
  OAI21_X1 U714 ( .B1(n1074), .B2(n404), .A(n162), .ZN(n862) );
  NAND2_X1 U715 ( .A1(coeffs_ff[8]), .A2(n1062), .ZN(n162) );
  OAI21_X1 U716 ( .B1(n1074), .B2(n405), .A(n163), .ZN(n863) );
  NAND2_X1 U717 ( .A1(coeffs_ff[7]), .A2(n1062), .ZN(n163) );
  OAI21_X1 U718 ( .B1(n1074), .B2(n406), .A(n164), .ZN(n864) );
  NAND2_X1 U719 ( .A1(coeffs_ff[6]), .A2(n1062), .ZN(n164) );
  OAI21_X1 U720 ( .B1(n1074), .B2(n407), .A(n165), .ZN(n865) );
  NAND2_X1 U721 ( .A1(coeffs_ff[5]), .A2(n1061), .ZN(n165) );
  OAI21_X1 U722 ( .B1(n1076), .B2(n408), .A(n166), .ZN(n866) );
  NAND2_X1 U723 ( .A1(coeffs_ff[4]), .A2(n1061), .ZN(n166) );
  OAI21_X1 U724 ( .B1(n1075), .B2(n409), .A(n167), .ZN(n867) );
  NAND2_X1 U725 ( .A1(coeffs_ff[3]), .A2(n1061), .ZN(n167) );
  OAI21_X1 U726 ( .B1(n1075), .B2(n410), .A(n168), .ZN(n868) );
  NAND2_X1 U727 ( .A1(coeffs_ff[2]), .A2(n1061), .ZN(n168) );
  OAI21_X1 U728 ( .B1(n1075), .B2(n411), .A(n169), .ZN(n869) );
  NAND2_X1 U729 ( .A1(coeffs_ff[1]), .A2(n1060), .ZN(n169) );
  OAI21_X1 U730 ( .B1(n1076), .B2(n412), .A(n170), .ZN(n870) );
  NAND2_X1 U731 ( .A1(coeffs_ff[0]), .A2(n1060), .ZN(n170) );
  OAI21_X1 U732 ( .B1(n1076), .B2(n413), .A(n171), .ZN(n871) );
  NAND2_X1 U733 ( .A1(coeffs_ff[47]), .A2(n1060), .ZN(n171) );
  OAI21_X1 U734 ( .B1(n1076), .B2(n414), .A(n172), .ZN(n872) );
  NAND2_X1 U735 ( .A1(coeffs_ff[46]), .A2(n1060), .ZN(n172) );
  OAI21_X1 U736 ( .B1(n1076), .B2(n415), .A(n173), .ZN(n873) );
  NAND2_X1 U737 ( .A1(coeffs_ff[45]), .A2(n1061), .ZN(n173) );
  OAI21_X1 U738 ( .B1(n1079), .B2(n479), .A(n237), .ZN(n937) );
  NAND2_X1 U739 ( .A1(coeffs_ff[77]), .A2(n1071), .ZN(n237) );
  OAI21_X1 U740 ( .B1(n1079), .B2(n480), .A(n238), .ZN(n938) );
  NAND2_X1 U741 ( .A1(coeffs_ff[76]), .A2(n1071), .ZN(n238) );
  OAI21_X1 U742 ( .B1(n1079), .B2(n481), .A(n239), .ZN(n939) );
  NAND2_X1 U743 ( .A1(coeffs_ff[75]), .A2(n1072), .ZN(n239) );
  OAI21_X1 U744 ( .B1(n1079), .B2(n482), .A(n240), .ZN(n940) );
  NAND2_X1 U745 ( .A1(coeffs_ff[74]), .A2(n1072), .ZN(n240) );
  OAI21_X1 U746 ( .B1(n1079), .B2(n483), .A(n241), .ZN(n941) );
  NAND2_X1 U747 ( .A1(coeffs_ff[73]), .A2(n1072), .ZN(n241) );
  OAI21_X1 U748 ( .B1(n1079), .B2(n484), .A(n242), .ZN(n942) );
  NAND2_X1 U749 ( .A1(coeffs_ff[72]), .A2(n1071), .ZN(n242) );
  OAI21_X1 U750 ( .B1(n1079), .B2(n485), .A(n243), .ZN(n943) );
  NAND2_X1 U751 ( .A1(coeffs_fb[23]), .A2(n1071), .ZN(n243) );
  OAI21_X1 U752 ( .B1(n1079), .B2(n486), .A(n244), .ZN(n944) );
  NAND2_X1 U753 ( .A1(coeffs_fb[22]), .A2(n1071), .ZN(n244) );
  OAI21_X1 U754 ( .B1(n1079), .B2(n487), .A(n245), .ZN(n945) );
  NAND2_X1 U755 ( .A1(coeffs_fb[21]), .A2(n1071), .ZN(n245) );
  OAI21_X1 U756 ( .B1(n1079), .B2(n488), .A(n246), .ZN(n946) );
  NAND2_X1 U757 ( .A1(coeffs_fb[20]), .A2(n1071), .ZN(n246) );
  OAI21_X1 U758 ( .B1(n1079), .B2(n489), .A(n247), .ZN(n947) );
  NAND2_X1 U759 ( .A1(coeffs_fb[19]), .A2(n1071), .ZN(n247) );
  OAI21_X1 U760 ( .B1(n1079), .B2(n490), .A(n248), .ZN(n948) );
  NAND2_X1 U761 ( .A1(coeffs_fb[18]), .A2(n1071), .ZN(n248) );
  OAI21_X1 U762 ( .B1(n1079), .B2(n491), .A(n249), .ZN(n949) );
  NAND2_X1 U763 ( .A1(coeffs_fb[17]), .A2(n1070), .ZN(n249) );
  OAI21_X1 U764 ( .B1(n1078), .B2(n492), .A(n250), .ZN(n950) );
  NAND2_X1 U765 ( .A1(coeffs_fb[16]), .A2(n1070), .ZN(n250) );
  OAI21_X1 U766 ( .B1(n1078), .B2(n493), .A(n251), .ZN(n951) );
  NAND2_X1 U767 ( .A1(coeffs_fb[15]), .A2(n1070), .ZN(n251) );
  OAI21_X1 U768 ( .B1(n1078), .B2(n495), .A(n253), .ZN(n953) );
  NAND2_X1 U769 ( .A1(coeffs_fb[13]), .A2(n1070), .ZN(n253) );
  OAI21_X1 U770 ( .B1(n1078), .B2(n496), .A(n254), .ZN(n954) );
  NAND2_X1 U771 ( .A1(coeffs_fb[12]), .A2(n1070), .ZN(n254) );
  OAI21_X1 U772 ( .B1(n1078), .B2(n497), .A(n255), .ZN(n955) );
  NAND2_X1 U773 ( .A1(coeffs_fb[11]), .A2(n1070), .ZN(n255) );
  OAI21_X1 U774 ( .B1(n1078), .B2(n498), .A(n256), .ZN(n956) );
  NAND2_X1 U775 ( .A1(coeffs_fb[10]), .A2(n1069), .ZN(n256) );
  OAI21_X1 U776 ( .B1(n1078), .B2(n499), .A(n257), .ZN(n957) );
  NAND2_X1 U777 ( .A1(coeffs_fb[9]), .A2(n1069), .ZN(n257) );
  OAI21_X1 U778 ( .B1(n1078), .B2(n500), .A(n258), .ZN(n958) );
  NAND2_X1 U779 ( .A1(coeffs_fb[8]), .A2(n1069), .ZN(n258) );
  OAI21_X1 U780 ( .B1(n1078), .B2(n501), .A(n259), .ZN(n959) );
  NAND2_X1 U781 ( .A1(coeffs_fb[7]), .A2(n1069), .ZN(n259) );
  OAI21_X1 U782 ( .B1(n1078), .B2(n502), .A(n260), .ZN(n960) );
  NAND2_X1 U783 ( .A1(coeffs_fb[6]), .A2(n1069), .ZN(n260) );
  OAI21_X1 U784 ( .B1(n1078), .B2(n503), .A(n261), .ZN(n961) );
  NAND2_X1 U785 ( .A1(coeffs_fb[5]), .A2(n1069), .ZN(n261) );
  OAI21_X1 U786 ( .B1(n1078), .B2(n504), .A(n262), .ZN(n962) );
  NAND2_X1 U787 ( .A1(coeffs_fb[4]), .A2(n1069), .ZN(n262) );
  OAI21_X1 U788 ( .B1(n1078), .B2(n505), .A(n263), .ZN(n963) );
  NAND2_X1 U789 ( .A1(coeffs_fb[3]), .A2(n1069), .ZN(n263) );
  OAI21_X1 U790 ( .B1(n1077), .B2(n506), .A(n264), .ZN(n964) );
  NAND2_X1 U791 ( .A1(coeffs_fb[2]), .A2(n1068), .ZN(n264) );
  OAI21_X1 U792 ( .B1(n1077), .B2(n507), .A(n265), .ZN(n965) );
  NAND2_X1 U793 ( .A1(coeffs_fb[1]), .A2(n1068), .ZN(n265) );
  OAI21_X1 U794 ( .B1(n1077), .B2(n508), .A(n266), .ZN(n966) );
  NAND2_X1 U795 ( .A1(coeffs_fb[0]), .A2(n1068), .ZN(n266) );
  OAI21_X1 U796 ( .B1(n1077), .B2(n509), .A(n267), .ZN(n967) );
  NAND2_X1 U797 ( .A1(coeffs_fb[47]), .A2(n1068), .ZN(n267) );
  OAI21_X1 U798 ( .B1(n1077), .B2(n510), .A(n268), .ZN(n968) );
  NAND2_X1 U799 ( .A1(coeffs_fb[46]), .A2(n1068), .ZN(n268) );
  OAI21_X1 U800 ( .B1(n1077), .B2(n511), .A(n269), .ZN(n969) );
  NAND2_X1 U801 ( .A1(coeffs_fb[45]), .A2(n1068), .ZN(n269) );
  OAI21_X1 U802 ( .B1(n1077), .B2(n512), .A(n270), .ZN(n970) );
  NAND2_X1 U803 ( .A1(coeffs_fb[44]), .A2(n1068), .ZN(n270) );
  OAI21_X1 U804 ( .B1(n1077), .B2(n513), .A(n271), .ZN(n971) );
  NAND2_X1 U805 ( .A1(coeffs_fb[43]), .A2(n1068), .ZN(n271) );
  OAI21_X1 U806 ( .B1(n1077), .B2(n514), .A(n272), .ZN(n972) );
  NAND2_X1 U807 ( .A1(coeffs_fb[42]), .A2(n1067), .ZN(n272) );
  OAI21_X1 U808 ( .B1(n1077), .B2(n515), .A(n273), .ZN(n973) );
  NAND2_X1 U809 ( .A1(coeffs_fb[41]), .A2(n1067), .ZN(n273) );
  OAI21_X1 U810 ( .B1(n1077), .B2(n516), .A(n274), .ZN(n974) );
  NAND2_X1 U811 ( .A1(coeffs_fb[40]), .A2(n1067), .ZN(n274) );
  OAI21_X1 U812 ( .B1(n1077), .B2(n517), .A(n275), .ZN(n975) );
  NAND2_X1 U813 ( .A1(coeffs_fb[39]), .A2(n1067), .ZN(n275) );
  OAI21_X1 U814 ( .B1(n1077), .B2(n518), .A(n276), .ZN(n976) );
  NAND2_X1 U815 ( .A1(coeffs_fb[38]), .A2(n1067), .ZN(n276) );
  OAI21_X1 U816 ( .B1(n1075), .B2(n277), .A(n33), .ZN(n978) );
  NAND2_X1 U817 ( .A1(coeffs_fb[36]), .A2(n1067), .ZN(n33) );
  OAI21_X1 U818 ( .B1(n1076), .B2(n278), .A(n34), .ZN(n979) );
  NAND2_X1 U819 ( .A1(coeffs_fb[35]), .A2(n1067), .ZN(n34) );
  OAI21_X1 U820 ( .B1(n1076), .B2(n279), .A(n35), .ZN(n980) );
  NAND2_X1 U821 ( .A1(coeffs_fb[34]), .A2(n1068), .ZN(n35) );
  OAI21_X1 U822 ( .B1(n1076), .B2(n280), .A(n36), .ZN(n981) );
  NAND2_X1 U823 ( .A1(coeffs_fb[33]), .A2(n1068), .ZN(n36) );
  OAI21_X1 U824 ( .B1(n1075), .B2(n281), .A(n37), .ZN(n982) );
  NAND2_X1 U825 ( .A1(coeffs_fb[32]), .A2(n1068), .ZN(n37) );
  OAI21_X1 U826 ( .B1(n1075), .B2(n282), .A(n38), .ZN(n983) );
  NAND2_X1 U827 ( .A1(coeffs_fb[31]), .A2(n1068), .ZN(n38) );
  OAI21_X1 U828 ( .B1(n1075), .B2(n283), .A(n39), .ZN(n984) );
  NAND2_X1 U829 ( .A1(coeffs_fb[30]), .A2(n1069), .ZN(n39) );
  OAI21_X1 U830 ( .B1(n1074), .B2(n284), .A(n40), .ZN(n985) );
  NAND2_X1 U831 ( .A1(coeffs_fb[29]), .A2(n1069), .ZN(n40) );
  OAI21_X1 U832 ( .B1(n1074), .B2(n285), .A(n41), .ZN(n986) );
  NAND2_X1 U833 ( .A1(coeffs_fb[28]), .A2(n1069), .ZN(n41) );
  OAI21_X1 U834 ( .B1(n1074), .B2(n286), .A(n42), .ZN(n987) );
  NAND2_X1 U835 ( .A1(coeffs_fb[27]), .A2(n1069), .ZN(n42) );
  OAI21_X1 U836 ( .B1(n1073), .B2(n287), .A(n43), .ZN(n988) );
  NAND2_X1 U837 ( .A1(coeffs_fb[26]), .A2(n1070), .ZN(n43) );
  OAI21_X1 U838 ( .B1(n1073), .B2(n288), .A(n44), .ZN(n989) );
  NAND2_X1 U839 ( .A1(coeffs_fb[25]), .A2(n1070), .ZN(n44) );
  OAI21_X1 U840 ( .B1(n1073), .B2(n289), .A(n45), .ZN(n990) );
  NAND2_X1 U841 ( .A1(coeffs_fb[24]), .A2(n1070), .ZN(n45) );
  OAI21_X1 U842 ( .B1(n1073), .B2(n290), .A(n46), .ZN(n991) );
  NAND2_X1 U843 ( .A1(dIn[11]), .A2(n1070), .ZN(n46) );
  OAI21_X1 U844 ( .B1(n1073), .B2(n292), .A(n48), .ZN(n993) );
  NAND2_X1 U845 ( .A1(dIn[9]), .A2(n1071), .ZN(n48) );
  OAI21_X1 U846 ( .B1(n1073), .B2(n293), .A(n49), .ZN(n994) );
  NAND2_X1 U847 ( .A1(dIn[8]), .A2(n1071), .ZN(n49) );
  OAI21_X1 U848 ( .B1(n1075), .B2(n294), .A(n50), .ZN(n995) );
  NAND2_X1 U849 ( .A1(dIn[7]), .A2(n1072), .ZN(n50) );
  OAI21_X1 U850 ( .B1(n1075), .B2(n295), .A(n51), .ZN(n996) );
  NAND2_X1 U851 ( .A1(dIn[6]), .A2(n1072), .ZN(n51) );
  OAI21_X1 U852 ( .B1(n1075), .B2(n296), .A(n52), .ZN(n997) );
  NAND2_X1 U853 ( .A1(dIn[5]), .A2(n1070), .ZN(n52) );
  OAI21_X1 U854 ( .B1(n1075), .B2(n297), .A(n53), .ZN(n998) );
  NAND2_X1 U855 ( .A1(dIn[4]), .A2(n1072), .ZN(n53) );
  OAI21_X1 U856 ( .B1(n1076), .B2(n298), .A(n54), .ZN(n999) );
  NAND2_X1 U857 ( .A1(dIn[3]), .A2(n1072), .ZN(n54) );
  OAI21_X1 U858 ( .B1(n1076), .B2(n299), .A(n55), .ZN(n1000) );
  NAND2_X1 U859 ( .A1(dIn[2]), .A2(n1067), .ZN(n55) );
  OAI21_X1 U860 ( .B1(n1076), .B2(n300), .A(n56), .ZN(n1001) );
  NAND2_X1 U861 ( .A1(dIn[1]), .A2(n1066), .ZN(n56) );
  OAI21_X1 U862 ( .B1(n1076), .B2(n301), .A(n57), .ZN(n1002) );
  NAND2_X1 U863 ( .A1(dIn[0]), .A2(n1066), .ZN(n57) );
  OAI21_X1 U864 ( .B1(n1072), .B2(n291), .A(n47), .ZN(n992) );
  NAND2_X1 U865 ( .A1(dIn[10]), .A2(n1071), .ZN(n47) );
  OAI21_X1 U866 ( .B1(n1083), .B2(n428), .A(n186), .ZN(n886) );
  NAND2_X1 U867 ( .A1(coeffs_ff[32]), .A2(n1067), .ZN(n186) );
  OAI21_X1 U868 ( .B1(n1083), .B2(n429), .A(n187), .ZN(n887) );
  NAND2_X1 U869 ( .A1(coeffs_ff[31]), .A2(n1061), .ZN(n187) );
  OAI21_X1 U870 ( .B1(n1083), .B2(n430), .A(n188), .ZN(n888) );
  NAND2_X1 U871 ( .A1(coeffs_ff[30]), .A2(n1061), .ZN(n188) );
  OAI21_X1 U872 ( .B1(n1083), .B2(n431), .A(n189), .ZN(n889) );
  NAND2_X1 U873 ( .A1(coeffs_ff[29]), .A2(n1061), .ZN(n189) );
  OAI21_X1 U874 ( .B1(n1083), .B2(n432), .A(n190), .ZN(n890) );
  NAND2_X1 U875 ( .A1(coeffs_ff[28]), .A2(n1062), .ZN(n190) );
  OAI21_X1 U876 ( .B1(n1083), .B2(n433), .A(n191), .ZN(n891) );
  NAND2_X1 U877 ( .A1(coeffs_ff[27]), .A2(n1062), .ZN(n191) );
  OAI21_X1 U878 ( .B1(n1083), .B2(n434), .A(n192), .ZN(n892) );
  NAND2_X1 U879 ( .A1(coeffs_ff[26]), .A2(n1062), .ZN(n192) );
  OAI21_X1 U880 ( .B1(n1083), .B2(n435), .A(n193), .ZN(n893) );
  NAND2_X1 U881 ( .A1(coeffs_ff[25]), .A2(n1062), .ZN(n193) );
  OAI21_X1 U882 ( .B1(n1083), .B2(n436), .A(n194), .ZN(n894) );
  NAND2_X1 U883 ( .A1(coeffs_ff[24]), .A2(n1062), .ZN(n194) );
  OAI21_X1 U884 ( .B1(n1083), .B2(n437), .A(n195), .ZN(n895) );
  NAND2_X1 U885 ( .A1(coeffs_ff[71]), .A2(n1062), .ZN(n195) );
  OAI21_X1 U886 ( .B1(n1083), .B2(n438), .A(n196), .ZN(n896) );
  NAND2_X1 U887 ( .A1(coeffs_ff[70]), .A2(n1062), .ZN(n196) );
  OAI21_X1 U888 ( .B1(n1083), .B2(n439), .A(n197), .ZN(n897) );
  NAND2_X1 U889 ( .A1(coeffs_ff[69]), .A2(n1062), .ZN(n197) );
  OAI21_X1 U890 ( .B1(n1083), .B2(n440), .A(n198), .ZN(n898) );
  NAND2_X1 U891 ( .A1(coeffs_ff[68]), .A2(n1063), .ZN(n198) );
  OAI21_X1 U892 ( .B1(n1082), .B2(n441), .A(n199), .ZN(n899) );
  NAND2_X1 U893 ( .A1(coeffs_ff[67]), .A2(n1063), .ZN(n199) );
  OAI21_X1 U894 ( .B1(n1082), .B2(n442), .A(n200), .ZN(n900) );
  NAND2_X1 U895 ( .A1(coeffs_ff[66]), .A2(n1063), .ZN(n200) );
  OAI21_X1 U896 ( .B1(n1082), .B2(n443), .A(n201), .ZN(n901) );
  NAND2_X1 U897 ( .A1(coeffs_ff[65]), .A2(n1063), .ZN(n201) );
  OAI21_X1 U898 ( .B1(n1082), .B2(n444), .A(n202), .ZN(n902) );
  NAND2_X1 U899 ( .A1(coeffs_ff[64]), .A2(n1063), .ZN(n202) );
  OAI21_X1 U900 ( .B1(n1082), .B2(n445), .A(n203), .ZN(n903) );
  NAND2_X1 U901 ( .A1(coeffs_ff[63]), .A2(n1063), .ZN(n203) );
  OAI21_X1 U902 ( .B1(n1082), .B2(n446), .A(n204), .ZN(n904) );
  NAND2_X1 U903 ( .A1(coeffs_ff[62]), .A2(n1063), .ZN(n204) );
  OAI21_X1 U904 ( .B1(n1082), .B2(n447), .A(n205), .ZN(n905) );
  NAND2_X1 U905 ( .A1(coeffs_ff[61]), .A2(n1063), .ZN(n205) );
  OAI21_X1 U906 ( .B1(n1082), .B2(n448), .A(n206), .ZN(n906) );
  NAND2_X1 U907 ( .A1(coeffs_ff[60]), .A2(n1064), .ZN(n206) );
  OAI21_X1 U908 ( .B1(n1082), .B2(n449), .A(n207), .ZN(n907) );
  NAND2_X1 U909 ( .A1(coeffs_ff[59]), .A2(n1064), .ZN(n207) );
  OAI21_X1 U910 ( .B1(n1082), .B2(n450), .A(n208), .ZN(n908) );
  NAND2_X1 U911 ( .A1(coeffs_ff[58]), .A2(n1064), .ZN(n208) );
  OAI21_X1 U912 ( .B1(n1082), .B2(n451), .A(n209), .ZN(n909) );
  NAND2_X1 U913 ( .A1(coeffs_ff[57]), .A2(n1064), .ZN(n209) );
  OAI21_X1 U914 ( .B1(n1082), .B2(n452), .A(n210), .ZN(n910) );
  NAND2_X1 U915 ( .A1(coeffs_ff[56]), .A2(n1064), .ZN(n210) );
  OAI21_X1 U916 ( .B1(n1082), .B2(n453), .A(n211), .ZN(n911) );
  NAND2_X1 U917 ( .A1(coeffs_ff[55]), .A2(n1064), .ZN(n211) );
  OAI21_X1 U918 ( .B1(n1081), .B2(n454), .A(n212), .ZN(n912) );
  NAND2_X1 U919 ( .A1(coeffs_ff[54]), .A2(n1064), .ZN(n212) );
  OAI21_X1 U920 ( .B1(n1081), .B2(n455), .A(n213), .ZN(n913) );
  NAND2_X1 U921 ( .A1(coeffs_ff[53]), .A2(n1064), .ZN(n213) );
  OAI21_X1 U922 ( .B1(n1081), .B2(n456), .A(n214), .ZN(n914) );
  NAND2_X1 U923 ( .A1(coeffs_ff[52]), .A2(n1065), .ZN(n214) );
  OAI21_X1 U924 ( .B1(n1081), .B2(n457), .A(n215), .ZN(n915) );
  NAND2_X1 U925 ( .A1(coeffs_ff[51]), .A2(n1065), .ZN(n215) );
  OAI21_X1 U926 ( .B1(n1081), .B2(n458), .A(n216), .ZN(n916) );
  NAND2_X1 U927 ( .A1(coeffs_ff[50]), .A2(n1065), .ZN(n216) );
  OAI21_X1 U928 ( .B1(n1081), .B2(n459), .A(n217), .ZN(n917) );
  NAND2_X1 U929 ( .A1(coeffs_ff[49]), .A2(n1065), .ZN(n217) );
  OAI21_X1 U930 ( .B1(n1081), .B2(n460), .A(n218), .ZN(n918) );
  NAND2_X1 U931 ( .A1(coeffs_ff[48]), .A2(n1065), .ZN(n218) );
  OAI21_X1 U932 ( .B1(n1081), .B2(n461), .A(n219), .ZN(n919) );
  NAND2_X1 U933 ( .A1(coeffs_ff[95]), .A2(n1065), .ZN(n219) );
  OAI21_X1 U934 ( .B1(n1081), .B2(n462), .A(n220), .ZN(n920) );
  NAND2_X1 U935 ( .A1(coeffs_ff[94]), .A2(n1065), .ZN(n220) );
  OAI21_X1 U936 ( .B1(n1081), .B2(n463), .A(n221), .ZN(n921) );
  NAND2_X1 U937 ( .A1(coeffs_ff[93]), .A2(n1065), .ZN(n221) );
  OAI21_X1 U938 ( .B1(n1081), .B2(n464), .A(n222), .ZN(n922) );
  NAND2_X1 U939 ( .A1(coeffs_ff[92]), .A2(n1066), .ZN(n222) );
  OAI21_X1 U940 ( .B1(n1081), .B2(n465), .A(n223), .ZN(n923) );
  NAND2_X1 U941 ( .A1(coeffs_ff[91]), .A2(n1066), .ZN(n223) );
  OAI21_X1 U942 ( .B1(n1081), .B2(n466), .A(n224), .ZN(n924) );
  NAND2_X1 U943 ( .A1(coeffs_ff[90]), .A2(n1066), .ZN(n224) );
  OAI21_X1 U944 ( .B1(n1080), .B2(n467), .A(n225), .ZN(n925) );
  NAND2_X1 U945 ( .A1(coeffs_ff[89]), .A2(n1066), .ZN(n225) );
  OAI21_X1 U946 ( .B1(n1080), .B2(n468), .A(n226), .ZN(n926) );
  NAND2_X1 U947 ( .A1(coeffs_ff[88]), .A2(n1066), .ZN(n226) );
  OAI21_X1 U948 ( .B1(n1080), .B2(n469), .A(n227), .ZN(n927) );
  NAND2_X1 U949 ( .A1(coeffs_ff[87]), .A2(n1066), .ZN(n227) );
  OAI21_X1 U950 ( .B1(n1080), .B2(n470), .A(n228), .ZN(n928) );
  NAND2_X1 U951 ( .A1(coeffs_ff[86]), .A2(n1066), .ZN(n228) );
  OAI21_X1 U952 ( .B1(n1080), .B2(n471), .A(n229), .ZN(n929) );
  NAND2_X1 U953 ( .A1(coeffs_ff[85]), .A2(n1066), .ZN(n229) );
  OAI21_X1 U954 ( .B1(n1080), .B2(n472), .A(n230), .ZN(n930) );
  NAND2_X1 U955 ( .A1(coeffs_ff[84]), .A2(n1067), .ZN(n230) );
  OAI21_X1 U956 ( .B1(n1080), .B2(n473), .A(n231), .ZN(n931) );
  NAND2_X1 U957 ( .A1(coeffs_ff[83]), .A2(n1067), .ZN(n231) );
  OAI21_X1 U958 ( .B1(n1080), .B2(n474), .A(n232), .ZN(n932) );
  NAND2_X1 U959 ( .A1(coeffs_ff[82]), .A2(n1067), .ZN(n232) );
  OAI21_X1 U960 ( .B1(n1080), .B2(n475), .A(n233), .ZN(n933) );
  NAND2_X1 U961 ( .A1(coeffs_ff[81]), .A2(n1072), .ZN(n233) );
  OAI21_X1 U962 ( .B1(n1080), .B2(n476), .A(n234), .ZN(n934) );
  NAND2_X1 U963 ( .A1(coeffs_ff[80]), .A2(n1072), .ZN(n234) );
  OAI21_X1 U964 ( .B1(n1080), .B2(n477), .A(n235), .ZN(n935) );
  NAND2_X1 U965 ( .A1(coeffs_ff[79]), .A2(n1072), .ZN(n235) );
  OAI21_X1 U966 ( .B1(n1080), .B2(n478), .A(n236), .ZN(n936) );
  NAND2_X1 U967 ( .A1(coeffs_ff[78]), .A2(n1072), .ZN(n236) );
  OAI21_X1 U968 ( .B1(n1080), .B2(n494), .A(n252), .ZN(n952) );
  NAND2_X1 U969 ( .A1(coeffs_fb[14]), .A2(n1070), .ZN(n252) );
  OAI21_X1 U970 ( .B1(n1084), .B2(n416), .A(n174), .ZN(n874) );
  NAND2_X1 U971 ( .A1(coeffs_ff[44]), .A2(n1060), .ZN(n174) );
  OAI21_X1 U972 ( .B1(n1084), .B2(n417), .A(n175), .ZN(n875) );
  NAND2_X1 U973 ( .A1(coeffs_ff[43]), .A2(n1060), .ZN(n175) );
  OAI21_X1 U974 ( .B1(n1084), .B2(n418), .A(n176), .ZN(n876) );
  NAND2_X1 U975 ( .A1(coeffs_ff[42]), .A2(n1060), .ZN(n176) );
  OAI21_X1 U976 ( .B1(n1084), .B2(n419), .A(n177), .ZN(n877) );
  NAND2_X1 U977 ( .A1(coeffs_ff[41]), .A2(n1060), .ZN(n177) );
  OAI21_X1 U978 ( .B1(n1084), .B2(n420), .A(n178), .ZN(n878) );
  NAND2_X1 U979 ( .A1(coeffs_ff[40]), .A2(n1060), .ZN(n178) );
  OAI21_X1 U980 ( .B1(n1084), .B2(n421), .A(n179), .ZN(n879) );
  NAND2_X1 U981 ( .A1(coeffs_ff[39]), .A2(n1060), .ZN(n179) );
  OAI21_X1 U982 ( .B1(n1084), .B2(n422), .A(n180), .ZN(n880) );
  NAND2_X1 U983 ( .A1(coeffs_ff[38]), .A2(n1060), .ZN(n180) );
  OAI21_X1 U984 ( .B1(n1084), .B2(n423), .A(n181), .ZN(n881) );
  NAND2_X1 U985 ( .A1(coeffs_ff[37]), .A2(n1060), .ZN(n181) );
  OAI21_X1 U986 ( .B1(n1084), .B2(n424), .A(n182), .ZN(n882) );
  NAND2_X1 U987 ( .A1(coeffs_ff[36]), .A2(n1061), .ZN(n182) );
  OAI21_X1 U988 ( .B1(n1084), .B2(n425), .A(n183), .ZN(n883) );
  NAND2_X1 U989 ( .A1(coeffs_ff[35]), .A2(n1061), .ZN(n183) );
  OAI21_X1 U990 ( .B1(n1084), .B2(n426), .A(n184), .ZN(n884) );
  NAND2_X1 U991 ( .A1(coeffs_ff[34]), .A2(n1061), .ZN(n184) );
  OAI21_X1 U992 ( .B1(n1084), .B2(n427), .A(n185), .ZN(n885) );
  NAND2_X1 U993 ( .A1(coeffs_ff[33]), .A2(n1061), .ZN(n185) );
  OAI21_X1 U994 ( .B1(n1076), .B2(n519), .A(n32), .ZN(n977) );
  NAND2_X1 U995 ( .A1(n1084), .A2(coeffs_fb[37]), .ZN(n32) );
  INV_X1 U996 ( .A(n142), .ZN(n812) );
  AOI22_X1 U997 ( .A1(n1033), .A2(DP_w_2_), .B1(n1039), .B2(DP_sw0_2_), .ZN(
        n142) );
  INV_X1 U998 ( .A(n130), .ZN(n782) );
  AOI22_X1 U999 ( .A1(n1032), .A2(DP_w_8_), .B1(n1042), .B2(DP_sw0_8_), .ZN(
        n130) );
  INV_X1 U1000 ( .A(n132), .ZN(n787) );
  AOI22_X1 U1001 ( .A1(n1032), .A2(DP_w_7_), .B1(n1041), .B2(DP_sw0_7_), .ZN(
        n132) );
  INV_X1 U1002 ( .A(n140), .ZN(n807) );
  AOI22_X1 U1003 ( .A1(n1033), .A2(DP_w_3_), .B1(n1039), .B2(DP_sw0_3_), .ZN(
        n140) );
  INV_X1 U1004 ( .A(n141), .ZN(n811) );
  AOI22_X1 U1005 ( .A1(n1033), .A2(DP_sw0_2_), .B1(n1039), .B2(DP_sw1_2_), 
        .ZN(n141) );
  INV_X1 U1006 ( .A(n123), .ZN(n766) );
  AOI22_X1 U1007 ( .A1(n1033), .A2(DP_sw0_11_), .B1(n1043), .B2(DP_sw1_11_), 
        .ZN(n123) );
  INV_X1 U1008 ( .A(n137), .ZN(n801) );
  AOI22_X1 U1009 ( .A1(n1033), .A2(DP_sw0_4_), .B1(n1040), .B2(DP_sw1_4_), 
        .ZN(n137) );
  INV_X1 U1010 ( .A(n139), .ZN(n806) );
  AOI22_X1 U1011 ( .A1(n1033), .A2(DP_sw0_3_), .B1(n1040), .B2(DP_sw1_3_), 
        .ZN(n139) );
  BUF_X1 U1012 ( .A(vIn), .Z(n1090) );
  INV_X1 U1013 ( .A(n144), .ZN(n817) );
  AOI22_X1 U1014 ( .A1(n1033), .A2(DP_w_1_), .B1(n1039), .B2(DP_sw0_1_), .ZN(
        n144) );
  INV_X1 U1015 ( .A(n143), .ZN(n816) );
  AOI22_X1 U1016 ( .A1(n1033), .A2(DP_sw0_1_), .B1(n1039), .B2(DP_sw1_1_), 
        .ZN(n143) );
  BUF_X1 U1017 ( .A(vIn), .Z(n1091) );
  INV_X1 U1018 ( .A(n145), .ZN(n820) );
  AOI22_X1 U1019 ( .A1(n1033), .A2(DP_w_0_), .B1(n1040), .B2(DP_sw0_0_), .ZN(
        n145) );
  INV_X1 U1020 ( .A(n99), .ZN(n706) );
  AOI22_X1 U1021 ( .A1(n1033), .A2(DP_sw0_23_), .B1(n1048), .B2(n1058), .ZN(
        n99) );
  BUF_X1 U1022 ( .A(rst_n), .Z(n1133) );
  BUF_X1 U1023 ( .A(rst_n), .Z(n1134) );
  BUF_X1 U1024 ( .A(rst_n), .Z(n1135) );
  BUF_X1 U1025 ( .A(rst_n), .Z(n1136) );
  BUF_X1 U1026 ( .A(rst_n), .Z(n1137) );
  BUF_X1 U1027 ( .A(rst_n), .Z(n1138) );
  BUF_X1 U1028 ( .A(rst_n), .Z(n1139) );
  INV_X1 U1029 ( .A(n1048), .ZN(n1031) );
  INV_X1 U1030 ( .A(n1049), .ZN(n1033) );
  INV_X1 U1031 ( .A(n1059), .ZN(n1058) );
  INV_X1 U1032 ( .A(DP_sw1_23_), .ZN(n1059) );
  CLKBUF_X1 U1033 ( .A(n1139), .Z(n1092) );
  CLKBUF_X1 U1034 ( .A(n1139), .Z(n1093) );
  CLKBUF_X1 U1035 ( .A(n1139), .Z(n1094) );
  CLKBUF_X1 U1036 ( .A(n1139), .Z(n1095) );
  CLKBUF_X1 U1037 ( .A(n1139), .Z(n1096) );
  CLKBUF_X1 U1038 ( .A(n1138), .Z(n1097) );
  CLKBUF_X1 U1039 ( .A(n1138), .Z(n1098) );
  CLKBUF_X1 U1040 ( .A(n1138), .Z(n1099) );
  CLKBUF_X1 U1041 ( .A(n1138), .Z(n1100) );
  CLKBUF_X1 U1042 ( .A(n1138), .Z(n1101) );
  CLKBUF_X1 U1043 ( .A(n1138), .Z(n1102) );
  CLKBUF_X1 U1044 ( .A(n1137), .Z(n1103) );
  CLKBUF_X1 U1045 ( .A(n1137), .Z(n1104) );
  CLKBUF_X1 U1046 ( .A(n1137), .Z(n1105) );
  CLKBUF_X1 U1047 ( .A(n1137), .Z(n1106) );
  CLKBUF_X1 U1048 ( .A(n1137), .Z(n1107) );
  CLKBUF_X1 U1049 ( .A(n1137), .Z(n1108) );
  CLKBUF_X1 U1050 ( .A(n1136), .Z(n1109) );
  CLKBUF_X1 U1051 ( .A(n1136), .Z(n1110) );
  CLKBUF_X1 U1052 ( .A(n1136), .Z(n1111) );
  CLKBUF_X1 U1053 ( .A(n1136), .Z(n1112) );
  CLKBUF_X1 U1054 ( .A(n1136), .Z(n1113) );
  CLKBUF_X1 U1055 ( .A(n1136), .Z(n1114) );
  CLKBUF_X1 U1056 ( .A(n1135), .Z(n1115) );
  CLKBUF_X1 U1057 ( .A(n1135), .Z(n1116) );
  CLKBUF_X1 U1058 ( .A(n1135), .Z(n1117) );
  CLKBUF_X1 U1059 ( .A(n1135), .Z(n1118) );
  CLKBUF_X1 U1060 ( .A(n1135), .Z(n1119) );
  CLKBUF_X1 U1061 ( .A(n1135), .Z(n1120) );
  CLKBUF_X1 U1062 ( .A(n1134), .Z(n1121) );
  CLKBUF_X1 U1063 ( .A(n1134), .Z(n1122) );
  CLKBUF_X1 U1064 ( .A(n1134), .Z(n1123) );
  CLKBUF_X1 U1065 ( .A(n1134), .Z(n1124) );
  CLKBUF_X1 U1066 ( .A(n1134), .Z(n1125) );
  CLKBUF_X1 U1067 ( .A(n1134), .Z(n1126) );
  CLKBUF_X1 U1068 ( .A(n1133), .Z(n1127) );
  CLKBUF_X1 U1069 ( .A(n1133), .Z(n1128) );
  CLKBUF_X1 U1070 ( .A(n1133), .Z(n1129) );
  CLKBUF_X1 U1071 ( .A(n1133), .Z(n1130) );
  CLKBUF_X1 U1072 ( .A(n1133), .Z(n1131) );
  CLKBUF_X1 U1073 ( .A(n1133), .Z(n1132) );
  INV_X1 U1074 ( .A(DP_y_23), .ZN(n1140) );
  NOR2_X1 U1075 ( .A1(DP_y_11_), .A2(n1140), .ZN(DP_N4) );
  INV_X1 U1076 ( .A(DP_y_11_), .ZN(n1141) );
  NOR2_X1 U1077 ( .A1(DP_y_23), .A2(n1141), .ZN(DP_N2) );
endmodule

